module rvecc_encode(
  input  [31:0] io_din,
  output [6:0]  io_ecc_out
);
  wire  w0_0 = io_din[0]; // @[el2_lib.scala 294:39]
  wire  w0_1 = io_din[1]; // @[el2_lib.scala 294:39]
  wire  w1_1 = io_din[2]; // @[el2_lib.scala 295:39]
  wire  w0_2 = io_din[3]; // @[el2_lib.scala 294:39]
  wire  w0_3 = io_din[4]; // @[el2_lib.scala 294:39]
  wire  w1_3 = io_din[5]; // @[el2_lib.scala 295:39]
  wire  w0_4 = io_din[6]; // @[el2_lib.scala 294:39]
  wire  w2_3 = io_din[7]; // @[el2_lib.scala 296:39]
  wire  w0_5 = io_din[8]; // @[el2_lib.scala 294:39]
  wire  w1_5 = io_din[9]; // @[el2_lib.scala 295:39]
  wire  w0_6 = io_din[10]; // @[el2_lib.scala 294:39]
  wire  w0_7 = io_din[11]; // @[el2_lib.scala 294:39]
  wire  w1_7 = io_din[12]; // @[el2_lib.scala 295:39]
  wire  w0_8 = io_din[13]; // @[el2_lib.scala 294:39]
  wire  w2_7 = io_din[14]; // @[el2_lib.scala 296:39]
  wire  w0_9 = io_din[15]; // @[el2_lib.scala 294:39]
  wire  w1_9 = io_din[16]; // @[el2_lib.scala 295:39]
  wire  w0_10 = io_din[17]; // @[el2_lib.scala 294:39]
  wire  w3_7 = io_din[18]; // @[el2_lib.scala 297:39]
  wire  w0_11 = io_din[19]; // @[el2_lib.scala 294:39]
  wire  w1_11 = io_din[20]; // @[el2_lib.scala 295:39]
  wire  w0_12 = io_din[21]; // @[el2_lib.scala 294:39]
  wire  w2_11 = io_din[22]; // @[el2_lib.scala 296:39]
  wire  w0_13 = io_din[23]; // @[el2_lib.scala 294:39]
  wire  w1_13 = io_din[24]; // @[el2_lib.scala 295:39]
  wire  w0_14 = io_din[25]; // @[el2_lib.scala 294:39]
  wire  w0_15 = io_din[26]; // @[el2_lib.scala 294:39]
  wire  w1_15 = io_din[27]; // @[el2_lib.scala 295:39]
  wire  w0_16 = io_din[28]; // @[el2_lib.scala 294:39]
  wire  w2_15 = io_din[29]; // @[el2_lib.scala 296:39]
  wire  w0_17 = io_din[30]; // @[el2_lib.scala 294:39]
  wire  w1_17 = io_din[31]; // @[el2_lib.scala 295:39]
  wire [5:0] _T_94 = {w1_17,w0_17,w2_15,w0_16,w1_15,w0_15}; // @[el2_lib.scala 301:22]
  wire  _T_95 = ^_T_94; // @[el2_lib.scala 301:29]
  wire [6:0] _T_101 = {w0_10,w1_9,w0_9,w2_7,w0_8,w1_7,w0_7}; // @[el2_lib.scala 301:39]
  wire [14:0] _T_109 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_101}; // @[el2_lib.scala 301:39]
  wire  _T_110 = ^_T_109; // @[el2_lib.scala 301:46]
  wire [6:0] _T_116 = {w0_6,w1_5,w0_5,w2_3,w0_4,w1_3,w0_3}; // @[el2_lib.scala 301:56]
  wire [14:0] _T_124 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_116}; // @[el2_lib.scala 301:56]
  wire  _T_125 = ^_T_124; // @[el2_lib.scala 301:63]
  wire [8:0] _T_133 = {w0_9,w2_7,w0_6,w1_5,w0_5,w2_3,w0_2,w1_1,w0_1}; // @[el2_lib.scala 301:73]
  wire [17:0] _T_142 = {w1_17,w0_17,w2_15,w0_14,w1_13,w0_13,w2_11,w0_10,w1_9,_T_133}; // @[el2_lib.scala 301:73]
  wire  _T_143 = ^_T_142; // @[el2_lib.scala 301:80]
  wire [8:0] _T_151 = {w0_8,w1_7,w0_6,w1_5,w0_4,w1_3,w0_2,w1_1,w0_0}; // @[el2_lib.scala 301:90]
  wire [17:0] _T_160 = {w1_17,w0_16,w1_15,w0_14,w1_13,w0_12,w1_11,w0_10,w1_9,_T_151}; // @[el2_lib.scala 301:90]
  wire  _T_161 = ^_T_160; // @[el2_lib.scala 301:97]
  wire [8:0] _T_169 = {w0_8,w0_7,w0_6,w0_5,w0_4,w0_3,w0_2,w0_1,w0_0}; // @[el2_lib.scala 301:107]
  wire [17:0] _T_178 = {w0_17,w0_16,w0_15,w0_14,w0_13,w0_12,w0_11,w0_10,w0_9,_T_169}; // @[el2_lib.scala 301:107]
  wire  _T_179 = ^_T_178; // @[el2_lib.scala 301:114]
  wire [5:0] w6 = {_T_95,_T_110,_T_125,_T_143,_T_161,_T_179}; // @[Cat.scala 29:58]
  wire  _T_184 = ^io_din; // @[el2_lib.scala 302:30]
  wire  _T_185 = ^w6; // @[el2_lib.scala 302:40]
  wire  _T_186 = _T_184 ^ _T_185; // @[el2_lib.scala 302:35]
  assign io_ecc_out = {_T_186,w6}; // @[el2_lib.scala 302:16]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [63:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] m1_io_din; // @[el2_ifu_mem_ctl.scala 635:18]
  wire [6:0] m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 635:18]
  wire [31:0] m2_io_din; // @[el2_ifu_mem_ctl.scala 637:18]
  wire [6:0] m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 637:18]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 184:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 319:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 320:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 320:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 252:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 546:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 548:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 186:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 307:34]
  wire [4:0] _GEN_464 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 667:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_464 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 667:53]
  wire [1:0] _GEN_465 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 670:91]
  wire [1:0] _T_2731 = ic_fetch_val_shift_right[3:2] & _GEN_465; // @[el2_ifu_mem_ctl.scala 670:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 321:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 274:46]
  wire [1:0] _GEN_466 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 670:113]
  wire [1:0] _T_2732 = _T_2731 & _GEN_466; // @[el2_ifu_mem_ctl.scala 670:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 656:59]
  wire [1:0] _GEN_467 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 670:130]
  wire [1:0] _T_2733 = _T_2732 | _GEN_467; // @[el2_ifu_mem_ctl.scala 670:130]
  wire  _T_2734 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 670:154]
  wire [1:0] _GEN_468 = {{1'd0}, _T_2734}; // @[el2_ifu_mem_ctl.scala 670:152]
  wire [1:0] _T_2735 = _T_2733 & _GEN_468; // @[el2_ifu_mem_ctl.scala 670:152]
  wire [1:0] _T_2724 = ic_fetch_val_shift_right[1:0] & _GEN_465; // @[el2_ifu_mem_ctl.scala 670:91]
  wire [1:0] _T_2725 = _T_2724 & _GEN_466; // @[el2_ifu_mem_ctl.scala 670:113]
  wire [1:0] _T_2726 = _T_2725 | _GEN_467; // @[el2_ifu_mem_ctl.scala 670:130]
  wire [1:0] _T_2728 = _T_2726 & _GEN_468; // @[el2_ifu_mem_ctl.scala 670:152]
  wire [3:0] iccm_ecc_word_enable = {_T_2735,_T_2728}; // @[Cat.scala 29:58]
  wire  _T_2835 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 334:30]
  wire  _T_2836 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 334:44]
  wire  _T_2837 = _T_2835 ^ _T_2836; // @[el2_lib.scala 334:35]
  wire [5:0] _T_2845 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 334:76]
  wire  _T_2846 = ^_T_2845; // @[el2_lib.scala 334:83]
  wire  _T_2847 = io_iccm_rd_data_ecc[37] ^ _T_2846; // @[el2_lib.scala 334:71]
  wire [6:0] _T_2854 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 334:103]
  wire [14:0] _T_2862 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2854}; // @[el2_lib.scala 334:103]
  wire  _T_2863 = ^_T_2862; // @[el2_lib.scala 334:110]
  wire  _T_2864 = io_iccm_rd_data_ecc[36] ^ _T_2863; // @[el2_lib.scala 334:98]
  wire [6:0] _T_2871 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 334:130]
  wire [14:0] _T_2879 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2871}; // @[el2_lib.scala 334:130]
  wire  _T_2880 = ^_T_2879; // @[el2_lib.scala 334:137]
  wire  _T_2881 = io_iccm_rd_data_ecc[35] ^ _T_2880; // @[el2_lib.scala 334:125]
  wire [8:0] _T_2890 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 334:157]
  wire [17:0] _T_2899 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2890}; // @[el2_lib.scala 334:157]
  wire  _T_2900 = ^_T_2899; // @[el2_lib.scala 334:164]
  wire  _T_2901 = io_iccm_rd_data_ecc[34] ^ _T_2900; // @[el2_lib.scala 334:152]
  wire [8:0] _T_2910 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 334:184]
  wire [17:0] _T_2919 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2910}; // @[el2_lib.scala 334:184]
  wire  _T_2920 = ^_T_2919; // @[el2_lib.scala 334:191]
  wire  _T_2921 = io_iccm_rd_data_ecc[33] ^ _T_2920; // @[el2_lib.scala 334:179]
  wire [8:0] _T_2930 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 334:211]
  wire [17:0] _T_2939 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_2930}; // @[el2_lib.scala 334:211]
  wire  _T_2940 = ^_T_2939; // @[el2_lib.scala 334:218]
  wire  _T_2941 = io_iccm_rd_data_ecc[32] ^ _T_2940; // @[el2_lib.scala 334:206]
  wire [6:0] _T_2947 = {_T_2837,_T_2847,_T_2864,_T_2881,_T_2901,_T_2921,_T_2941}; // @[Cat.scala 29:58]
  wire  _T_2948 = _T_2947 != 7'h0; // @[el2_lib.scala 335:44]
  wire  _T_2949 = iccm_ecc_word_enable[0] & _T_2948; // @[el2_lib.scala 335:32]
  wire  _T_2951 = _T_2949 & _T_2947[6]; // @[el2_lib.scala 335:53]
  wire  _T_3220 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 334:30]
  wire  _T_3221 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 334:44]
  wire  _T_3222 = _T_3220 ^ _T_3221; // @[el2_lib.scala 334:35]
  wire [5:0] _T_3230 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 334:76]
  wire  _T_3231 = ^_T_3230; // @[el2_lib.scala 334:83]
  wire  _T_3232 = io_iccm_rd_data_ecc[76] ^ _T_3231; // @[el2_lib.scala 334:71]
  wire [6:0] _T_3239 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 334:103]
  wire [14:0] _T_3247 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3239}; // @[el2_lib.scala 334:103]
  wire  _T_3248 = ^_T_3247; // @[el2_lib.scala 334:110]
  wire  _T_3249 = io_iccm_rd_data_ecc[75] ^ _T_3248; // @[el2_lib.scala 334:98]
  wire [6:0] _T_3256 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 334:130]
  wire [14:0] _T_3264 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3256}; // @[el2_lib.scala 334:130]
  wire  _T_3265 = ^_T_3264; // @[el2_lib.scala 334:137]
  wire  _T_3266 = io_iccm_rd_data_ecc[74] ^ _T_3265; // @[el2_lib.scala 334:125]
  wire [8:0] _T_3275 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 334:157]
  wire [17:0] _T_3284 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3275}; // @[el2_lib.scala 334:157]
  wire  _T_3285 = ^_T_3284; // @[el2_lib.scala 334:164]
  wire  _T_3286 = io_iccm_rd_data_ecc[73] ^ _T_3285; // @[el2_lib.scala 334:152]
  wire [8:0] _T_3295 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 334:184]
  wire [17:0] _T_3304 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3295}; // @[el2_lib.scala 334:184]
  wire  _T_3305 = ^_T_3304; // @[el2_lib.scala 334:191]
  wire  _T_3306 = io_iccm_rd_data_ecc[72] ^ _T_3305; // @[el2_lib.scala 334:179]
  wire [8:0] _T_3315 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 334:211]
  wire [17:0] _T_3324 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3315}; // @[el2_lib.scala 334:211]
  wire  _T_3325 = ^_T_3324; // @[el2_lib.scala 334:218]
  wire  _T_3326 = io_iccm_rd_data_ecc[71] ^ _T_3325; // @[el2_lib.scala 334:206]
  wire [6:0] _T_3332 = {_T_3222,_T_3232,_T_3249,_T_3266,_T_3286,_T_3306,_T_3326}; // @[Cat.scala 29:58]
  wire  _T_3333 = _T_3332 != 7'h0; // @[el2_lib.scala 335:44]
  wire  _T_3334 = iccm_ecc_word_enable[1] & _T_3333; // @[el2_lib.scala 335:32]
  wire  _T_3336 = _T_3334 & _T_3332[6]; // @[el2_lib.scala 335:53]
  wire [1:0] iccm_single_ecc_error = {_T_2951,_T_3336}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 189:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 630:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 190:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 191:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 475:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 191:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 191:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 191:72]
  wire  _T_2490 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2495 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2515 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 525:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 389:42]
  wire  _T_2517 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 525:79]
  wire  _T_2518 = _T_2515 | _T_2517; // @[el2_ifu_mem_ctl.scala 525:56]
  wire  _T_2519 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 525:122]
  wire  _T_2520 = ~_T_2519; // @[el2_ifu_mem_ctl.scala 525:101]
  wire  _T_2521 = _T_2518 & _T_2520; // @[el2_ifu_mem_ctl.scala 525:99]
  wire  _T_2522 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2536 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 532:45]
  wire  _T_2537 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 532:69]
  wire  _T_2538 = _T_2536 & _T_2537; // @[el2_ifu_mem_ctl.scala 532:67]
  wire  _T_2539 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_2522 ? _T_2538 : _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2495 ? _T_2521 : _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2490 ? 1'h0 : _GEN_59; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 191:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 193:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 193:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 282:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 282:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 702:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 282:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 273:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 273:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 323:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 273:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 273:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 282:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 282:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 282:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 282:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 282:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 545:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 587:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 614:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 309:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 595:56]
  wire  _T_2641 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 612:69]
  wire  _T_2642 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 612:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2641 : _T_2642; // @[el2_ifu_mem_ctl.scala 612:28]
  wire  _T_2588 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 591:68]
  wire  _T_2589 = ic_act_miss_f | _T_2588; // @[el2_ifu_mem_ctl.scala 591:48]
  wire  bus_reset_data_beat_cnt = _T_2589 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 591:91]
  wire  _T_2585 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 590:50]
  wire  _T_2586 = bus_ifu_wr_en_ff & _T_2585; // @[el2_ifu_mem_ctl.scala 590:48]
  wire  _T_2587 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 590:72]
  wire  bus_inc_data_beat_cnt = _T_2586 & _T_2587; // @[el2_ifu_mem_ctl.scala 590:70]
  wire [2:0] _T_2593 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 594:115]
  wire [2:0] _T_2595 = bus_inc_data_beat_cnt ? _T_2593 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2590 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 592:32]
  wire  _T_2591 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 592:57]
  wire  bus_hold_data_beat_cnt = _T_2590 & _T_2591; // @[el2_ifu_mem_ctl.scala 592:55]
  wire [2:0] _T_2596 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2595 | _T_2596; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 193:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 193:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 194:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 193:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 194:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 200:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 200:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 425:45]
  wire  _T_2120 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 446:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 402:60]
  wire  _T_2151 = _T_2120 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2124 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 446:127]
  wire  _T_2152 = _T_2124 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2159 = _T_2151 | _T_2152; // @[Mux.scala 27:72]
  wire  _T_2128 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 446:127]
  wire  _T_2153 = _T_2128 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2160 = _T_2159 | _T_2153; // @[Mux.scala 27:72]
  wire  _T_2132 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 446:127]
  wire  _T_2154 = _T_2132 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2161 = _T_2160 | _T_2154; // @[Mux.scala 27:72]
  wire  _T_2136 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 446:127]
  wire  _T_2155 = _T_2136 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2162 = _T_2161 | _T_2155; // @[Mux.scala 27:72]
  wire  _T_2140 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 446:127]
  wire  _T_2156 = _T_2140 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2163 = _T_2162 | _T_2156; // @[Mux.scala 27:72]
  wire  _T_2144 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 446:127]
  wire  _T_2157 = _T_2144 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2164 = _T_2163 | _T_2157; // @[Mux.scala 27:72]
  wire  _T_2148 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 446:127]
  wire  _T_2158 = _T_2148 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2164 | _T_2158; // @[Mux.scala 27:72]
  wire  _T_2206 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 448:69]
  wire  _T_2207 = ic_miss_buff_data_valid_bypass_index & _T_2206; // @[el2_ifu_mem_ctl.scala 448:67]
  wire  _T_2209 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 448:91]
  wire  _T_2210 = _T_2207 & _T_2209; // @[el2_ifu_mem_ctl.scala 448:89]
  wire  _T_2215 = _T_2207 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 449:65]
  wire  _T_2216 = _T_2210 | _T_2215; // @[el2_ifu_mem_ctl.scala 448:112]
  wire  _T_2218 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 450:43]
  wire  _T_2221 = _T_2218 & _T_2209; // @[el2_ifu_mem_ctl.scala 450:65]
  wire  _T_2222 = _T_2216 | _T_2221; // @[el2_ifu_mem_ctl.scala 449:88]
  wire  _T_2226 = _T_2218 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 451:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 428:75]
  wire  _T_2166 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2190 = _T_2166 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2169 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2191 = _T_2169 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2190 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2172 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2192 = _T_2172 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2199 = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2193 = _T_2175 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2199 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2178 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2194 = _T_2178 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2181 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2195 = _T_2181 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2184 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2196 = _T_2184 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2187 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 447:110]
  wire  _T_2197 = _T_2187 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2227 = _T_2226 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 451:87]
  wire  _T_2228 = _T_2222 | _T_2227; // @[el2_ifu_mem_ctl.scala 450:88]
  wire  _T_2232 = ic_miss_buff_data_valid_bypass_index & _T_2148; // @[el2_ifu_mem_ctl.scala 452:43]
  wire  miss_buff_hit_unq_f = _T_2228 | _T_2232; // @[el2_ifu_mem_ctl.scala 451:131]
  wire  _T_2248 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 457:55]
  wire  _T_2249 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 457:87]
  wire  _T_2250 = _T_2248 | _T_2249; // @[el2_ifu_mem_ctl.scala 457:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2250; // @[el2_ifu_mem_ctl.scala 457:41]
  wire  _T_2233 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 454:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 310:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 445:51]
  wire  _T_2234 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 454:68]
  wire  _T_2235 = miss_buff_hit_unq_f & _T_2234; // @[el2_ifu_mem_ctl.scala 454:66]
  wire  stream_hit_f = _T_2233 & _T_2235; // @[el2_ifu_mem_ctl.scala 454:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 277:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 277:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 277:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 597:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 624:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 204:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 204:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 204:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 204:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 204:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 205:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 206:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 206:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 207:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 208:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 208:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 208:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 196:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 208:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 208:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 208:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 209:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 209:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 209:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 209:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 210:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 211:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 211:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 211:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 209:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 208:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 207:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 206:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 205:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 204:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2245 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 456:60]
  wire  _T_2246 = _T_2245 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 456:94]
  wire  stream_eol_f = _T_2246 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 456:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 219:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 219:87]
  wire  _T_113 = _T_111 & _T_2587; // @[el2_ifu_mem_ctl.scala 219:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 219:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 223:48]
  wire  _T_126 = _T_124 & _T_2587; // @[el2_ifu_mem_ctl.scala 223:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 223:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 283:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 283:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 283:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 283:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 284:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 283:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 284:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 337:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 284:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 284:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 284:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 227:50]
  wire  _T_137 = _T_135 & _T_2587; // @[el2_ifu_mem_ctl.scala 227:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 285:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 286:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 285:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:35]
  wire  _T_143 = _T_141 & _T_2587; // @[el2_ifu_mem_ctl.scala 228:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 228:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 227:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 233:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 232:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 232:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 237:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 237:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 194:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 194:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 194:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 194:91]
  wire  _T_30 = ic_act_miss_f & _T_2587; // @[el2_ifu_mem_ctl.scala 201:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 212:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 212:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 212:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 212:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 212:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 216:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 216:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 216:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 220:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 220:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 224:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 224:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 229:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 229:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 229:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 234:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 234:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 253:95]
  wire  _T_175 = _T_2248 & _T_174; // @[el2_ifu_mem_ctl.scala 253:93]
  wire  crit_wd_byp_ok_ff = _T_2249 | _T_175; // @[el2_ifu_mem_ctl.scala 253:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 254:36]
  wire  _T_180 = _T_2248 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 254:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 254:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 254:70]
  wire  _T_184 = _T_2248 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 255:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 255:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 254:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 255:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 256:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 256:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 255:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 258:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 258:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 266:35]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 736:14]
  wire  _T_4399 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_4527 = _T_4399 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4400 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_4528 = _T_4400 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_4655 = _T_4527 | _T_4528; // @[Mux.scala 27:72]
  wire  _T_4401 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_4529 = _T_4401 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_4656 = _T_4655 | _T_4529; // @[Mux.scala 27:72]
  wire  _T_4402 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_4530 = _T_4402 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_4657 = _T_4656 | _T_4530; // @[Mux.scala 27:72]
  wire  _T_4403 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_4531 = _T_4403 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_4658 = _T_4657 | _T_4531; // @[Mux.scala 27:72]
  wire  _T_4404 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_4532 = _T_4404 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_4659 = _T_4658 | _T_4532; // @[Mux.scala 27:72]
  wire  _T_4405 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_4533 = _T_4405 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_4660 = _T_4659 | _T_4533; // @[Mux.scala 27:72]
  wire  _T_4406 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_4534 = _T_4406 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_4661 = _T_4660 | _T_4534; // @[Mux.scala 27:72]
  wire  _T_4407 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_4535 = _T_4407 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_4662 = _T_4661 | _T_4535; // @[Mux.scala 27:72]
  wire  _T_4408 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_4536 = _T_4408 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_4663 = _T_4662 | _T_4536; // @[Mux.scala 27:72]
  wire  _T_4409 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_4537 = _T_4409 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_4664 = _T_4663 | _T_4537; // @[Mux.scala 27:72]
  wire  _T_4410 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_4538 = _T_4410 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_4665 = _T_4664 | _T_4538; // @[Mux.scala 27:72]
  wire  _T_4411 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_4539 = _T_4411 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_4666 = _T_4665 | _T_4539; // @[Mux.scala 27:72]
  wire  _T_4412 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_4540 = _T_4412 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_4667 = _T_4666 | _T_4540; // @[Mux.scala 27:72]
  wire  _T_4413 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_4541 = _T_4413 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_4668 = _T_4667 | _T_4541; // @[Mux.scala 27:72]
  wire  _T_4414 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_4542 = _T_4414 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_4669 = _T_4668 | _T_4542; // @[Mux.scala 27:72]
  wire  _T_4415 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_4543 = _T_4415 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_4670 = _T_4669 | _T_4543; // @[Mux.scala 27:72]
  wire  _T_4416 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_4544 = _T_4416 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_4671 = _T_4670 | _T_4544; // @[Mux.scala 27:72]
  wire  _T_4417 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_4545 = _T_4417 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_4672 = _T_4671 | _T_4545; // @[Mux.scala 27:72]
  wire  _T_4418 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_4546 = _T_4418 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_4673 = _T_4672 | _T_4546; // @[Mux.scala 27:72]
  wire  _T_4419 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_4547 = _T_4419 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_4674 = _T_4673 | _T_4547; // @[Mux.scala 27:72]
  wire  _T_4420 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_4548 = _T_4420 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_4675 = _T_4674 | _T_4548; // @[Mux.scala 27:72]
  wire  _T_4421 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_4549 = _T_4421 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_4676 = _T_4675 | _T_4549; // @[Mux.scala 27:72]
  wire  _T_4422 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_4550 = _T_4422 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_4677 = _T_4676 | _T_4550; // @[Mux.scala 27:72]
  wire  _T_4423 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_4551 = _T_4423 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_4678 = _T_4677 | _T_4551; // @[Mux.scala 27:72]
  wire  _T_4424 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_4552 = _T_4424 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_4679 = _T_4678 | _T_4552; // @[Mux.scala 27:72]
  wire  _T_4425 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_4553 = _T_4425 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_4680 = _T_4679 | _T_4553; // @[Mux.scala 27:72]
  wire  _T_4426 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_4554 = _T_4426 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_4681 = _T_4680 | _T_4554; // @[Mux.scala 27:72]
  wire  _T_4427 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_4555 = _T_4427 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_4682 = _T_4681 | _T_4555; // @[Mux.scala 27:72]
  wire  _T_4428 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_4556 = _T_4428 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_4683 = _T_4682 | _T_4556; // @[Mux.scala 27:72]
  wire  _T_4429 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_4557 = _T_4429 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_4684 = _T_4683 | _T_4557; // @[Mux.scala 27:72]
  wire  _T_4430 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_4558 = _T_4430 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_4685 = _T_4684 | _T_4558; // @[Mux.scala 27:72]
  wire  _T_4431 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_4559 = _T_4431 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_4686 = _T_4685 | _T_4559; // @[Mux.scala 27:72]
  wire  _T_4432 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_4560 = _T_4432 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_4687 = _T_4686 | _T_4560; // @[Mux.scala 27:72]
  wire  _T_4433 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_4561 = _T_4433 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_4688 = _T_4687 | _T_4561; // @[Mux.scala 27:72]
  wire  _T_4434 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_4562 = _T_4434 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_4689 = _T_4688 | _T_4562; // @[Mux.scala 27:72]
  wire  _T_4435 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_4563 = _T_4435 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_4690 = _T_4689 | _T_4563; // @[Mux.scala 27:72]
  wire  _T_4436 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_4564 = _T_4436 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_4691 = _T_4690 | _T_4564; // @[Mux.scala 27:72]
  wire  _T_4437 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_4565 = _T_4437 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_4692 = _T_4691 | _T_4565; // @[Mux.scala 27:72]
  wire  _T_4438 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_4566 = _T_4438 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_4693 = _T_4692 | _T_4566; // @[Mux.scala 27:72]
  wire  _T_4439 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_4567 = _T_4439 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_4694 = _T_4693 | _T_4567; // @[Mux.scala 27:72]
  wire  _T_4440 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_4568 = _T_4440 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_4695 = _T_4694 | _T_4568; // @[Mux.scala 27:72]
  wire  _T_4441 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_4569 = _T_4441 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_4696 = _T_4695 | _T_4569; // @[Mux.scala 27:72]
  wire  _T_4442 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_4570 = _T_4442 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_4697 = _T_4696 | _T_4570; // @[Mux.scala 27:72]
  wire  _T_4443 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_4571 = _T_4443 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_4698 = _T_4697 | _T_4571; // @[Mux.scala 27:72]
  wire  _T_4444 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_4572 = _T_4444 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_4699 = _T_4698 | _T_4572; // @[Mux.scala 27:72]
  wire  _T_4445 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_4573 = _T_4445 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_4700 = _T_4699 | _T_4573; // @[Mux.scala 27:72]
  wire  _T_4446 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_4574 = _T_4446 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_4701 = _T_4700 | _T_4574; // @[Mux.scala 27:72]
  wire  _T_4447 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_4575 = _T_4447 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_4702 = _T_4701 | _T_4575; // @[Mux.scala 27:72]
  wire  _T_4448 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_4576 = _T_4448 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_4703 = _T_4702 | _T_4576; // @[Mux.scala 27:72]
  wire  _T_4449 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_4577 = _T_4449 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_4704 = _T_4703 | _T_4577; // @[Mux.scala 27:72]
  wire  _T_4450 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_4578 = _T_4450 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_4705 = _T_4704 | _T_4578; // @[Mux.scala 27:72]
  wire  _T_4451 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_4579 = _T_4451 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_4706 = _T_4705 | _T_4579; // @[Mux.scala 27:72]
  wire  _T_4452 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_4580 = _T_4452 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_4707 = _T_4706 | _T_4580; // @[Mux.scala 27:72]
  wire  _T_4453 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_4581 = _T_4453 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_4708 = _T_4707 | _T_4581; // @[Mux.scala 27:72]
  wire  _T_4454 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_4582 = _T_4454 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_4709 = _T_4708 | _T_4582; // @[Mux.scala 27:72]
  wire  _T_4455 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_4583 = _T_4455 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_4710 = _T_4709 | _T_4583; // @[Mux.scala 27:72]
  wire  _T_4456 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_4584 = _T_4456 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_4711 = _T_4710 | _T_4584; // @[Mux.scala 27:72]
  wire  _T_4457 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_4585 = _T_4457 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_4712 = _T_4711 | _T_4585; // @[Mux.scala 27:72]
  wire  _T_4458 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_4586 = _T_4458 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_4713 = _T_4712 | _T_4586; // @[Mux.scala 27:72]
  wire  _T_4459 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_4587 = _T_4459 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_4714 = _T_4713 | _T_4587; // @[Mux.scala 27:72]
  wire  _T_4460 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_4588 = _T_4460 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_4715 = _T_4714 | _T_4588; // @[Mux.scala 27:72]
  wire  _T_4461 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_4589 = _T_4461 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_4716 = _T_4715 | _T_4589; // @[Mux.scala 27:72]
  wire  _T_4462 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_4590 = _T_4462 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_4717 = _T_4716 | _T_4590; // @[Mux.scala 27:72]
  wire  _T_4463 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_4591 = _T_4463 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_4718 = _T_4717 | _T_4591; // @[Mux.scala 27:72]
  wire  _T_4464 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_4592 = _T_4464 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_4719 = _T_4718 | _T_4592; // @[Mux.scala 27:72]
  wire  _T_4465 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_4593 = _T_4465 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_4720 = _T_4719 | _T_4593; // @[Mux.scala 27:72]
  wire  _T_4466 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_4594 = _T_4466 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_4721 = _T_4720 | _T_4594; // @[Mux.scala 27:72]
  wire  _T_4467 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_4595 = _T_4467 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_4722 = _T_4721 | _T_4595; // @[Mux.scala 27:72]
  wire  _T_4468 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_4596 = _T_4468 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_4723 = _T_4722 | _T_4596; // @[Mux.scala 27:72]
  wire  _T_4469 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_4597 = _T_4469 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_4724 = _T_4723 | _T_4597; // @[Mux.scala 27:72]
  wire  _T_4470 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_4598 = _T_4470 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_4725 = _T_4724 | _T_4598; // @[Mux.scala 27:72]
  wire  _T_4471 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_4599 = _T_4471 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_4726 = _T_4725 | _T_4599; // @[Mux.scala 27:72]
  wire  _T_4472 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_4600 = _T_4472 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_4727 = _T_4726 | _T_4600; // @[Mux.scala 27:72]
  wire  _T_4473 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_4601 = _T_4473 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_4728 = _T_4727 | _T_4601; // @[Mux.scala 27:72]
  wire  _T_4474 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_4602 = _T_4474 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_4729 = _T_4728 | _T_4602; // @[Mux.scala 27:72]
  wire  _T_4475 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_4603 = _T_4475 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_4730 = _T_4729 | _T_4603; // @[Mux.scala 27:72]
  wire  _T_4476 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_4604 = _T_4476 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_4731 = _T_4730 | _T_4604; // @[Mux.scala 27:72]
  wire  _T_4477 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_4605 = _T_4477 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_4732 = _T_4731 | _T_4605; // @[Mux.scala 27:72]
  wire  _T_4478 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_4606 = _T_4478 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_4733 = _T_4732 | _T_4606; // @[Mux.scala 27:72]
  wire  _T_4479 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_4607 = _T_4479 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_4734 = _T_4733 | _T_4607; // @[Mux.scala 27:72]
  wire  _T_4480 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_4608 = _T_4480 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_4735 = _T_4734 | _T_4608; // @[Mux.scala 27:72]
  wire  _T_4481 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_4609 = _T_4481 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_4736 = _T_4735 | _T_4609; // @[Mux.scala 27:72]
  wire  _T_4482 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_4610 = _T_4482 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_4737 = _T_4736 | _T_4610; // @[Mux.scala 27:72]
  wire  _T_4483 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_4611 = _T_4483 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_4738 = _T_4737 | _T_4611; // @[Mux.scala 27:72]
  wire  _T_4484 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_4612 = _T_4484 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_4739 = _T_4738 | _T_4612; // @[Mux.scala 27:72]
  wire  _T_4485 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_4613 = _T_4485 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_4740 = _T_4739 | _T_4613; // @[Mux.scala 27:72]
  wire  _T_4486 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_4614 = _T_4486 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_4741 = _T_4740 | _T_4614; // @[Mux.scala 27:72]
  wire  _T_4487 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_4615 = _T_4487 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_4742 = _T_4741 | _T_4615; // @[Mux.scala 27:72]
  wire  _T_4488 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_4616 = _T_4488 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_4743 = _T_4742 | _T_4616; // @[Mux.scala 27:72]
  wire  _T_4489 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_4617 = _T_4489 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_4744 = _T_4743 | _T_4617; // @[Mux.scala 27:72]
  wire  _T_4490 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_4618 = _T_4490 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_4745 = _T_4744 | _T_4618; // @[Mux.scala 27:72]
  wire  _T_4491 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_4619 = _T_4491 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_4746 = _T_4745 | _T_4619; // @[Mux.scala 27:72]
  wire  _T_4492 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_4620 = _T_4492 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_4747 = _T_4746 | _T_4620; // @[Mux.scala 27:72]
  wire  _T_4493 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_4621 = _T_4493 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_4748 = _T_4747 | _T_4621; // @[Mux.scala 27:72]
  wire  _T_4494 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_4622 = _T_4494 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_4749 = _T_4748 | _T_4622; // @[Mux.scala 27:72]
  wire  _T_4495 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_4623 = _T_4495 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_4750 = _T_4749 | _T_4623; // @[Mux.scala 27:72]
  wire  _T_4496 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_4624 = _T_4496 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_4751 = _T_4750 | _T_4624; // @[Mux.scala 27:72]
  wire  _T_4497 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_4625 = _T_4497 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_4752 = _T_4751 | _T_4625; // @[Mux.scala 27:72]
  wire  _T_4498 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_4626 = _T_4498 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_4753 = _T_4752 | _T_4626; // @[Mux.scala 27:72]
  wire  _T_4499 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_4627 = _T_4499 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_4754 = _T_4753 | _T_4627; // @[Mux.scala 27:72]
  wire  _T_4500 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_4628 = _T_4500 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_4755 = _T_4754 | _T_4628; // @[Mux.scala 27:72]
  wire  _T_4501 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_4629 = _T_4501 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_4756 = _T_4755 | _T_4629; // @[Mux.scala 27:72]
  wire  _T_4502 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_4630 = _T_4502 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_4757 = _T_4756 | _T_4630; // @[Mux.scala 27:72]
  wire  _T_4503 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_4631 = _T_4503 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_4758 = _T_4757 | _T_4631; // @[Mux.scala 27:72]
  wire  _T_4504 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_4632 = _T_4504 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_4759 = _T_4758 | _T_4632; // @[Mux.scala 27:72]
  wire  _T_4505 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_4633 = _T_4505 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_4760 = _T_4759 | _T_4633; // @[Mux.scala 27:72]
  wire  _T_4506 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_4634 = _T_4506 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_4761 = _T_4760 | _T_4634; // @[Mux.scala 27:72]
  wire  _T_4507 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_4635 = _T_4507 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_4762 = _T_4761 | _T_4635; // @[Mux.scala 27:72]
  wire  _T_4508 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_4636 = _T_4508 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_4763 = _T_4762 | _T_4636; // @[Mux.scala 27:72]
  wire  _T_4509 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_4637 = _T_4509 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_4764 = _T_4763 | _T_4637; // @[Mux.scala 27:72]
  wire  _T_4510 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_4638 = _T_4510 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_4765 = _T_4764 | _T_4638; // @[Mux.scala 27:72]
  wire  _T_4511 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_4639 = _T_4511 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_4766 = _T_4765 | _T_4639; // @[Mux.scala 27:72]
  wire  _T_4512 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_4640 = _T_4512 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_4767 = _T_4766 | _T_4640; // @[Mux.scala 27:72]
  wire  _T_4513 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_4641 = _T_4513 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_4768 = _T_4767 | _T_4641; // @[Mux.scala 27:72]
  wire  _T_4514 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_4642 = _T_4514 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_4769 = _T_4768 | _T_4642; // @[Mux.scala 27:72]
  wire  _T_4515 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_4643 = _T_4515 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_4770 = _T_4769 | _T_4643; // @[Mux.scala 27:72]
  wire  _T_4516 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_4644 = _T_4516 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_4771 = _T_4770 | _T_4644; // @[Mux.scala 27:72]
  wire  _T_4517 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_4645 = _T_4517 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_4772 = _T_4771 | _T_4645; // @[Mux.scala 27:72]
  wire  _T_4518 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_4646 = _T_4518 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_4773 = _T_4772 | _T_4646; // @[Mux.scala 27:72]
  wire  _T_4519 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_4647 = _T_4519 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_4774 = _T_4773 | _T_4647; // @[Mux.scala 27:72]
  wire  _T_4520 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_4648 = _T_4520 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_4775 = _T_4774 | _T_4648; // @[Mux.scala 27:72]
  wire  _T_4521 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_4649 = _T_4521 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_4776 = _T_4775 | _T_4649; // @[Mux.scala 27:72]
  wire  _T_4522 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_4650 = _T_4522 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_4777 = _T_4776 | _T_4650; // @[Mux.scala 27:72]
  wire  _T_4523 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_4651 = _T_4523 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_4778 = _T_4777 | _T_4651; // @[Mux.scala 27:72]
  wire  _T_4524 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_4652 = _T_4524 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_4779 = _T_4778 | _T_4652; // @[Mux.scala 27:72]
  wire  _T_4525 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_4653 = _T_4525 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_4780 = _T_4779 | _T_4653; // @[Mux.scala 27:72]
  wire  _T_4526 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 732:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_4654 = _T_4526 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_4780 | _T_4654; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 261:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 261:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:29]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 263:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 265:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 270:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 275:59]
  wire  _T_214 = _T_212 | _T_2233; // @[el2_ifu_mem_ctl.scala 275:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 275:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 281:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 281:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 281:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 281:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 288:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 288:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 288:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 289:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 289:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 292:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 292:135]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2662 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 620:48]
  wire  _T_2663 = _T_2662 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 620:52]
  wire  bus_ifu_wr_data_error_ff = _T_2663 & miss_pending; // @[el2_ifu_mem_ctl.scala 620:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 365:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 364:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 292:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 292:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 295:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 295:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 296:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 315:30]
  wire  _T_9988 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 788:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 316:24]
  wire  _T_9990 = _T_9988 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 788:51]
  wire  _T_9992 = _T_9990 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 788:67]
  wire  _T_9994 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 788:86]
  wire  replace_way_mb_any_0 = _T_9992 | _T_9994; // @[el2_ifu_mem_ctl.scala 788:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9997 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 789:50]
  wire  _T_9999 = _T_9997 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 789:66]
  wire  _T_10001 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 789:85]
  wire  _T_10003 = _T_10001 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 789:100]
  wire  replace_way_mb_any_1 = _T_9999 | _T_10003; // @[el2_ifu_mem_ctl.scala 789:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 300:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 300:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 301:56]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 304:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 304:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 305:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 304:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 304:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 306:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 314:23]
  wire  _T_313 = _T_2248 & flush_final_f; // @[el2_ifu_mem_ctl.scala 318:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 318:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 318:53]
  wire  _T_2240 = ~_T_2235; // @[el2_ifu_mem_ctl.scala 455:46]
  wire  _T_2241 = _T_2233 & _T_2240; // @[el2_ifu_mem_ctl.scala 455:44]
  wire  stream_miss_f = _T_2241 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 455:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 318:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 318:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 324:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_2233; // @[el2_ifu_mem_ctl.scala 326:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 326:82]
  wire  _T_2254 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 460:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2254}; // @[Cat.scala 29:58]
  wire  _T_2255 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2279 = _T_2255 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2258 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2280 = _T_2258 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2287 = _T_2279 | _T_2280; // @[Mux.scala 27:72]
  wire  _T_2261 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2281 = _T_2261 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2287 | _T_2281; // @[Mux.scala 27:72]
  wire  _T_2264 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2282 = _T_2264 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2288 | _T_2282; // @[Mux.scala 27:72]
  wire  _T_2267 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2283 = _T_2267 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2289 | _T_2283; // @[Mux.scala 27:72]
  wire  _T_2270 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2284 = _T_2270 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2290 | _T_2284; // @[Mux.scala 27:72]
  wire  _T_2273 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2285 = _T_2273 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2291 | _T_2285; // @[Mux.scala 27:72]
  wire  _T_2276 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 461:81]
  wire  _T_2286 = _T_2276 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2292 | _T_2286; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 462:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 330:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 330:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 617:61]
  wire  _T_2656 = ic_act_miss_f_delayed & _T_2249; // @[el2_ifu_mem_ctl.scala 618:53]
  wire  reset_tag_valid_for_miss = _T_2656 & _T_17; // @[el2_ifu_mem_ctl.scala 618:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 330:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 332:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 334:84]
  wire  _T_2650 = ~_T_2662; // @[el2_ifu_mem_ctl.scala 615:84]
  wire  _T_2651 = _T_100 & _T_2650; // @[el2_ifu_mem_ctl.scala 615:82]
  wire  bus_ifu_wr_en_ff_q = _T_2651 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 615:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 334:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 335:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_567 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 417:13]
  wire  _T_568 = ^_T_567; // @[el2_lib.scala 417:20]
  wire [6:0] _T_574 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 417:30]
  wire [7:0] _T_581 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 417:30]
  wire [14:0] _T_582 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_574}; // @[el2_lib.scala 417:30]
  wire [7:0] _T_589 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 417:30]
  wire [30:0] _T_598 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_582}; // @[el2_lib.scala 417:30]
  wire  _T_599 = ^_T_598; // @[el2_lib.scala 417:37]
  wire [6:0] _T_605 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 417:47]
  wire [14:0] _T_613 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_605}; // @[el2_lib.scala 417:47]
  wire [30:0] _T_629 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_613}; // @[el2_lib.scala 417:47]
  wire  _T_630 = ^_T_629; // @[el2_lib.scala 417:54]
  wire [6:0] _T_636 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 417:64]
  wire [14:0] _T_644 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_636}; // @[el2_lib.scala 417:64]
  wire [30:0] _T_660 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_581,_T_644}; // @[el2_lib.scala 417:64]
  wire  _T_661 = ^_T_660; // @[el2_lib.scala 417:71]
  wire [7:0] _T_668 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 417:81]
  wire [16:0] _T_677 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_668}; // @[el2_lib.scala 417:81]
  wire [8:0] _T_685 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 417:81]
  wire [17:0] _T_694 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_685}; // @[el2_lib.scala 417:81]
  wire [34:0] _T_695 = {_T_694,_T_677}; // @[el2_lib.scala 417:81]
  wire  _T_696 = ^_T_695; // @[el2_lib.scala 417:88]
  wire [7:0] _T_703 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 417:98]
  wire [16:0] _T_712 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_703}; // @[el2_lib.scala 417:98]
  wire [8:0] _T_720 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 417:98]
  wire [17:0] _T_729 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_720}; // @[el2_lib.scala 417:98]
  wire [34:0] _T_730 = {_T_729,_T_712}; // @[el2_lib.scala 417:98]
  wire  _T_731 = ^_T_730; // @[el2_lib.scala 417:105]
  wire [7:0] _T_738 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 417:115]
  wire [16:0] _T_747 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_738}; // @[el2_lib.scala 417:115]
  wire [8:0] _T_755 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 417:115]
  wire [17:0] _T_764 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_755}; // @[el2_lib.scala 417:115]
  wire [34:0] _T_765 = {_T_764,_T_747}; // @[el2_lib.scala 417:115]
  wire  _T_766 = ^_T_765; // @[el2_lib.scala 417:122]
  wire [3:0] _T_2295 = {ifu_bus_rid_ff[2:1],_T_2254,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2296 = _T_2295 == 4'h0; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2343 = _T_2296 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2299 = _T_2295 == 4'h1; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2344 = _T_2299 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2343 | _T_2344; // @[Mux.scala 27:72]
  wire  _T_2302 = _T_2295 == 4'h2; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2345 = _T_2302 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2360 = _T_2359 | _T_2345; // @[Mux.scala 27:72]
  wire  _T_2305 = _T_2295 == 4'h3; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2346 = _T_2305 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2360 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2308 = _T_2295 == 4'h4; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2347 = _T_2308 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire  _T_2311 = _T_2295 == 4'h5; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2348 = _T_2311 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2363 = _T_2362 | _T_2348; // @[Mux.scala 27:72]
  wire  _T_2314 = _T_2295 == 4'h6; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2349 = _T_2314 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2364 = _T_2363 | _T_2349; // @[Mux.scala 27:72]
  wire  _T_2317 = _T_2295 == 4'h7; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2350 = _T_2317 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2365 = _T_2364 | _T_2350; // @[Mux.scala 27:72]
  wire  _T_2320 = _T_2295 == 4'h8; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2351 = _T_2320 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2366 = _T_2365 | _T_2351; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2295 == 4'h9; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2352 = _T_2323 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2367 = _T_2366 | _T_2352; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2295 == 4'ha; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2353 = _T_2326 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2368 = _T_2367 | _T_2353; // @[Mux.scala 27:72]
  wire  _T_2329 = _T_2295 == 4'hb; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2354 = _T_2329 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2369 = _T_2368 | _T_2354; // @[Mux.scala 27:72]
  wire  _T_2332 = _T_2295 == 4'hc; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2355 = _T_2332 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 27:72]
  wire  _T_2335 = _T_2295 == 4'hd; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2356 = _T_2335 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2371 = _T_2370 | _T_2356; // @[Mux.scala 27:72]
  wire  _T_2338 = _T_2295 == 4'he; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2357 = _T_2338 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2372 = _T_2371 | _T_2357; // @[Mux.scala 27:72]
  wire  _T_2341 = _T_2295 == 4'hf; // @[el2_ifu_mem_ctl.scala 463:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2358 = _T_2341 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2373 = _T_2372 | _T_2358; // @[Mux.scala 27:72]
  wire [3:0] _T_2375 = {ifu_bus_rid_ff[2:1],_T_2254,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2376 = _T_2375 == 4'h0; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2423 = _T_2376 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2375 == 4'h1; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2424 = _T_2379 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2439 = _T_2423 | _T_2424; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2375 == 4'h2; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2425 = _T_2382 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2440 = _T_2439 | _T_2425; // @[Mux.scala 27:72]
  wire  _T_2385 = _T_2375 == 4'h3; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2426 = _T_2385 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2441 = _T_2440 | _T_2426; // @[Mux.scala 27:72]
  wire  _T_2388 = _T_2375 == 4'h4; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2427 = _T_2388 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2442 = _T_2441 | _T_2427; // @[Mux.scala 27:72]
  wire  _T_2391 = _T_2375 == 4'h5; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2428 = _T_2391 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2443 = _T_2442 | _T_2428; // @[Mux.scala 27:72]
  wire  _T_2394 = _T_2375 == 4'h6; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2429 = _T_2394 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2444 = _T_2443 | _T_2429; // @[Mux.scala 27:72]
  wire  _T_2397 = _T_2375 == 4'h7; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2430 = _T_2397 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2445 = _T_2444 | _T_2430; // @[Mux.scala 27:72]
  wire  _T_2400 = _T_2375 == 4'h8; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2431 = _T_2400 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2446 = _T_2445 | _T_2431; // @[Mux.scala 27:72]
  wire  _T_2403 = _T_2375 == 4'h9; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2432 = _T_2403 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2447 = _T_2446 | _T_2432; // @[Mux.scala 27:72]
  wire  _T_2406 = _T_2375 == 4'ha; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2433 = _T_2406 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2448 = _T_2447 | _T_2433; // @[Mux.scala 27:72]
  wire  _T_2409 = _T_2375 == 4'hb; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2434 = _T_2409 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2449 = _T_2448 | _T_2434; // @[Mux.scala 27:72]
  wire  _T_2412 = _T_2375 == 4'hc; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2435 = _T_2412 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2450 = _T_2449 | _T_2435; // @[Mux.scala 27:72]
  wire  _T_2415 = _T_2375 == 4'hd; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2436 = _T_2415 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2451 = _T_2450 | _T_2436; // @[Mux.scala 27:72]
  wire  _T_2418 = _T_2375 == 4'he; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2437 = _T_2418 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2452 = _T_2451 | _T_2437; // @[Mux.scala 27:72]
  wire  _T_2421 = _T_2375 == 4'hf; // @[el2_ifu_mem_ctl.scala 464:66]
  wire [31:0] _T_2438 = _T_2421 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2453 = _T_2452 | _T_2438; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [6:0] _T_989 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 417:13]
  wire  _T_990 = ^_T_989; // @[el2_lib.scala 417:20]
  wire [6:0] _T_996 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 417:30]
  wire [7:0] _T_1003 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 417:30]
  wire [14:0] _T_1004 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_996}; // @[el2_lib.scala 417:30]
  wire [7:0] _T_1011 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 417:30]
  wire [30:0] _T_1020 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1004}; // @[el2_lib.scala 417:30]
  wire  _T_1021 = ^_T_1020; // @[el2_lib.scala 417:37]
  wire [6:0] _T_1027 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 417:47]
  wire [14:0] _T_1035 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1027}; // @[el2_lib.scala 417:47]
  wire [30:0] _T_1051 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1035}; // @[el2_lib.scala 417:47]
  wire  _T_1052 = ^_T_1051; // @[el2_lib.scala 417:54]
  wire [6:0] _T_1058 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 417:64]
  wire [14:0] _T_1066 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1058}; // @[el2_lib.scala 417:64]
  wire [30:0] _T_1082 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1003,_T_1066}; // @[el2_lib.scala 417:64]
  wire  _T_1083 = ^_T_1082; // @[el2_lib.scala 417:71]
  wire [7:0] _T_1090 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 417:81]
  wire [16:0] _T_1099 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1090}; // @[el2_lib.scala 417:81]
  wire [8:0] _T_1107 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 417:81]
  wire [17:0] _T_1116 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1107}; // @[el2_lib.scala 417:81]
  wire [34:0] _T_1117 = {_T_1116,_T_1099}; // @[el2_lib.scala 417:81]
  wire  _T_1118 = ^_T_1117; // @[el2_lib.scala 417:88]
  wire [7:0] _T_1125 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 417:98]
  wire [16:0] _T_1134 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1125}; // @[el2_lib.scala 417:98]
  wire [8:0] _T_1142 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 417:98]
  wire [17:0] _T_1151 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1142}; // @[el2_lib.scala 417:98]
  wire [34:0] _T_1152 = {_T_1151,_T_1134}; // @[el2_lib.scala 417:98]
  wire  _T_1153 = ^_T_1152; // @[el2_lib.scala 417:105]
  wire [7:0] _T_1160 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 417:115]
  wire [16:0] _T_1169 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1160}; // @[el2_lib.scala 417:115]
  wire [8:0] _T_1177 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 417:115]
  wire [17:0] _T_1186 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1177}; // @[el2_lib.scala 417:115]
  wire [34:0] _T_1187 = {_T_1186,_T_1169}; // @[el2_lib.scala 417:115]
  wire  _T_1188 = ^_T_1187; // @[el2_lib.scala 417:122]
  wire [70:0] _T_1233 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1232 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [141:0] _T_1234 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff,_T_1232}; // @[Cat.scala 29:58]
  wire [141:0] _T_1237 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453,_T_1233}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1234 : _T_1237; // @[el2_ifu_mem_ctl.scala 356:28]
  wire  _T_1196 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 346:56]
  wire  _T_1197 = _T_1196 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 346:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 410:28]
  wire  _T_1413 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 613:35]
  wire  _T_1282 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1339 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 401:118]
  wire  _T_1340 = ic_miss_buff_data_valid[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1340; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1436 = _T_1413 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1343 = ic_miss_buff_data_valid[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1343; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1437 = _T_1416 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1444 = _T_1436 | _T_1437; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  _T_1284 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1346 = ic_miss_buff_data_valid[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1346; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1438 = _T_1419 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1444 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1349 = ic_miss_buff_data_valid[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1349; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1439 = _T_1422 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1425 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1352 = ic_miss_buff_data_valid[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1352; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1440 = _T_1425 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1428 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1355 = ic_miss_buff_data_valid[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1355; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1441 = _T_1428 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1431 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1358 = ic_miss_buff_data_valid[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1358; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1442 = _T_1431 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1434 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 412:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 395:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 395:73]
  wire  _T_1361 = ic_miss_buff_data_valid[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 401:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1361; // @[el2_ifu_mem_ctl.scala 401:88]
  wire  _T_1443 = _T_1434 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1452 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 413:58]
  wire  _T_1453 = bypass_valid_value_check & _T_1452; // @[el2_ifu_mem_ctl.scala 413:56]
  wire  _T_1455 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 413:77]
  wire  _T_1456 = _T_1453 & _T_1455; // @[el2_ifu_mem_ctl.scala 413:75]
  wire  _T_1461 = _T_1453 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 414:75]
  wire  _T_1462 = _T_1456 | _T_1461; // @[el2_ifu_mem_ctl.scala 413:95]
  wire  _T_1464 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 415:56]
  wire  _T_1467 = _T_1464 & _T_1455; // @[el2_ifu_mem_ctl.scala 415:74]
  wire  _T_1468 = _T_1462 | _T_1467; // @[el2_ifu_mem_ctl.scala 414:94]
  wire  _T_1472 = _T_1464 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 416:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 411:70]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1489 = _T_1473 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1490 = _T_1475 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1497 = _T_1489 | _T_1490; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1491 = _T_1477 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1498 = _T_1497 | _T_1491; // @[Mux.scala 27:72]
  wire  _T_1479 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1492 = _T_1479 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1498 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1481 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1493 = _T_1481 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1499 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1483 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1494 = _T_1483 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1500 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1485 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1495 = _T_1485 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1501 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1487 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 416:132]
  wire  _T_1496 = _T_1487 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1502 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1472 & _T_1503; // @[el2_ifu_mem_ctl.scala 416:69]
  wire  _T_1506 = _T_1468 | _T_1505; // @[el2_ifu_mem_ctl.scala 415:94]
  wire [4:0] _GEN_473 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 417:95]
  wire  _T_1509 = _GEN_473 == 5'h1f; // @[el2_ifu_mem_ctl.scala 417:95]
  wire  _T_1510 = bypass_valid_value_check & _T_1509; // @[el2_ifu_mem_ctl.scala 417:56]
  wire  bypass_data_ready_in = _T_1506 | _T_1510; // @[el2_ifu_mem_ctl.scala 416:181]
  wire  _T_1511 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 421:53]
  wire  _T_1512 = _T_1511 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 421:73]
  wire  _T_1514 = _T_1512 & _T_317; // @[el2_ifu_mem_ctl.scala 421:96]
  wire  _T_1516 = _T_1514 & _T_58; // @[el2_ifu_mem_ctl.scala 421:118]
  wire  _T_1518 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 422:73]
  wire  _T_1520 = _T_1518 & _T_317; // @[el2_ifu_mem_ctl.scala 422:96]
  wire  _T_1522 = _T_1520 & _T_58; // @[el2_ifu_mem_ctl.scala 422:118]
  wire  _T_1523 = _T_1516 | _T_1522; // @[el2_ifu_mem_ctl.scala 421:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 424:58]
  wire  _T_1524 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 423:54]
  wire  _T_1525 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 423:76]
  wire  _T_1526 = _T_1524 & _T_1525; // @[el2_ifu_mem_ctl.scala 423:74]
  wire  _T_1528 = _T_1526 & _T_317; // @[el2_ifu_mem_ctl.scala 423:96]
  wire  ic_crit_wd_rdy_new_in = _T_1523 | _T_1528; // @[el2_ifu_mem_ctl.scala 422:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 623:43]
  wire  _T_1249 = ic_crit_wd_rdy | _T_2233; // @[el2_ifu_mem_ctl.scala 369:38]
  wire  _T_1251 = _T_1249 | _T_2249; // @[el2_ifu_mem_ctl.scala 369:64]
  wire  _T_1252 = ~_T_1251; // @[el2_ifu_mem_ctl.scala 369:21]
  wire  _T_1253 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 369:98]
  wire  sel_ic_data = _T_1252 & _T_1253; // @[el2_ifu_mem_ctl.scala 369:96]
  wire  _T_2456 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 468:44]
  wire  _T_1622 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 435:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 407:60]
  wire  _T_1566 = _T_1413 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1416 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1566 | _T_1567; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1419 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1574 | _T_1568; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1422 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1575 | _T_1569; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1425 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1570; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1428 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1571; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1431 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1572; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1434 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1579 | _T_1573; // @[Mux.scala 27:72]
  wire  _T_1605 = _T_2166 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1606 = _T_2169 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1613 = _T_1605 | _T_1606; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_2172 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1614 = _T_1613 | _T_1607; // @[Mux.scala 27:72]
  wire  _T_1608 = _T_2175 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1615 = _T_1614 | _T_1608; // @[Mux.scala 27:72]
  wire  _T_1609 = _T_2178 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1616 = _T_1615 | _T_1609; // @[Mux.scala 27:72]
  wire  _T_1610 = _T_2181 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1617 = _T_1616 | _T_1610; // @[Mux.scala 27:72]
  wire  _T_1611 = _T_2184 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1618 = _T_1617 | _T_1611; // @[Mux.scala 27:72]
  wire  _T_1612 = _T_2187 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1618 | _T_1612; // @[Mux.scala 27:72]
  wire  _T_1623 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 437:70]
  wire  ifu_byp_data_err_new = _T_1622 ? ic_miss_buff_data_error_bypass : _T_1623; // @[el2_ifu_mem_ctl.scala 435:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 380:42]
  wire  _T_2457 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 468:91]
  wire  _T_2458 = ~_T_2457; // @[el2_ifu_mem_ctl.scala 468:60]
  wire  ic_rd_parity_final_err = _T_2456 & _T_2458; // @[el2_ifu_mem_ctl.scala 468:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9606 = _T_4399 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 763:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9608 = _T_4400 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9861 = _T_9606 | _T_9608; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9610 = _T_4401 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9862 = _T_9861 | _T_9610; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9612 = _T_4402 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9863 = _T_9862 | _T_9612; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9614 = _T_4403 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9864 = _T_9863 | _T_9614; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9616 = _T_4404 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9865 = _T_9864 | _T_9616; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9618 = _T_4405 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9866 = _T_9865 | _T_9618; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9620 = _T_4406 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9867 = _T_9866 | _T_9620; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9622 = _T_4407 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9868 = _T_9867 | _T_9622; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9624 = _T_4408 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9869 = _T_9868 | _T_9624; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9626 = _T_4409 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9870 = _T_9869 | _T_9626; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9628 = _T_4410 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9871 = _T_9870 | _T_9628; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9630 = _T_4411 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9872 = _T_9871 | _T_9630; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9632 = _T_4412 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9873 = _T_9872 | _T_9632; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9634 = _T_4413 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9874 = _T_9873 | _T_9634; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9636 = _T_4414 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9875 = _T_9874 | _T_9636; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9638 = _T_4415 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9876 = _T_9875 | _T_9638; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9640 = _T_4416 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9877 = _T_9876 | _T_9640; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9642 = _T_4417 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9878 = _T_9877 | _T_9642; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9644 = _T_4418 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9879 = _T_9878 | _T_9644; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9646 = _T_4419 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9880 = _T_9879 | _T_9646; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9648 = _T_4420 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9881 = _T_9880 | _T_9648; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9650 = _T_4421 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9882 = _T_9881 | _T_9650; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9652 = _T_4422 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9883 = _T_9882 | _T_9652; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9654 = _T_4423 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9884 = _T_9883 | _T_9654; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9656 = _T_4424 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9885 = _T_9884 | _T_9656; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9658 = _T_4425 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9886 = _T_9885 | _T_9658; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9660 = _T_4426 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9887 = _T_9886 | _T_9660; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9662 = _T_4427 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9888 = _T_9887 | _T_9662; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9664 = _T_4428 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9889 = _T_9888 | _T_9664; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9666 = _T_4429 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9890 = _T_9889 | _T_9666; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9668 = _T_4430 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9891 = _T_9890 | _T_9668; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9670 = _T_4431 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9892 = _T_9891 | _T_9670; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9672 = _T_4432 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9893 = _T_9892 | _T_9672; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9674 = _T_4433 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9894 = _T_9893 | _T_9674; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9676 = _T_4434 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9895 = _T_9894 | _T_9676; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9678 = _T_4435 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9896 = _T_9895 | _T_9678; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9680 = _T_4436 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9897 = _T_9896 | _T_9680; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9682 = _T_4437 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9898 = _T_9897 | _T_9682; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9684 = _T_4438 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9899 = _T_9898 | _T_9684; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9686 = _T_4439 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9900 = _T_9899 | _T_9686; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9688 = _T_4440 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9901 = _T_9900 | _T_9688; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9690 = _T_4441 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9902 = _T_9901 | _T_9690; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9692 = _T_4442 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9903 = _T_9902 | _T_9692; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9694 = _T_4443 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9904 = _T_9903 | _T_9694; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9696 = _T_4444 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9905 = _T_9904 | _T_9696; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9698 = _T_4445 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9906 = _T_9905 | _T_9698; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9700 = _T_4446 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9907 = _T_9906 | _T_9700; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9702 = _T_4447 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9908 = _T_9907 | _T_9702; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9704 = _T_4448 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9909 = _T_9908 | _T_9704; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9706 = _T_4449 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9910 = _T_9909 | _T_9706; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9708 = _T_4450 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9911 = _T_9910 | _T_9708; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9710 = _T_4451 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9912 = _T_9911 | _T_9710; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9712 = _T_4452 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9913 = _T_9912 | _T_9712; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9714 = _T_4453 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9914 = _T_9913 | _T_9714; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9716 = _T_4454 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9915 = _T_9914 | _T_9716; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9718 = _T_4455 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9916 = _T_9915 | _T_9718; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9720 = _T_4456 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9917 = _T_9916 | _T_9720; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9722 = _T_4457 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9918 = _T_9917 | _T_9722; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9724 = _T_4458 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9919 = _T_9918 | _T_9724; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9726 = _T_4459 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9920 = _T_9919 | _T_9726; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9728 = _T_4460 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9921 = _T_9920 | _T_9728; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9730 = _T_4461 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9922 = _T_9921 | _T_9730; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9732 = _T_4462 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9923 = _T_9922 | _T_9732; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9734 = _T_4463 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9924 = _T_9923 | _T_9734; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9736 = _T_4464 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9925 = _T_9924 | _T_9736; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9738 = _T_4465 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9926 = _T_9925 | _T_9738; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9740 = _T_4466 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9927 = _T_9926 | _T_9740; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9742 = _T_4467 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9928 = _T_9927 | _T_9742; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9744 = _T_4468 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9929 = _T_9928 | _T_9744; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9746 = _T_4469 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9930 = _T_9929 | _T_9746; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9748 = _T_4470 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9931 = _T_9930 | _T_9748; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9750 = _T_4471 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9932 = _T_9931 | _T_9750; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9752 = _T_4472 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9933 = _T_9932 | _T_9752; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9754 = _T_4473 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9934 = _T_9933 | _T_9754; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9756 = _T_4474 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9935 = _T_9934 | _T_9756; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9758 = _T_4475 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9936 = _T_9935 | _T_9758; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9760 = _T_4476 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9937 = _T_9936 | _T_9760; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9762 = _T_4477 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9938 = _T_9937 | _T_9762; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9764 = _T_4478 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9939 = _T_9938 | _T_9764; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9766 = _T_4479 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9940 = _T_9939 | _T_9766; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9768 = _T_4480 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9941 = _T_9940 | _T_9768; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9770 = _T_4481 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9942 = _T_9941 | _T_9770; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9772 = _T_4482 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9943 = _T_9942 | _T_9772; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9774 = _T_4483 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9944 = _T_9943 | _T_9774; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9776 = _T_4484 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9945 = _T_9944 | _T_9776; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9778 = _T_4485 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9946 = _T_9945 | _T_9778; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9780 = _T_4486 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9947 = _T_9946 | _T_9780; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9782 = _T_4487 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9948 = _T_9947 | _T_9782; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9784 = _T_4488 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9949 = _T_9948 | _T_9784; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9786 = _T_4489 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9950 = _T_9949 | _T_9786; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9788 = _T_4490 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9951 = _T_9950 | _T_9788; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9790 = _T_4491 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9952 = _T_9951 | _T_9790; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9792 = _T_4492 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9953 = _T_9952 | _T_9792; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9794 = _T_4493 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9954 = _T_9953 | _T_9794; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9796 = _T_4494 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9955 = _T_9954 | _T_9796; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9798 = _T_4495 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9956 = _T_9955 | _T_9798; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9800 = _T_4496 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9957 = _T_9956 | _T_9800; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9802 = _T_4497 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9958 = _T_9957 | _T_9802; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9804 = _T_4498 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9959 = _T_9958 | _T_9804; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9806 = _T_4499 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9960 = _T_9959 | _T_9806; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9808 = _T_4500 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9961 = _T_9960 | _T_9808; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9810 = _T_4501 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9962 = _T_9961 | _T_9810; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9812 = _T_4502 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9963 = _T_9962 | _T_9812; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9814 = _T_4503 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9964 = _T_9963 | _T_9814; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9816 = _T_4504 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9965 = _T_9964 | _T_9816; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9818 = _T_4505 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9966 = _T_9965 | _T_9818; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9820 = _T_4506 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9967 = _T_9966 | _T_9820; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9822 = _T_4507 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9968 = _T_9967 | _T_9822; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9824 = _T_4508 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9969 = _T_9968 | _T_9824; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9826 = _T_4509 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9970 = _T_9969 | _T_9826; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9828 = _T_4510 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9971 = _T_9970 | _T_9828; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9830 = _T_4511 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9972 = _T_9971 | _T_9830; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9832 = _T_4512 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9973 = _T_9972 | _T_9832; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9834 = _T_4513 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9974 = _T_9973 | _T_9834; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9836 = _T_4514 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9975 = _T_9974 | _T_9836; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9838 = _T_4515 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9976 = _T_9975 | _T_9838; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9840 = _T_4516 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9977 = _T_9976 | _T_9840; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9842 = _T_4517 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9978 = _T_9977 | _T_9842; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9844 = _T_4518 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9979 = _T_9978 | _T_9844; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9846 = _T_4519 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9980 = _T_9979 | _T_9846; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9848 = _T_4520 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9981 = _T_9980 | _T_9848; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9850 = _T_4521 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9982 = _T_9981 | _T_9850; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9852 = _T_4522 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9983 = _T_9982 | _T_9852; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9854 = _T_4523 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9984 = _T_9983 | _T_9854; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9856 = _T_4524 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9985 = _T_9984 | _T_9856; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9858 = _T_4525 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9986 = _T_9985 | _T_9858; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9860 = _T_4526 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9987 = _T_9986 | _T_9860; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9223 = _T_4399 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 763:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9225 = _T_4400 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9478 = _T_9223 | _T_9225; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9227 = _T_4401 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9479 = _T_9478 | _T_9227; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9229 = _T_4402 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9480 = _T_9479 | _T_9229; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9231 = _T_4403 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9481 = _T_9480 | _T_9231; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9233 = _T_4404 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9482 = _T_9481 | _T_9233; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9235 = _T_4405 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9483 = _T_9482 | _T_9235; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9237 = _T_4406 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9484 = _T_9483 | _T_9237; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9239 = _T_4407 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9485 = _T_9484 | _T_9239; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9241 = _T_4408 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9486 = _T_9485 | _T_9241; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9243 = _T_4409 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9487 = _T_9486 | _T_9243; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9245 = _T_4410 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9488 = _T_9487 | _T_9245; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9247 = _T_4411 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9489 = _T_9488 | _T_9247; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9249 = _T_4412 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9490 = _T_9489 | _T_9249; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9251 = _T_4413 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9491 = _T_9490 | _T_9251; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9253 = _T_4414 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9492 = _T_9491 | _T_9253; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9255 = _T_4415 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9493 = _T_9492 | _T_9255; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9257 = _T_4416 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9494 = _T_9493 | _T_9257; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9259 = _T_4417 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9495 = _T_9494 | _T_9259; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9261 = _T_4418 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9496 = _T_9495 | _T_9261; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9263 = _T_4419 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9497 = _T_9496 | _T_9263; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9265 = _T_4420 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9498 = _T_9497 | _T_9265; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9267 = _T_4421 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9499 = _T_9498 | _T_9267; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9269 = _T_4422 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9500 = _T_9499 | _T_9269; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9271 = _T_4423 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9501 = _T_9500 | _T_9271; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9273 = _T_4424 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9502 = _T_9501 | _T_9273; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9275 = _T_4425 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9503 = _T_9502 | _T_9275; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9277 = _T_4426 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9504 = _T_9503 | _T_9277; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9279 = _T_4427 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9505 = _T_9504 | _T_9279; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9281 = _T_4428 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9506 = _T_9505 | _T_9281; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9283 = _T_4429 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9507 = _T_9506 | _T_9283; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9285 = _T_4430 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9508 = _T_9507 | _T_9285; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9287 = _T_4431 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9509 = _T_9508 | _T_9287; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9289 = _T_4432 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9510 = _T_9509 | _T_9289; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9291 = _T_4433 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9511 = _T_9510 | _T_9291; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9293 = _T_4434 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9512 = _T_9511 | _T_9293; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9295 = _T_4435 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9513 = _T_9512 | _T_9295; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9297 = _T_4436 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9514 = _T_9513 | _T_9297; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9299 = _T_4437 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9515 = _T_9514 | _T_9299; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9301 = _T_4438 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9516 = _T_9515 | _T_9301; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9303 = _T_4439 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9517 = _T_9516 | _T_9303; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9305 = _T_4440 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9518 = _T_9517 | _T_9305; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9307 = _T_4441 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9519 = _T_9518 | _T_9307; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9309 = _T_4442 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9520 = _T_9519 | _T_9309; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9311 = _T_4443 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9521 = _T_9520 | _T_9311; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9313 = _T_4444 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9522 = _T_9521 | _T_9313; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9315 = _T_4445 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9523 = _T_9522 | _T_9315; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9317 = _T_4446 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9524 = _T_9523 | _T_9317; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9319 = _T_4447 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9525 = _T_9524 | _T_9319; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9321 = _T_4448 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9526 = _T_9525 | _T_9321; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9323 = _T_4449 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9527 = _T_9526 | _T_9323; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9325 = _T_4450 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9528 = _T_9527 | _T_9325; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9327 = _T_4451 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9529 = _T_9528 | _T_9327; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9329 = _T_4452 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9530 = _T_9529 | _T_9329; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9331 = _T_4453 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9531 = _T_9530 | _T_9331; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9333 = _T_4454 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9532 = _T_9531 | _T_9333; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9335 = _T_4455 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9533 = _T_9532 | _T_9335; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9337 = _T_4456 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9534 = _T_9533 | _T_9337; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9339 = _T_4457 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9535 = _T_9534 | _T_9339; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9341 = _T_4458 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9536 = _T_9535 | _T_9341; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9343 = _T_4459 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9537 = _T_9536 | _T_9343; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9345 = _T_4460 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9538 = _T_9537 | _T_9345; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9347 = _T_4461 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9539 = _T_9538 | _T_9347; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9349 = _T_4462 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9540 = _T_9539 | _T_9349; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9351 = _T_4463 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9541 = _T_9540 | _T_9351; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9353 = _T_4464 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9542 = _T_9541 | _T_9353; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9355 = _T_4465 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9543 = _T_9542 | _T_9355; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9357 = _T_4466 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9544 = _T_9543 | _T_9357; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9359 = _T_4467 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9545 = _T_9544 | _T_9359; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9361 = _T_4468 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9546 = _T_9545 | _T_9361; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9363 = _T_4469 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9547 = _T_9546 | _T_9363; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9365 = _T_4470 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9548 = _T_9547 | _T_9365; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9367 = _T_4471 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9549 = _T_9548 | _T_9367; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9369 = _T_4472 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9550 = _T_9549 | _T_9369; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9371 = _T_4473 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9551 = _T_9550 | _T_9371; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9373 = _T_4474 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9552 = _T_9551 | _T_9373; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9375 = _T_4475 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9553 = _T_9552 | _T_9375; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9377 = _T_4476 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9554 = _T_9553 | _T_9377; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9379 = _T_4477 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9555 = _T_9554 | _T_9379; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9381 = _T_4478 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9556 = _T_9555 | _T_9381; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9383 = _T_4479 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9557 = _T_9556 | _T_9383; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9385 = _T_4480 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9558 = _T_9557 | _T_9385; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9387 = _T_4481 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9559 = _T_9558 | _T_9387; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9389 = _T_4482 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9560 = _T_9559 | _T_9389; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9391 = _T_4483 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9561 = _T_9560 | _T_9391; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9393 = _T_4484 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9562 = _T_9561 | _T_9393; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9395 = _T_4485 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9563 = _T_9562 | _T_9395; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9397 = _T_4486 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9564 = _T_9563 | _T_9397; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9399 = _T_4487 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9565 = _T_9564 | _T_9399; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9401 = _T_4488 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9566 = _T_9565 | _T_9401; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9403 = _T_4489 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9567 = _T_9566 | _T_9403; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9405 = _T_4490 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9568 = _T_9567 | _T_9405; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9407 = _T_4491 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9569 = _T_9568 | _T_9407; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9409 = _T_4492 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9570 = _T_9569 | _T_9409; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9411 = _T_4493 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9571 = _T_9570 | _T_9411; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9413 = _T_4494 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9572 = _T_9571 | _T_9413; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9415 = _T_4495 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9573 = _T_9572 | _T_9415; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9417 = _T_4496 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9574 = _T_9573 | _T_9417; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9419 = _T_4497 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9575 = _T_9574 | _T_9419; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9421 = _T_4498 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9576 = _T_9575 | _T_9421; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9423 = _T_4499 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9577 = _T_9576 | _T_9423; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9425 = _T_4500 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9578 = _T_9577 | _T_9425; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9427 = _T_4501 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9579 = _T_9578 | _T_9427; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9429 = _T_4502 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9580 = _T_9579 | _T_9429; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9431 = _T_4503 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9581 = _T_9580 | _T_9431; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9433 = _T_4504 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9582 = _T_9581 | _T_9433; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9435 = _T_4505 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9583 = _T_9582 | _T_9435; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9437 = _T_4506 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9584 = _T_9583 | _T_9437; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9439 = _T_4507 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9585 = _T_9584 | _T_9439; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9441 = _T_4508 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9586 = _T_9585 | _T_9441; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9443 = _T_4509 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9587 = _T_9586 | _T_9443; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9445 = _T_4510 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9588 = _T_9587 | _T_9445; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9447 = _T_4511 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9589 = _T_9588 | _T_9447; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9449 = _T_4512 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9590 = _T_9589 | _T_9449; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9451 = _T_4513 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9591 = _T_9590 | _T_9451; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9453 = _T_4514 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9592 = _T_9591 | _T_9453; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9455 = _T_4515 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9593 = _T_9592 | _T_9455; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9457 = _T_4516 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9594 = _T_9593 | _T_9457; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9459 = _T_4517 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9595 = _T_9594 | _T_9459; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9461 = _T_4518 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9596 = _T_9595 | _T_9461; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9463 = _T_4519 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9597 = _T_9596 | _T_9463; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9465 = _T_4520 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9598 = _T_9597 | _T_9465; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9467 = _T_4521 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9599 = _T_9598 | _T_9467; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9469 = _T_4522 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9600 = _T_9599 | _T_9469; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9471 = _T_4523 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9601 = _T_9600 | _T_9471; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9473 = _T_4524 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9602 = _T_9601 | _T_9473; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9475 = _T_4525 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9603 = _T_9602 | _T_9475; // @[el2_ifu_mem_ctl.scala 763:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9477 = _T_4526 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 763:10]
  wire  _T_9604 = _T_9603 | _T_9477; // @[el2_ifu_mem_ctl.scala 763:91]
  wire [1:0] ic_tag_valid_unq = {_T_9987,_T_9604}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 837:54]
  wire [1:0] _T_10027 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10028 = ic_debug_way_ff & _T_10027; // @[el2_ifu_mem_ctl.scala 818:67]
  wire [1:0] _T_10029 = ic_tag_valid_unq & _T_10028; // @[el2_ifu_mem_ctl.scala 818:48]
  wire  ic_debug_tag_val_rd_out = |_T_10029; // @[el2_ifu_mem_ctl.scala 818:115]
  wire [65:0] _T_1208 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1209; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2591; // @[el2_ifu_mem_ctl.scala 363:80]
  wire  _T_1247 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 368:98]
  wire  sel_byp_data = _T_1251 & _T_1247; // @[el2_ifu_mem_ctl.scala 368:96]
  wire [63:0] _T_1258 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1259 = _T_1258 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 375:69]
  wire [63:0] _T_1261 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2113 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 443:31]
  wire  _T_1626 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 439:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1627 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1675 = _T_1627 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1630 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1676 = _T_1630 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1675 | _T_1676; // @[Mux.scala 27:72]
  wire  _T_1633 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1677 = _T_1633 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1692 = _T_1691 | _T_1677; // @[Mux.scala 27:72]
  wire  _T_1636 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1678 = _T_1636 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1692 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1639 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1679 = _T_1639 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire  _T_1642 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1680 = _T_1642 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1695 = _T_1694 | _T_1680; // @[Mux.scala 27:72]
  wire  _T_1645 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1681 = _T_1645 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1696 = _T_1695 | _T_1681; // @[Mux.scala 27:72]
  wire  _T_1648 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1682 = _T_1648 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1697 = _T_1696 | _T_1682; // @[Mux.scala 27:72]
  wire  _T_1651 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1683 = _T_1651 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1698 = _T_1697 | _T_1683; // @[Mux.scala 27:72]
  wire  _T_1654 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1684 = _T_1654 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1699 = _T_1698 | _T_1684; // @[Mux.scala 27:72]
  wire  _T_1657 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1685 = _T_1657 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1700 = _T_1699 | _T_1685; // @[Mux.scala 27:72]
  wire  _T_1660 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1686 = _T_1660 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1701 = _T_1700 | _T_1686; // @[Mux.scala 27:72]
  wire  _T_1663 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1687 = _T_1663 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1702 = _T_1701 | _T_1687; // @[Mux.scala 27:72]
  wire  _T_1666 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1688 = _T_1666 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1703 = _T_1702 | _T_1688; // @[Mux.scala 27:72]
  wire  _T_1669 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1689 = _T_1669 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1704 = _T_1703 | _T_1689; // @[Mux.scala 27:72]
  wire  _T_1672 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 440:73]
  wire [15:0] _T_1690 = _T_1672 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1705 = _T_1704 | _T_1690; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1707 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1755 = _T_1707 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1710 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1756 = _T_1710 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1755 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1713 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1757 = _T_1713 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1772 = _T_1771 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1716 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1758 = _T_1716 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1772 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1719 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1759 = _T_1719 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1722 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1760 = _T_1722 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1775 = _T_1774 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1725 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1761 = _T_1725 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1776 = _T_1775 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1728 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1762 = _T_1728 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1777 = _T_1776 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1731 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1763 = _T_1731 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1778 = _T_1777 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1734 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1764 = _T_1734 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1779 = _T_1778 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1737 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1765 = _T_1737 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1780 = _T_1779 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1740 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1766 = _T_1740 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1781 = _T_1780 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1743 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1767 = _T_1743 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1782 = _T_1781 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1746 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1768 = _T_1746 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1783 = _T_1782 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1749 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1769 = _T_1749 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1784 = _T_1783 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1752 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 440:179]
  wire [31:0] _T_1770 = _T_1752 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1785 = _T_1784 | _T_1770; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1787 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1835 = _T_1787 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1790 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1836 = _T_1790 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1835 | _T_1836; // @[Mux.scala 27:72]
  wire  _T_1793 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1837 = _T_1793 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1852 = _T_1851 | _T_1837; // @[Mux.scala 27:72]
  wire  _T_1796 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1838 = _T_1796 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1852 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1799 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1839 = _T_1799 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire  _T_1802 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1840 = _T_1802 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1855 = _T_1854 | _T_1840; // @[Mux.scala 27:72]
  wire  _T_1805 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1841 = _T_1805 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1856 = _T_1855 | _T_1841; // @[Mux.scala 27:72]
  wire  _T_1808 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1842 = _T_1808 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1857 = _T_1856 | _T_1842; // @[Mux.scala 27:72]
  wire  _T_1811 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1843 = _T_1811 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1858 = _T_1857 | _T_1843; // @[Mux.scala 27:72]
  wire  _T_1814 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1844 = _T_1814 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1859 = _T_1858 | _T_1844; // @[Mux.scala 27:72]
  wire  _T_1817 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1845 = _T_1817 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1860 = _T_1859 | _T_1845; // @[Mux.scala 27:72]
  wire  _T_1820 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1846 = _T_1820 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1861 = _T_1860 | _T_1846; // @[Mux.scala 27:72]
  wire  _T_1823 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1847 = _T_1823 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1862 = _T_1861 | _T_1847; // @[Mux.scala 27:72]
  wire  _T_1826 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1848 = _T_1826 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1863 = _T_1862 | _T_1848; // @[Mux.scala 27:72]
  wire  _T_1829 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1849 = _T_1829 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1864 = _T_1863 | _T_1849; // @[Mux.scala 27:72]
  wire  _T_1832 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 440:285]
  wire [31:0] _T_1850 = _T_1832 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1865 = _T_1864 | _T_1850; // @[Mux.scala 27:72]
  wire [79:0] _T_1868 = {_T_1705,_T_1785,_T_1865}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1869 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1917 = _T_1869 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1918 = _T_1872 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1917 | _T_1918; // @[Mux.scala 27:72]
  wire  _T_1875 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1919 = _T_1875 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1934 = _T_1933 | _T_1919; // @[Mux.scala 27:72]
  wire  _T_1878 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1920 = _T_1878 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1934 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1881 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1921 = _T_1881 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire  _T_1884 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1922 = _T_1884 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1937 = _T_1936 | _T_1922; // @[Mux.scala 27:72]
  wire  _T_1887 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1923 = _T_1887 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1938 = _T_1937 | _T_1923; // @[Mux.scala 27:72]
  wire  _T_1890 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1924 = _T_1890 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1939 = _T_1938 | _T_1924; // @[Mux.scala 27:72]
  wire  _T_1893 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1925 = _T_1893 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1940 = _T_1939 | _T_1925; // @[Mux.scala 27:72]
  wire  _T_1896 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1926 = _T_1896 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1941 = _T_1940 | _T_1926; // @[Mux.scala 27:72]
  wire  _T_1899 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1927 = _T_1899 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1942 = _T_1941 | _T_1927; // @[Mux.scala 27:72]
  wire  _T_1902 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1928 = _T_1902 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1943 = _T_1942 | _T_1928; // @[Mux.scala 27:72]
  wire  _T_1905 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1929 = _T_1905 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1944 = _T_1943 | _T_1929; // @[Mux.scala 27:72]
  wire  _T_1908 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1930 = _T_1908 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1945 = _T_1944 | _T_1930; // @[Mux.scala 27:72]
  wire  _T_1911 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1931 = _T_1911 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1946 = _T_1945 | _T_1931; // @[Mux.scala 27:72]
  wire  _T_1914 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1932 = _T_1914 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1947 = _T_1946 | _T_1932; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1627 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1630 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_1997 | _T_1998; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1633 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_2013 | _T_1999; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1636 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_2014 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1639 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1642 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2017 = _T_2016 | _T_2002; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_1645 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2018 = _T_2017 | _T_2003; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_1648 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2019 = _T_2018 | _T_2004; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_1651 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2020 = _T_2019 | _T_2005; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_1654 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2021 = _T_2020 | _T_2006; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_1657 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2022 = _T_2021 | _T_2007; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_1660 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2023 = _T_2022 | _T_2008; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_1663 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2024 = _T_2023 | _T_2009; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_1666 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2025 = _T_2024 | _T_2010; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_1669 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2026 = _T_2025 | _T_2011; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_1672 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2027 = _T_2026 | _T_2012; // @[Mux.scala 27:72]
  wire [79:0] _T_2110 = {_T_1947,_T_2027,_T_1785}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1626 ? _T_1868 : _T_2110; // @[el2_ifu_mem_ctl.scala 439:37]
  wire [79:0] _T_2115 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2113 ? ic_byp_data_only_pre_new : _T_2115; // @[el2_ifu_mem_ctl.scala 443:30]
  wire [79:0] _GEN_474 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 375:114]
  wire [79:0] _T_1262 = _GEN_474 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 375:114]
  wire [79:0] _GEN_475 = {{16'd0}, _T_1259}; // @[el2_ifu_mem_ctl.scala 375:88]
  wire [79:0] ic_premux_data_temp = _GEN_475 | _T_1262; // @[el2_ifu_mem_ctl.scala 375:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 382:38]
  wire [1:0] _T_1271 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 386:8]
  wire  _T_1273 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 388:45]
  wire  _T_1275 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 388:80]
  wire  _T_1276 = ~_T_1275; // @[el2_ifu_mem_ctl.scala 388:71]
  wire  _T_1277 = _T_1273 & _T_1276; // @[el2_ifu_mem_ctl.scala 388:69]
  wire  _T_1278 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 388:131]
  wire  _T_1279 = _T_1277 & _T_1278; // @[el2_ifu_mem_ctl.scala 388:114]
  wire [7:0] _T_1368 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1373 = ic_miss_buff_data_error[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  _T_2659 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 619:47]
  wire  _T_2660 = _T_2659 & _T_13; // @[el2_ifu_mem_ctl.scala 619:50]
  wire  bus_ifu_wr_data_error = _T_2660 & miss_pending; // @[el2_ifu_mem_ctl.scala 619:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1373; // @[el2_ifu_mem_ctl.scala 405:72]
  wire  _T_1377 = ic_miss_buff_data_error[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1377; // @[el2_ifu_mem_ctl.scala 405:72]
  wire  _T_1381 = ic_miss_buff_data_error[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1381; // @[el2_ifu_mem_ctl.scala 405:72]
  wire  _T_1385 = ic_miss_buff_data_error[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1385; // @[el2_ifu_mem_ctl.scala 405:72]
  wire  _T_1389 = ic_miss_buff_data_error[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1389; // @[el2_ifu_mem_ctl.scala 405:72]
  wire  _T_1393 = ic_miss_buff_data_error[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1393; // @[el2_ifu_mem_ctl.scala 405:72]
  wire  _T_1397 = ic_miss_buff_data_error[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1397; // @[el2_ifu_mem_ctl.scala 405:72]
  wire  _T_1401 = ic_miss_buff_data_error[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1401; // @[el2_ifu_mem_ctl.scala 405:72]
  wire [7:0] _T_1408 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2465 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2473 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 488:65]
  wire  _T_2474 = _T_2473 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 488:88]
  wire  _T_2476 = _T_2474 & _T_2587; // @[el2_ifu_mem_ctl.scala 488:112]
  wire  _T_2477 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2478 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 493:50]
  wire  _T_2480 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2486 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2488 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_2486 | _T_2488; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2480 ? _T_2478 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_2477 ? _T_2478 : _GEN_41; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2465 ? _T_2476 : _GEN_43; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2465 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2479 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 494:56]
  wire  _GEN_44 = _T_2477 & _T_2479; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2465 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 479:58]
  wire  _T_2462 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 478:49]
  wire  _T_2467 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 487:87]
  wire  _T_2481 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 497:54]
  wire  _T_2482 = _T_2481 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 497:84]
  wire  _T_2491 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 518:66]
  wire  _T_2492 = io_dec_tlu_flush_err_wb & _T_2491; // @[el2_ifu_mem_ctl.scala 518:52]
  wire  _T_2494 = _T_2492 & _T_2587; // @[el2_ifu_mem_ctl.scala 518:81]
  wire  _T_2496 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 521:59]
  wire  _T_2497 = _T_2496 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 521:86]
  wire  _T_2511 = _T_2496 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 524:81]
  wire  _T_2512 = _T_2511 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 524:103]
  wire  _T_2513 = _T_2512 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 524:126]
  wire  _T_2533 = _T_2511 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 531:103]
  wire  _T_2540 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 536:62]
  wire  _T_2541 = io_dec_tlu_flush_lower_wb & _T_2540; // @[el2_ifu_mem_ctl.scala 536:60]
  wire  _T_2542 = _T_2541 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 536:88]
  wire  _T_2543 = _T_2542 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 536:115]
  wire  _GEN_51 = _T_2539 & _T_2497; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_2522 ? _T_2533 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_2522 | _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2495 ? _T_2513 : _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_2495 | _GEN_56; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2490 ? _T_2494 : _GEN_58; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2555 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 553:64]
  wire  _T_2557 = _T_2555 & _T_2587; // @[el2_ifu_mem_ctl.scala 553:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2559 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 553:133]
  wire  _T_2560 = _T_2559 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 553:164]
  wire  _T_2561 = _T_2560 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 553:184]
  wire  _T_2562 = _T_2561 & miss_pending; // @[el2_ifu_mem_ctl.scala 553:204]
  wire  _T_2563 = ~_T_2562; // @[el2_ifu_mem_ctl.scala 553:112]
  wire  ifc_bus_ic_req_ff_in = _T_2557 & _T_2563; // @[el2_ifu_mem_ctl.scala 553:110]
  wire  _T_2564 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 554:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 585:45]
  wire  _T_2581 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 588:35]
  wire  _T_2582 = _T_2581 & miss_pending; // @[el2_ifu_mem_ctl.scala 588:53]
  wire  bus_cmd_sent = _T_2582 & _T_2587; // @[el2_ifu_mem_ctl.scala 588:68]
  wire [2:0] _T_2572 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2574 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2576 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 586:51]
  wire  _T_2602 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 596:73]
  wire  _T_2603 = _T_2588 & _T_2602; // @[el2_ifu_mem_ctl.scala 596:71]
  wire  _T_2605 = last_data_recieved_ff & _T_1339; // @[el2_ifu_mem_ctl.scala 596:114]
  wire  last_data_recieved_in = _T_2603 | _T_2605; // @[el2_ifu_mem_ctl.scala 596:89]
  wire [2:0] _T_2611 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 601:45]
  wire  _T_2614 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 602:81]
  wire  _T_2615 = _T_2614 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 602:97]
  wire  _T_2617 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 604:48]
  wire  _T_2618 = _T_2617 & miss_pending; // @[el2_ifu_mem_ctl.scala 604:68]
  wire  bus_inc_cmd_beat_cnt = _T_2618 & _T_2587; // @[el2_ifu_mem_ctl.scala 604:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 606:57]
  wire  _T_2622 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 607:31]
  wire  _T_2623 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 607:71]
  wire  _T_2624 = _T_2623 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 607:87]
  wire  _T_2625 = ~_T_2624; // @[el2_ifu_mem_ctl.scala 607:55]
  wire  bus_hold_cmd_beat_cnt = _T_2622 & _T_2625; // @[el2_ifu_mem_ctl.scala 607:53]
  wire  _T_2626 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 608:46]
  wire  bus_cmd_beat_en = _T_2626 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 608:62]
  wire [2:0] _T_2629 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 610:46]
  wire [2:0] _T_2631 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2632 = bus_inc_cmd_beat_cnt ? _T_2629 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2633 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2635 = _T_2631 | _T_2632; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2635 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2639 = _T_2615 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 611:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 622:62]
  wire  _T_2667 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 627:50]
  wire  _T_2668 = io_ifc_dma_access_ok & _T_2667; // @[el2_ifu_mem_ctl.scala 627:47]
  wire  _T_2669 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 627:70]
  wire  ifc_dma_access_ok_d = _T_2668 & _T_2669; // @[el2_ifu_mem_ctl.scala 627:68]
  wire  _T_2673 = _T_2668 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 628:72]
  wire  _T_2674 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 628:111]
  wire  _T_2675 = _T_2673 & _T_2674; // @[el2_ifu_mem_ctl.scala 628:97]
  wire  ifc_dma_access_q_ok = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 628:127]
  wire  _T_2678 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 631:40]
  wire  _T_2679 = _T_2678 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 631:58]
  wire  _T_2682 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 632:60]
  wire  _T_2683 = _T_2678 & _T_2682; // @[el2_ifu_mem_ctl.scala 632:58]
  wire  _T_2684 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 632:104]
  wire [2:0] _T_2689 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [13:0] dma_mem_ecc = {m2_io_ecc_out,m1_io_ecc_out}; // @[Cat.scala 29:58]
  wire  _T_2694 = ~_T_2678; // @[el2_ifu_mem_ctl.scala 641:45]
  wire  _T_2695 = iccm_correct_ecc & _T_2694; // @[el2_ifu_mem_ctl.scala 641:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_2696 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_2703 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 655:53]
  wire  _T_3035 = _T_2947[5:0] == 6'h27; // @[el2_lib.scala 340:41]
  wire  _T_3033 = _T_2947[5:0] == 6'h26; // @[el2_lib.scala 340:41]
  wire  _T_3031 = _T_2947[5:0] == 6'h25; // @[el2_lib.scala 340:41]
  wire  _T_3029 = _T_2947[5:0] == 6'h24; // @[el2_lib.scala 340:41]
  wire  _T_3027 = _T_2947[5:0] == 6'h23; // @[el2_lib.scala 340:41]
  wire  _T_3025 = _T_2947[5:0] == 6'h22; // @[el2_lib.scala 340:41]
  wire  _T_3023 = _T_2947[5:0] == 6'h21; // @[el2_lib.scala 340:41]
  wire  _T_3021 = _T_2947[5:0] == 6'h20; // @[el2_lib.scala 340:41]
  wire  _T_3019 = _T_2947[5:0] == 6'h1f; // @[el2_lib.scala 340:41]
  wire  _T_3017 = _T_2947[5:0] == 6'h1e; // @[el2_lib.scala 340:41]
  wire [9:0] _T_3093 = {_T_3035,_T_3033,_T_3031,_T_3029,_T_3027,_T_3025,_T_3023,_T_3021,_T_3019,_T_3017}; // @[el2_lib.scala 343:69]
  wire  _T_3015 = _T_2947[5:0] == 6'h1d; // @[el2_lib.scala 340:41]
  wire  _T_3013 = _T_2947[5:0] == 6'h1c; // @[el2_lib.scala 340:41]
  wire  _T_3011 = _T_2947[5:0] == 6'h1b; // @[el2_lib.scala 340:41]
  wire  _T_3009 = _T_2947[5:0] == 6'h1a; // @[el2_lib.scala 340:41]
  wire  _T_3007 = _T_2947[5:0] == 6'h19; // @[el2_lib.scala 340:41]
  wire  _T_3005 = _T_2947[5:0] == 6'h18; // @[el2_lib.scala 340:41]
  wire  _T_3003 = _T_2947[5:0] == 6'h17; // @[el2_lib.scala 340:41]
  wire  _T_3001 = _T_2947[5:0] == 6'h16; // @[el2_lib.scala 340:41]
  wire  _T_2999 = _T_2947[5:0] == 6'h15; // @[el2_lib.scala 340:41]
  wire  _T_2997 = _T_2947[5:0] == 6'h14; // @[el2_lib.scala 340:41]
  wire [9:0] _T_3084 = {_T_3015,_T_3013,_T_3011,_T_3009,_T_3007,_T_3005,_T_3003,_T_3001,_T_2999,_T_2997}; // @[el2_lib.scala 343:69]
  wire  _T_2995 = _T_2947[5:0] == 6'h13; // @[el2_lib.scala 340:41]
  wire  _T_2993 = _T_2947[5:0] == 6'h12; // @[el2_lib.scala 340:41]
  wire  _T_2991 = _T_2947[5:0] == 6'h11; // @[el2_lib.scala 340:41]
  wire  _T_2989 = _T_2947[5:0] == 6'h10; // @[el2_lib.scala 340:41]
  wire  _T_2987 = _T_2947[5:0] == 6'hf; // @[el2_lib.scala 340:41]
  wire  _T_2985 = _T_2947[5:0] == 6'he; // @[el2_lib.scala 340:41]
  wire  _T_2983 = _T_2947[5:0] == 6'hd; // @[el2_lib.scala 340:41]
  wire  _T_2981 = _T_2947[5:0] == 6'hc; // @[el2_lib.scala 340:41]
  wire  _T_2979 = _T_2947[5:0] == 6'hb; // @[el2_lib.scala 340:41]
  wire  _T_2977 = _T_2947[5:0] == 6'ha; // @[el2_lib.scala 340:41]
  wire [9:0] _T_3074 = {_T_2995,_T_2993,_T_2991,_T_2989,_T_2987,_T_2985,_T_2983,_T_2981,_T_2979,_T_2977}; // @[el2_lib.scala 343:69]
  wire  _T_2975 = _T_2947[5:0] == 6'h9; // @[el2_lib.scala 340:41]
  wire  _T_2973 = _T_2947[5:0] == 6'h8; // @[el2_lib.scala 340:41]
  wire  _T_2971 = _T_2947[5:0] == 6'h7; // @[el2_lib.scala 340:41]
  wire  _T_2969 = _T_2947[5:0] == 6'h6; // @[el2_lib.scala 340:41]
  wire  _T_2967 = _T_2947[5:0] == 6'h5; // @[el2_lib.scala 340:41]
  wire  _T_2965 = _T_2947[5:0] == 6'h4; // @[el2_lib.scala 340:41]
  wire  _T_2963 = _T_2947[5:0] == 6'h3; // @[el2_lib.scala 340:41]
  wire  _T_2961 = _T_2947[5:0] == 6'h2; // @[el2_lib.scala 340:41]
  wire  _T_2959 = _T_2947[5:0] == 6'h1; // @[el2_lib.scala 340:41]
  wire [18:0] _T_3075 = {_T_3074,_T_2975,_T_2973,_T_2971,_T_2969,_T_2967,_T_2965,_T_2963,_T_2961,_T_2959}; // @[el2_lib.scala 343:69]
  wire [38:0] _T_3095 = {_T_3093,_T_3084,_T_3075}; // @[el2_lib.scala 343:69]
  wire [7:0] _T_3050 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3056 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3050}; // @[Cat.scala 29:58]
  wire [38:0] _T_3096 = _T_3095 ^ _T_3056; // @[el2_lib.scala 343:76]
  wire [38:0] _T_3097 = _T_2951 ? _T_3096 : _T_3056; // @[el2_lib.scala 343:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3097[37:32],_T_3097[30:16],_T_3097[14:8],_T_3097[6:4],_T_3097[2]}; // @[Cat.scala 29:58]
  wire  _T_3420 = _T_3332[5:0] == 6'h27; // @[el2_lib.scala 340:41]
  wire  _T_3418 = _T_3332[5:0] == 6'h26; // @[el2_lib.scala 340:41]
  wire  _T_3416 = _T_3332[5:0] == 6'h25; // @[el2_lib.scala 340:41]
  wire  _T_3414 = _T_3332[5:0] == 6'h24; // @[el2_lib.scala 340:41]
  wire  _T_3412 = _T_3332[5:0] == 6'h23; // @[el2_lib.scala 340:41]
  wire  _T_3410 = _T_3332[5:0] == 6'h22; // @[el2_lib.scala 340:41]
  wire  _T_3408 = _T_3332[5:0] == 6'h21; // @[el2_lib.scala 340:41]
  wire  _T_3406 = _T_3332[5:0] == 6'h20; // @[el2_lib.scala 340:41]
  wire  _T_3404 = _T_3332[5:0] == 6'h1f; // @[el2_lib.scala 340:41]
  wire  _T_3402 = _T_3332[5:0] == 6'h1e; // @[el2_lib.scala 340:41]
  wire [9:0] _T_3478 = {_T_3420,_T_3418,_T_3416,_T_3414,_T_3412,_T_3410,_T_3408,_T_3406,_T_3404,_T_3402}; // @[el2_lib.scala 343:69]
  wire  _T_3400 = _T_3332[5:0] == 6'h1d; // @[el2_lib.scala 340:41]
  wire  _T_3398 = _T_3332[5:0] == 6'h1c; // @[el2_lib.scala 340:41]
  wire  _T_3396 = _T_3332[5:0] == 6'h1b; // @[el2_lib.scala 340:41]
  wire  _T_3394 = _T_3332[5:0] == 6'h1a; // @[el2_lib.scala 340:41]
  wire  _T_3392 = _T_3332[5:0] == 6'h19; // @[el2_lib.scala 340:41]
  wire  _T_3390 = _T_3332[5:0] == 6'h18; // @[el2_lib.scala 340:41]
  wire  _T_3388 = _T_3332[5:0] == 6'h17; // @[el2_lib.scala 340:41]
  wire  _T_3386 = _T_3332[5:0] == 6'h16; // @[el2_lib.scala 340:41]
  wire  _T_3384 = _T_3332[5:0] == 6'h15; // @[el2_lib.scala 340:41]
  wire  _T_3382 = _T_3332[5:0] == 6'h14; // @[el2_lib.scala 340:41]
  wire [9:0] _T_3469 = {_T_3400,_T_3398,_T_3396,_T_3394,_T_3392,_T_3390,_T_3388,_T_3386,_T_3384,_T_3382}; // @[el2_lib.scala 343:69]
  wire  _T_3380 = _T_3332[5:0] == 6'h13; // @[el2_lib.scala 340:41]
  wire  _T_3378 = _T_3332[5:0] == 6'h12; // @[el2_lib.scala 340:41]
  wire  _T_3376 = _T_3332[5:0] == 6'h11; // @[el2_lib.scala 340:41]
  wire  _T_3374 = _T_3332[5:0] == 6'h10; // @[el2_lib.scala 340:41]
  wire  _T_3372 = _T_3332[5:0] == 6'hf; // @[el2_lib.scala 340:41]
  wire  _T_3370 = _T_3332[5:0] == 6'he; // @[el2_lib.scala 340:41]
  wire  _T_3368 = _T_3332[5:0] == 6'hd; // @[el2_lib.scala 340:41]
  wire  _T_3366 = _T_3332[5:0] == 6'hc; // @[el2_lib.scala 340:41]
  wire  _T_3364 = _T_3332[5:0] == 6'hb; // @[el2_lib.scala 340:41]
  wire  _T_3362 = _T_3332[5:0] == 6'ha; // @[el2_lib.scala 340:41]
  wire [9:0] _T_3459 = {_T_3380,_T_3378,_T_3376,_T_3374,_T_3372,_T_3370,_T_3368,_T_3366,_T_3364,_T_3362}; // @[el2_lib.scala 343:69]
  wire  _T_3360 = _T_3332[5:0] == 6'h9; // @[el2_lib.scala 340:41]
  wire  _T_3358 = _T_3332[5:0] == 6'h8; // @[el2_lib.scala 340:41]
  wire  _T_3356 = _T_3332[5:0] == 6'h7; // @[el2_lib.scala 340:41]
  wire  _T_3354 = _T_3332[5:0] == 6'h6; // @[el2_lib.scala 340:41]
  wire  _T_3352 = _T_3332[5:0] == 6'h5; // @[el2_lib.scala 340:41]
  wire  _T_3350 = _T_3332[5:0] == 6'h4; // @[el2_lib.scala 340:41]
  wire  _T_3348 = _T_3332[5:0] == 6'h3; // @[el2_lib.scala 340:41]
  wire  _T_3346 = _T_3332[5:0] == 6'h2; // @[el2_lib.scala 340:41]
  wire  _T_3344 = _T_3332[5:0] == 6'h1; // @[el2_lib.scala 340:41]
  wire [18:0] _T_3460 = {_T_3459,_T_3360,_T_3358,_T_3356,_T_3354,_T_3352,_T_3350,_T_3348,_T_3346,_T_3344}; // @[el2_lib.scala 343:69]
  wire [38:0] _T_3480 = {_T_3478,_T_3469,_T_3460}; // @[el2_lib.scala 343:69]
  wire [7:0] _T_3435 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3441 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3435}; // @[Cat.scala 29:58]
  wire [38:0] _T_3481 = _T_3480 ^ _T_3441; // @[el2_lib.scala 343:76]
  wire [38:0] _T_3482 = _T_3336 ? _T_3481 : _T_3441; // @[el2_lib.scala 343:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3482[37:32],_T_3482[30:16],_T_3482[14:8],_T_3482[6:4],_T_3482[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 647:35]
  wire  _T_2955 = ~_T_2947[6]; // @[el2_lib.scala 336:55]
  wire  _T_2956 = _T_2949 & _T_2955; // @[el2_lib.scala 336:53]
  wire  _T_3340 = ~_T_3332[6]; // @[el2_lib.scala 336:55]
  wire  _T_3341 = _T_3334 & _T_3340; // @[el2_lib.scala 336:53]
  wire [1:0] iccm_double_ecc_error = {_T_2956,_T_3341}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 649:53]
  wire [63:0] _T_2707 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_2708 = {iccm_dma_rdata_1_muxed,_T_3097[37:32],_T_3097[30:16],_T_3097[14:8],_T_3097[6:4],_T_3097[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 651:54]
  reg [2:0] iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 652:74]
  reg  iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 657:76]
  reg [63:0] iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 661:75]
  wire  _T_2713 = _T_2678 & _T_2667; // @[el2_ifu_mem_ctl.scala 664:65]
  wire  _T_2716 = _T_2694 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 665:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_2717 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_2719 = _T_2716 ? {{1'd0}, _T_2717} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 665:8]
  wire [31:0] _T_2720 = _T_2713 ? io_dma_mem_addr : {{16'd0}, _T_2719}; // @[el2_ifu_mem_ctl.scala 664:25]
  wire  _T_3109 = _T_2947 == 7'h40; // @[el2_lib.scala 346:62]
  wire  _T_3110 = _T_3097[38] ^ _T_3109; // @[el2_lib.scala 346:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3110,_T_3097[31],_T_3097[15],_T_3097[7],_T_3097[3],_T_3097[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3494 = _T_3332 == 7'h40; // @[el2_lib.scala 346:62]
  wire  _T_3495 = _T_3482[38] ^ _T_3494; // @[el2_lib.scala 346:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3495,_T_3482[31],_T_3482[15],_T_3482[7],_T_3482[3],_T_3482[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3511 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 677:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 679:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 680:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 688:62]
  wire  _T_3519 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 682:76]
  wire  _T_3520 = io_iccm_rd_ecc_single_err & _T_3519; // @[el2_ifu_mem_ctl.scala 682:74]
  wire  _T_3522 = _T_3520 & _T_317; // @[el2_ifu_mem_ctl.scala 682:104]
  wire  iccm_ecc_write_status = _T_3522 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 682:127]
  wire  _T_3523 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 683:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3523 & _T_317; // @[el2_ifu_mem_ctl.scala 683:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 687:51]
  wire [13:0] _T_3528 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 686:102]
  wire [38:0] _T_3532 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3537 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 691:41]
  wire  _T_3538 = io_ifc_fetch_req_bf & _T_3537; // @[el2_ifu_mem_ctl.scala 691:39]
  wire  _T_3539 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 691:72]
  wire  _T_3540 = _T_3538 & _T_3539; // @[el2_ifu_mem_ctl.scala 691:70]
  wire  _T_3542 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 692:34]
  wire  _T_3543 = _T_2233 & _T_3542; // @[el2_ifu_mem_ctl.scala 692:32]
  wire  _T_3546 = _T_2249 & _T_3542; // @[el2_ifu_mem_ctl.scala 693:37]
  wire  _T_3547 = _T_3543 | _T_3546; // @[el2_ifu_mem_ctl.scala 692:88]
  wire  _T_3548 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 694:19]
  wire  _T_3550 = _T_3548 & _T_3542; // @[el2_ifu_mem_ctl.scala 694:41]
  wire  _T_3551 = _T_3547 | _T_3550; // @[el2_ifu_mem_ctl.scala 693:88]
  wire  _T_3552 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 695:19]
  wire  _T_3554 = _T_3552 & _T_3542; // @[el2_ifu_mem_ctl.scala 695:35]
  wire  _T_3555 = _T_3551 | _T_3554; // @[el2_ifu_mem_ctl.scala 694:88]
  wire  _T_3558 = _T_2248 & _T_3542; // @[el2_ifu_mem_ctl.scala 696:38]
  wire  _T_3559 = _T_3555 | _T_3558; // @[el2_ifu_mem_ctl.scala 695:88]
  wire  _T_3561 = _T_2249 & miss_state_en; // @[el2_ifu_mem_ctl.scala 697:37]
  wire  _T_3562 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 697:71]
  wire  _T_3563 = _T_3561 & _T_3562; // @[el2_ifu_mem_ctl.scala 697:54]
  wire  _T_3564 = _T_3559 | _T_3563; // @[el2_ifu_mem_ctl.scala 696:57]
  wire  _T_3565 = ~_T_3564; // @[el2_ifu_mem_ctl.scala 692:5]
  wire  _T_3566 = _T_3540 & _T_3565; // @[el2_ifu_mem_ctl.scala 691:96]
  wire  _T_3567 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 698:28]
  wire  _T_3569 = _T_3567 & _T_3537; // @[el2_ifu_mem_ctl.scala 698:50]
  wire  _T_3571 = _T_3569 & _T_3539; // @[el2_ifu_mem_ctl.scala 698:81]
  wire [1:0] _T_3574 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10012 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 795:74]
  wire  bus_wren_1 = _T_10012 & miss_pending; // @[el2_ifu_mem_ctl.scala 795:98]
  wire  _T_10011 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 795:74]
  wire  bus_wren_0 = _T_10011 & miss_pending; // @[el2_ifu_mem_ctl.scala 795:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3580 = ~_T_108; // @[el2_ifu_mem_ctl.scala 701:106]
  wire  _T_3581 = _T_2233 & _T_3580; // @[el2_ifu_mem_ctl.scala 701:104]
  wire  _T_3582 = _T_2249 | _T_3581; // @[el2_ifu_mem_ctl.scala 701:77]
  wire  _T_3586 = ~_T_51; // @[el2_ifu_mem_ctl.scala 701:172]
  wire  _T_3587 = _T_3582 & _T_3586; // @[el2_ifu_mem_ctl.scala 701:170]
  wire  _T_3588 = ~_T_3587; // @[el2_ifu_mem_ctl.scala 701:44]
  wire  _T_3592 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 704:64]
  wire  _T_3593 = ~_T_3592; // @[el2_ifu_mem_ctl.scala 704:50]
  wire  _T_3594 = _T_276 & _T_3593; // @[el2_ifu_mem_ctl.scala 704:48]
  wire  _T_3595 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 704:81]
  wire  ic_valid = _T_3594 & _T_3595; // @[el2_ifu_mem_ctl.scala 704:79]
  wire  _T_3597 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 705:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 708:14]
  wire  _T_3600 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 711:74]
  wire  _T_10009 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 794:45]
  wire  way_status_wr_en = _T_10009 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 794:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3600; // @[el2_ifu_mem_ctl.scala 711:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 713:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 790:41]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 721:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 723:132]
  wire  _T_3620 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3621 = _T_3620 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3622 = _T_3621 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3625 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3626 = _T_3625 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3627 = _T_3626 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3630 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3631 = _T_3630 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3632 = _T_3631 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3635 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3636 = _T_3635 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3637 = _T_3636 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3640 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3641 = _T_3640 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3642 = _T_3641 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3645 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3646 = _T_3645 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3647 = _T_3646 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3650 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3651 = _T_3650 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3652 = _T_3651 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3655 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 727:100]
  wire  _T_3656 = _T_3655 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 727:108]
  wire  _T_3657 = _T_3656 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3662 = _T_3621 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3667 = _T_3626 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3672 = _T_3631 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3677 = _T_3636 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3682 = _T_3641 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3687 = _T_3646 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3692 = _T_3651 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3697 = _T_3656 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3702 = _T_3621 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3707 = _T_3626 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3712 = _T_3631 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3717 = _T_3636 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3722 = _T_3641 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3727 = _T_3646 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3732 = _T_3651 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3737 = _T_3656 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3742 = _T_3621 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3747 = _T_3626 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3752 = _T_3631 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3757 = _T_3636 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3762 = _T_3641 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3767 = _T_3646 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3772 = _T_3651 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3777 = _T_3656 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3782 = _T_3621 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3787 = _T_3626 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3792 = _T_3631 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3797 = _T_3636 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3802 = _T_3641 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3807 = _T_3646 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3812 = _T_3651 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3817 = _T_3656 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3822 = _T_3621 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3827 = _T_3626 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3832 = _T_3631 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3837 = _T_3636 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3842 = _T_3641 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3847 = _T_3646 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3852 = _T_3651 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3857 = _T_3656 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3862 = _T_3621 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3867 = _T_3626 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3872 = _T_3631 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3877 = _T_3636 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3882 = _T_3641 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3887 = _T_3646 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3892 = _T_3651 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3897 = _T_3656 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3902 = _T_3621 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3907 = _T_3626 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3912 = _T_3631 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3917 = _T_3636 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3922 = _T_3641 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3927 = _T_3646 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3932 = _T_3651 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3937 = _T_3656 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3942 = _T_3621 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3947 = _T_3626 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3952 = _T_3631 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3957 = _T_3636 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3962 = _T_3641 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3967 = _T_3646 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3972 = _T_3651 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3977 = _T_3656 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3982 = _T_3621 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3987 = _T_3626 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3992 = _T_3631 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_3997 = _T_3636 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4002 = _T_3641 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4007 = _T_3646 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4012 = _T_3651 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4017 = _T_3656 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4022 = _T_3621 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4027 = _T_3626 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4032 = _T_3631 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4037 = _T_3636 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4042 = _T_3641 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4047 = _T_3646 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4052 = _T_3651 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4057 = _T_3656 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4062 = _T_3621 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4067 = _T_3626 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4072 = _T_3631 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4077 = _T_3636 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4082 = _T_3641 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4087 = _T_3646 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4092 = _T_3651 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4097 = _T_3656 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4102 = _T_3621 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4107 = _T_3626 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4112 = _T_3631 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4117 = _T_3636 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4122 = _T_3641 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4127 = _T_3646 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4132 = _T_3651 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4137 = _T_3656 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4142 = _T_3621 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4147 = _T_3626 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4152 = _T_3631 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4157 = _T_3636 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4162 = _T_3641 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4167 = _T_3646 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4172 = _T_3651 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4177 = _T_3656 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4182 = _T_3621 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4187 = _T_3626 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4192 = _T_3631 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4197 = _T_3636 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4202 = _T_3641 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4207 = _T_3646 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4212 = _T_3651 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4217 = _T_3656 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4222 = _T_3621 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4227 = _T_3626 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4232 = _T_3631 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4237 = _T_3636 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4242 = _T_3641 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4247 = _T_3646 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4252 = _T_3651 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_4257 = _T_3656 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 727:131]
  wire  _T_10015 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 797:84]
  wire  _T_10016 = _T_10015 & miss_pending; // @[el2_ifu_mem_ctl.scala 797:108]
  wire  bus_wren_last_1 = _T_10016 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 797:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 798:84]
  wire  _T_10018 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 799:73]
  wire  _T_10013 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 797:84]
  wire  _T_10014 = _T_10013 & miss_pending; // @[el2_ifu_mem_ctl.scala 797:108]
  wire  bus_wren_last_0 = _T_10014 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 797:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 798:84]
  wire  _T_10017 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 799:73]
  wire [1:0] ifu_tag_wren = {_T_10018,_T_10017}; // @[Cat.scala 29:58]
  wire [1:0] _T_10053 = _T_3600 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10053 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 833:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 740:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 742:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 746:14]
  wire  _T_4791 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 750:78]
  wire  _T_4793 = _T_4791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4795 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 751:70]
  wire  _T_4797 = _T_4795 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4798 = _T_4793 | _T_4797; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4799 = _T_4798 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire  _T_4803 = _T_4791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4807 = _T_4795 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4808 = _T_4803 | _T_4807; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4809 = _T_4808 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire [1:0] tag_valid_clken_0 = {_T_4809,_T_4799}; // @[Cat.scala 29:58]
  wire  _T_4811 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 750:78]
  wire  _T_4813 = _T_4811 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4815 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 751:70]
  wire  _T_4817 = _T_4815 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4818 = _T_4813 | _T_4817; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4819 = _T_4818 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire  _T_4823 = _T_4811 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4827 = _T_4815 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4828 = _T_4823 | _T_4827; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4829 = _T_4828 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire [1:0] tag_valid_clken_1 = {_T_4829,_T_4819}; // @[Cat.scala 29:58]
  wire  _T_4831 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 750:78]
  wire  _T_4833 = _T_4831 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4835 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 751:70]
  wire  _T_4837 = _T_4835 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4838 = _T_4833 | _T_4837; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4839 = _T_4838 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire  _T_4843 = _T_4831 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4847 = _T_4835 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4848 = _T_4843 | _T_4847; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4849 = _T_4848 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire [1:0] tag_valid_clken_2 = {_T_4849,_T_4839}; // @[Cat.scala 29:58]
  wire  _T_4851 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 750:78]
  wire  _T_4853 = _T_4851 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4855 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 751:70]
  wire  _T_4857 = _T_4855 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4858 = _T_4853 | _T_4857; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4859 = _T_4858 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire  _T_4863 = _T_4851 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:87]
  wire  _T_4867 = _T_4855 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:79]
  wire  _T_4868 = _T_4863 | _T_4867; // @[el2_ifu_mem_ctl.scala 750:109]
  wire  _T_4869 = _T_4868 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:102]
  wire [1:0] tag_valid_clken_3 = {_T_4869,_T_4859}; // @[Cat.scala 29:58]
  wire  _T_4872 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 759:66]
  wire  _T_4873 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 759:93]
  wire  _T_4874 = _T_4872 & _T_4873; // @[el2_ifu_mem_ctl.scala 759:91]
  wire  _T_4877 = _T_4399 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4878 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4880 = _T_4878 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_4881 = _T_4877 | _T_4880; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_4882 = _T_4881 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_4884 = _T_4882 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_4894 = _T_4400 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4895 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4897 = _T_4895 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_4898 = _T_4894 | _T_4897; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_4899 = _T_4898 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_4901 = _T_4899 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_4911 = _T_4401 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4912 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4914 = _T_4912 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_4915 = _T_4911 | _T_4914; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_4916 = _T_4915 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_4918 = _T_4916 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_4928 = _T_4402 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4929 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4931 = _T_4929 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_4932 = _T_4928 | _T_4931; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_4933 = _T_4932 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_4935 = _T_4933 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_4945 = _T_4403 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4946 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4948 = _T_4946 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_4949 = _T_4945 | _T_4948; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_4950 = _T_4949 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_4952 = _T_4950 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_4962 = _T_4404 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4963 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4965 = _T_4963 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_4966 = _T_4962 | _T_4965; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_4967 = _T_4966 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_4969 = _T_4967 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_4979 = _T_4405 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4980 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4982 = _T_4980 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_4983 = _T_4979 | _T_4982; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_4984 = _T_4983 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_4986 = _T_4984 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_4996 = _T_4406 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_4997 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_4999 = _T_4997 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5000 = _T_4996 | _T_4999; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5001 = _T_5000 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5003 = _T_5001 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5013 = _T_4407 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5014 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5016 = _T_5014 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5017 = _T_5013 | _T_5016; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5018 = _T_5017 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5020 = _T_5018 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5030 = _T_4408 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5031 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5033 = _T_5031 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5034 = _T_5030 | _T_5033; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5035 = _T_5034 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5037 = _T_5035 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5047 = _T_4409 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5048 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5050 = _T_5048 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5051 = _T_5047 | _T_5050; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5052 = _T_5051 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5054 = _T_5052 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5064 = _T_4410 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5065 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5067 = _T_5065 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5068 = _T_5064 | _T_5067; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5069 = _T_5068 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5071 = _T_5069 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5081 = _T_4411 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5082 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5084 = _T_5082 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5085 = _T_5081 | _T_5084; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5086 = _T_5085 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5088 = _T_5086 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5098 = _T_4412 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5099 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5101 = _T_5099 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5102 = _T_5098 | _T_5101; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5103 = _T_5102 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5105 = _T_5103 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5115 = _T_4413 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5116 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5118 = _T_5116 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5119 = _T_5115 | _T_5118; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5120 = _T_5119 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5122 = _T_5120 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5132 = _T_4414 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5133 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5135 = _T_5133 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5136 = _T_5132 | _T_5135; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5137 = _T_5136 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5139 = _T_5137 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5149 = _T_4415 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5150 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5152 = _T_5150 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5153 = _T_5149 | _T_5152; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5154 = _T_5153 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5156 = _T_5154 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5166 = _T_4416 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5167 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5169 = _T_5167 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5170 = _T_5166 | _T_5169; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5171 = _T_5170 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5173 = _T_5171 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5183 = _T_4417 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5184 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5186 = _T_5184 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5187 = _T_5183 | _T_5186; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5188 = _T_5187 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5190 = _T_5188 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5200 = _T_4418 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5201 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5203 = _T_5201 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5204 = _T_5200 | _T_5203; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5205 = _T_5204 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5207 = _T_5205 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5217 = _T_4419 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5218 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5220 = _T_5218 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5221 = _T_5217 | _T_5220; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5222 = _T_5221 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5224 = _T_5222 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5234 = _T_4420 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5235 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5237 = _T_5235 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5238 = _T_5234 | _T_5237; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5239 = _T_5238 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5241 = _T_5239 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5251 = _T_4421 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5252 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5254 = _T_5252 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5255 = _T_5251 | _T_5254; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5256 = _T_5255 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5258 = _T_5256 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5268 = _T_4422 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5269 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5271 = _T_5269 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5272 = _T_5268 | _T_5271; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5273 = _T_5272 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5275 = _T_5273 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5285 = _T_4423 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5286 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5288 = _T_5286 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5289 = _T_5285 | _T_5288; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5290 = _T_5289 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5292 = _T_5290 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5302 = _T_4424 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5303 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5305 = _T_5303 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5306 = _T_5302 | _T_5305; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5307 = _T_5306 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5309 = _T_5307 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5319 = _T_4425 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5320 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5322 = _T_5320 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5323 = _T_5319 | _T_5322; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5324 = _T_5323 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5326 = _T_5324 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5336 = _T_4426 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5337 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5339 = _T_5337 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5340 = _T_5336 | _T_5339; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5341 = _T_5340 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5343 = _T_5341 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5353 = _T_4427 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5354 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5356 = _T_5354 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5357 = _T_5353 | _T_5356; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5358 = _T_5357 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5360 = _T_5358 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5370 = _T_4428 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5371 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5373 = _T_5371 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5374 = _T_5370 | _T_5373; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5375 = _T_5374 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5377 = _T_5375 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5387 = _T_4429 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5388 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5390 = _T_5388 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5391 = _T_5387 | _T_5390; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5392 = _T_5391 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5394 = _T_5392 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5404 = _T_4430 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5405 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5407 = _T_5405 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5408 = _T_5404 | _T_5407; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5409 = _T_5408 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5411 = _T_5409 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5421 = _T_4399 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5424 = _T_4878 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5425 = _T_5421 | _T_5424; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5426 = _T_5425 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5428 = _T_5426 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5438 = _T_4400 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5441 = _T_4895 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5442 = _T_5438 | _T_5441; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5443 = _T_5442 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5445 = _T_5443 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5455 = _T_4401 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5458 = _T_4912 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5459 = _T_5455 | _T_5458; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5460 = _T_5459 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5462 = _T_5460 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5472 = _T_4402 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5475 = _T_4929 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5476 = _T_5472 | _T_5475; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5477 = _T_5476 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5479 = _T_5477 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5489 = _T_4403 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5492 = _T_4946 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5493 = _T_5489 | _T_5492; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5494 = _T_5493 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5496 = _T_5494 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5506 = _T_4404 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5509 = _T_4963 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5510 = _T_5506 | _T_5509; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5511 = _T_5510 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5513 = _T_5511 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5523 = _T_4405 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5526 = _T_4980 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5527 = _T_5523 | _T_5526; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5528 = _T_5527 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5530 = _T_5528 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5540 = _T_4406 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5543 = _T_4997 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5544 = _T_5540 | _T_5543; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5545 = _T_5544 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5547 = _T_5545 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5557 = _T_4407 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5560 = _T_5014 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5561 = _T_5557 | _T_5560; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5562 = _T_5561 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5564 = _T_5562 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5574 = _T_4408 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5577 = _T_5031 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5578 = _T_5574 | _T_5577; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5579 = _T_5578 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5581 = _T_5579 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5591 = _T_4409 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5594 = _T_5048 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5595 = _T_5591 | _T_5594; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5596 = _T_5595 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5598 = _T_5596 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5608 = _T_4410 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5611 = _T_5065 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5612 = _T_5608 | _T_5611; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5613 = _T_5612 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5615 = _T_5613 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5625 = _T_4411 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5628 = _T_5082 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5629 = _T_5625 | _T_5628; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5630 = _T_5629 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5632 = _T_5630 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5642 = _T_4412 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5645 = _T_5099 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5646 = _T_5642 | _T_5645; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5647 = _T_5646 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5649 = _T_5647 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5659 = _T_4413 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5662 = _T_5116 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5663 = _T_5659 | _T_5662; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5664 = _T_5663 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5666 = _T_5664 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5676 = _T_4414 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5679 = _T_5133 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5680 = _T_5676 | _T_5679; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5681 = _T_5680 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5683 = _T_5681 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5693 = _T_4415 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5696 = _T_5150 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5697 = _T_5693 | _T_5696; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5698 = _T_5697 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5700 = _T_5698 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5710 = _T_4416 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5713 = _T_5167 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5714 = _T_5710 | _T_5713; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5715 = _T_5714 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5717 = _T_5715 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5727 = _T_4417 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5730 = _T_5184 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5731 = _T_5727 | _T_5730; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5732 = _T_5731 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5734 = _T_5732 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5744 = _T_4418 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5747 = _T_5201 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5748 = _T_5744 | _T_5747; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5749 = _T_5748 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5751 = _T_5749 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5761 = _T_4419 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5764 = _T_5218 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5765 = _T_5761 | _T_5764; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5766 = _T_5765 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5768 = _T_5766 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5778 = _T_4420 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5781 = _T_5235 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5782 = _T_5778 | _T_5781; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5783 = _T_5782 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5785 = _T_5783 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5795 = _T_4421 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5798 = _T_5252 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5799 = _T_5795 | _T_5798; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5800 = _T_5799 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5802 = _T_5800 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5812 = _T_4422 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5815 = _T_5269 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5816 = _T_5812 | _T_5815; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5817 = _T_5816 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5819 = _T_5817 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5829 = _T_4423 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5832 = _T_5286 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5833 = _T_5829 | _T_5832; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5834 = _T_5833 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5836 = _T_5834 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5846 = _T_4424 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5849 = _T_5303 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5850 = _T_5846 | _T_5849; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5851 = _T_5850 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5853 = _T_5851 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5863 = _T_4425 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5866 = _T_5320 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5867 = _T_5863 | _T_5866; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5868 = _T_5867 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5870 = _T_5868 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5880 = _T_4426 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5883 = _T_5337 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5884 = _T_5880 | _T_5883; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5885 = _T_5884 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5887 = _T_5885 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5897 = _T_4427 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5900 = _T_5354 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5901 = _T_5897 | _T_5900; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5902 = _T_5901 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5904 = _T_5902 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5914 = _T_4428 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5917 = _T_5371 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5918 = _T_5914 | _T_5917; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5919 = _T_5918 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5921 = _T_5919 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5931 = _T_4429 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5934 = _T_5388 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5935 = _T_5931 | _T_5934; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5936 = _T_5935 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5938 = _T_5936 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5948 = _T_4430 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5951 = _T_5405 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5952 = _T_5948 | _T_5951; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5953 = _T_5952 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5955 = _T_5953 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5965 = _T_4431 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5966 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5968 = _T_5966 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5969 = _T_5965 | _T_5968; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5970 = _T_5969 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5972 = _T_5970 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5982 = _T_4432 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_5983 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_5985 = _T_5983 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_5986 = _T_5982 | _T_5985; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_5987 = _T_5986 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_5989 = _T_5987 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_5999 = _T_4433 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6000 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6002 = _T_6000 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6003 = _T_5999 | _T_6002; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6004 = _T_6003 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6006 = _T_6004 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6016 = _T_4434 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6017 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6019 = _T_6017 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6020 = _T_6016 | _T_6019; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6021 = _T_6020 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6023 = _T_6021 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6033 = _T_4435 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6034 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6036 = _T_6034 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6037 = _T_6033 | _T_6036; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6038 = _T_6037 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6040 = _T_6038 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6050 = _T_4436 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6051 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6053 = _T_6051 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6054 = _T_6050 | _T_6053; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6055 = _T_6054 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6057 = _T_6055 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6067 = _T_4437 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6068 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6070 = _T_6068 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6071 = _T_6067 | _T_6070; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6072 = _T_6071 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6074 = _T_6072 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6084 = _T_4438 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6085 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6087 = _T_6085 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6088 = _T_6084 | _T_6087; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6089 = _T_6088 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6091 = _T_6089 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6101 = _T_4439 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6102 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6104 = _T_6102 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6105 = _T_6101 | _T_6104; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6106 = _T_6105 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6108 = _T_6106 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6118 = _T_4440 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6119 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6121 = _T_6119 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6122 = _T_6118 | _T_6121; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6123 = _T_6122 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6125 = _T_6123 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6135 = _T_4441 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6136 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6138 = _T_6136 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6139 = _T_6135 | _T_6138; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6140 = _T_6139 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6142 = _T_6140 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6152 = _T_4442 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6153 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6155 = _T_6153 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6156 = _T_6152 | _T_6155; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6157 = _T_6156 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6159 = _T_6157 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6169 = _T_4443 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6170 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6172 = _T_6170 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6173 = _T_6169 | _T_6172; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6174 = _T_6173 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6176 = _T_6174 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6186 = _T_4444 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6187 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6189 = _T_6187 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6190 = _T_6186 | _T_6189; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6191 = _T_6190 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6193 = _T_6191 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6203 = _T_4445 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6204 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6206 = _T_6204 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6207 = _T_6203 | _T_6206; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6208 = _T_6207 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6210 = _T_6208 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6220 = _T_4446 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6221 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6223 = _T_6221 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6224 = _T_6220 | _T_6223; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6225 = _T_6224 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6227 = _T_6225 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6237 = _T_4447 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6238 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6240 = _T_6238 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6241 = _T_6237 | _T_6240; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6242 = _T_6241 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6244 = _T_6242 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6254 = _T_4448 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6255 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6257 = _T_6255 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6258 = _T_6254 | _T_6257; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6259 = _T_6258 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6261 = _T_6259 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6271 = _T_4449 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6272 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6274 = _T_6272 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6275 = _T_6271 | _T_6274; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6276 = _T_6275 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6278 = _T_6276 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6288 = _T_4450 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6289 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6291 = _T_6289 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6292 = _T_6288 | _T_6291; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6293 = _T_6292 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6295 = _T_6293 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6305 = _T_4451 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6306 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6308 = _T_6306 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6309 = _T_6305 | _T_6308; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6310 = _T_6309 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6312 = _T_6310 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6322 = _T_4452 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6323 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6325 = _T_6323 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6326 = _T_6322 | _T_6325; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6327 = _T_6326 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6329 = _T_6327 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6339 = _T_4453 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6340 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6342 = _T_6340 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6343 = _T_6339 | _T_6342; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6344 = _T_6343 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6346 = _T_6344 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6356 = _T_4454 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6357 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6359 = _T_6357 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6360 = _T_6356 | _T_6359; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6361 = _T_6360 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6363 = _T_6361 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6373 = _T_4455 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6374 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6376 = _T_6374 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6377 = _T_6373 | _T_6376; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6378 = _T_6377 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6380 = _T_6378 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6390 = _T_4456 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6391 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6393 = _T_6391 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6394 = _T_6390 | _T_6393; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6395 = _T_6394 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6397 = _T_6395 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6407 = _T_4457 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6408 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6410 = _T_6408 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6411 = _T_6407 | _T_6410; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6412 = _T_6411 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6414 = _T_6412 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6424 = _T_4458 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6425 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6427 = _T_6425 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6428 = _T_6424 | _T_6427; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6429 = _T_6428 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6431 = _T_6429 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6441 = _T_4459 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6442 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6444 = _T_6442 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6445 = _T_6441 | _T_6444; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6446 = _T_6445 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6448 = _T_6446 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6458 = _T_4460 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6459 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6461 = _T_6459 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6462 = _T_6458 | _T_6461; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6463 = _T_6462 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6465 = _T_6463 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6475 = _T_4461 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6476 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6478 = _T_6476 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6479 = _T_6475 | _T_6478; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6480 = _T_6479 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6482 = _T_6480 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6492 = _T_4462 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6493 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_6495 = _T_6493 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6496 = _T_6492 | _T_6495; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6497 = _T_6496 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6499 = _T_6497 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6509 = _T_4431 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6512 = _T_5966 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6513 = _T_6509 | _T_6512; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6514 = _T_6513 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6516 = _T_6514 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6526 = _T_4432 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6529 = _T_5983 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6530 = _T_6526 | _T_6529; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6531 = _T_6530 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6533 = _T_6531 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6543 = _T_4433 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6546 = _T_6000 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6547 = _T_6543 | _T_6546; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6548 = _T_6547 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6550 = _T_6548 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6560 = _T_4434 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6563 = _T_6017 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6564 = _T_6560 | _T_6563; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6565 = _T_6564 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6567 = _T_6565 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6577 = _T_4435 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6580 = _T_6034 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6581 = _T_6577 | _T_6580; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6582 = _T_6581 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6584 = _T_6582 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6594 = _T_4436 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6597 = _T_6051 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6598 = _T_6594 | _T_6597; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6599 = _T_6598 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6601 = _T_6599 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6611 = _T_4437 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6614 = _T_6068 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6615 = _T_6611 | _T_6614; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6616 = _T_6615 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6618 = _T_6616 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6628 = _T_4438 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6631 = _T_6085 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6632 = _T_6628 | _T_6631; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6633 = _T_6632 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6635 = _T_6633 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6645 = _T_4439 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6648 = _T_6102 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6649 = _T_6645 | _T_6648; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6650 = _T_6649 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6652 = _T_6650 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6662 = _T_4440 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6665 = _T_6119 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6666 = _T_6662 | _T_6665; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6667 = _T_6666 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6669 = _T_6667 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6679 = _T_4441 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6682 = _T_6136 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6683 = _T_6679 | _T_6682; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6684 = _T_6683 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6686 = _T_6684 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6696 = _T_4442 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6699 = _T_6153 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6700 = _T_6696 | _T_6699; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6701 = _T_6700 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6703 = _T_6701 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6713 = _T_4443 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6716 = _T_6170 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6717 = _T_6713 | _T_6716; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6718 = _T_6717 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6720 = _T_6718 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6730 = _T_4444 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6733 = _T_6187 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6734 = _T_6730 | _T_6733; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6735 = _T_6734 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6737 = _T_6735 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6747 = _T_4445 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6750 = _T_6204 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6751 = _T_6747 | _T_6750; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6752 = _T_6751 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6754 = _T_6752 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6764 = _T_4446 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6767 = _T_6221 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6768 = _T_6764 | _T_6767; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6769 = _T_6768 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6771 = _T_6769 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6781 = _T_4447 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6784 = _T_6238 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6785 = _T_6781 | _T_6784; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6786 = _T_6785 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6788 = _T_6786 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6798 = _T_4448 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6801 = _T_6255 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6802 = _T_6798 | _T_6801; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6803 = _T_6802 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6805 = _T_6803 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6815 = _T_4449 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6818 = _T_6272 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6819 = _T_6815 | _T_6818; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6820 = _T_6819 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6822 = _T_6820 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6832 = _T_4450 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6835 = _T_6289 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6836 = _T_6832 | _T_6835; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6837 = _T_6836 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6839 = _T_6837 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6849 = _T_4451 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6852 = _T_6306 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6853 = _T_6849 | _T_6852; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6854 = _T_6853 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6856 = _T_6854 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6866 = _T_4452 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6869 = _T_6323 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6870 = _T_6866 | _T_6869; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6871 = _T_6870 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6873 = _T_6871 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6883 = _T_4453 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6886 = _T_6340 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6887 = _T_6883 | _T_6886; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6888 = _T_6887 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6890 = _T_6888 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6900 = _T_4454 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6903 = _T_6357 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6904 = _T_6900 | _T_6903; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6905 = _T_6904 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6907 = _T_6905 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6917 = _T_4455 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6920 = _T_6374 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6921 = _T_6917 | _T_6920; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6922 = _T_6921 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6924 = _T_6922 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6934 = _T_4456 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6937 = _T_6391 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6938 = _T_6934 | _T_6937; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6939 = _T_6938 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6941 = _T_6939 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6951 = _T_4457 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6954 = _T_6408 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6955 = _T_6951 | _T_6954; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6956 = _T_6955 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6958 = _T_6956 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6968 = _T_4458 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6971 = _T_6425 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6972 = _T_6968 | _T_6971; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6973 = _T_6972 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6975 = _T_6973 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_6985 = _T_4459 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_6988 = _T_6442 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_6989 = _T_6985 | _T_6988; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_6990 = _T_6989 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_6992 = _T_6990 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7002 = _T_4460 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7005 = _T_6459 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7006 = _T_7002 | _T_7005; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7007 = _T_7006 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7009 = _T_7007 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7019 = _T_4461 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7022 = _T_6476 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7023 = _T_7019 | _T_7022; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7024 = _T_7023 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7026 = _T_7024 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7036 = _T_4462 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7039 = _T_6493 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7040 = _T_7036 | _T_7039; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7041 = _T_7040 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7043 = _T_7041 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7053 = _T_4463 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7054 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7056 = _T_7054 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7057 = _T_7053 | _T_7056; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7058 = _T_7057 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7060 = _T_7058 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7070 = _T_4464 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7071 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7073 = _T_7071 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7074 = _T_7070 | _T_7073; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7075 = _T_7074 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7077 = _T_7075 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7087 = _T_4465 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7088 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7090 = _T_7088 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7091 = _T_7087 | _T_7090; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7092 = _T_7091 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7094 = _T_7092 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7104 = _T_4466 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7105 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7107 = _T_7105 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7108 = _T_7104 | _T_7107; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7109 = _T_7108 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7111 = _T_7109 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7121 = _T_4467 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7122 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7124 = _T_7122 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7125 = _T_7121 | _T_7124; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7126 = _T_7125 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7128 = _T_7126 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7138 = _T_4468 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7139 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7141 = _T_7139 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7142 = _T_7138 | _T_7141; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7143 = _T_7142 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7145 = _T_7143 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7155 = _T_4469 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7156 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7158 = _T_7156 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7159 = _T_7155 | _T_7158; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7160 = _T_7159 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7162 = _T_7160 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7172 = _T_4470 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7173 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7175 = _T_7173 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7176 = _T_7172 | _T_7175; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7177 = _T_7176 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7179 = _T_7177 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7189 = _T_4471 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7190 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7192 = _T_7190 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7193 = _T_7189 | _T_7192; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7194 = _T_7193 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7196 = _T_7194 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7206 = _T_4472 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7207 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7209 = _T_7207 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7210 = _T_7206 | _T_7209; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7211 = _T_7210 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7213 = _T_7211 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7223 = _T_4473 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7224 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7226 = _T_7224 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7227 = _T_7223 | _T_7226; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7228 = _T_7227 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7230 = _T_7228 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7240 = _T_4474 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7241 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7243 = _T_7241 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7244 = _T_7240 | _T_7243; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7245 = _T_7244 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7247 = _T_7245 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7257 = _T_4475 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7258 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7260 = _T_7258 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7261 = _T_7257 | _T_7260; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7262 = _T_7261 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7264 = _T_7262 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7274 = _T_4476 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7275 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7277 = _T_7275 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7278 = _T_7274 | _T_7277; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7279 = _T_7278 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7281 = _T_7279 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7291 = _T_4477 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7292 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7294 = _T_7292 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7295 = _T_7291 | _T_7294; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7296 = _T_7295 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7298 = _T_7296 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7308 = _T_4478 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7309 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7311 = _T_7309 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7312 = _T_7308 | _T_7311; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7313 = _T_7312 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7315 = _T_7313 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7325 = _T_4479 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7326 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7328 = _T_7326 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7329 = _T_7325 | _T_7328; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7330 = _T_7329 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7332 = _T_7330 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7342 = _T_4480 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7343 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7345 = _T_7343 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7346 = _T_7342 | _T_7345; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7347 = _T_7346 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7349 = _T_7347 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7359 = _T_4481 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7360 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7362 = _T_7360 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7363 = _T_7359 | _T_7362; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7364 = _T_7363 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7366 = _T_7364 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7376 = _T_4482 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7377 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7379 = _T_7377 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7380 = _T_7376 | _T_7379; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7381 = _T_7380 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7383 = _T_7381 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7393 = _T_4483 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7394 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7396 = _T_7394 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7397 = _T_7393 | _T_7396; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7398 = _T_7397 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7400 = _T_7398 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7410 = _T_4484 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7411 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7413 = _T_7411 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7414 = _T_7410 | _T_7413; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7415 = _T_7414 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7417 = _T_7415 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7427 = _T_4485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7428 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7430 = _T_7428 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7431 = _T_7427 | _T_7430; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7432 = _T_7431 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7434 = _T_7432 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7444 = _T_4486 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7445 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7447 = _T_7445 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7448 = _T_7444 | _T_7447; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7449 = _T_7448 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7451 = _T_7449 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7461 = _T_4487 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7462 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7464 = _T_7462 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7465 = _T_7461 | _T_7464; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7466 = _T_7465 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7468 = _T_7466 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7478 = _T_4488 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7479 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7481 = _T_7479 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7482 = _T_7478 | _T_7481; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7483 = _T_7482 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7485 = _T_7483 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7495 = _T_4489 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7496 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7498 = _T_7496 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7499 = _T_7495 | _T_7498; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7500 = _T_7499 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7502 = _T_7500 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7512 = _T_4490 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7513 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7515 = _T_7513 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7516 = _T_7512 | _T_7515; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7517 = _T_7516 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7519 = _T_7517 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7529 = _T_4491 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7530 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7532 = _T_7530 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7533 = _T_7529 | _T_7532; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7534 = _T_7533 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7536 = _T_7534 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7546 = _T_4492 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7547 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7549 = _T_7547 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7550 = _T_7546 | _T_7549; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7551 = _T_7550 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7553 = _T_7551 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7563 = _T_4493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7564 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7566 = _T_7564 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7567 = _T_7563 | _T_7566; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7568 = _T_7567 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7570 = _T_7568 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7580 = _T_4494 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7581 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_7583 = _T_7581 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7584 = _T_7580 | _T_7583; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7585 = _T_7584 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7587 = _T_7585 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7597 = _T_4463 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7600 = _T_7054 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7601 = _T_7597 | _T_7600; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7602 = _T_7601 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7604 = _T_7602 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7614 = _T_4464 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7617 = _T_7071 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7618 = _T_7614 | _T_7617; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7619 = _T_7618 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7621 = _T_7619 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7631 = _T_4465 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7634 = _T_7088 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7635 = _T_7631 | _T_7634; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7636 = _T_7635 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7638 = _T_7636 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7648 = _T_4466 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7651 = _T_7105 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7652 = _T_7648 | _T_7651; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7653 = _T_7652 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7655 = _T_7653 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7665 = _T_4467 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7668 = _T_7122 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7669 = _T_7665 | _T_7668; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7670 = _T_7669 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7672 = _T_7670 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7682 = _T_4468 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7685 = _T_7139 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7686 = _T_7682 | _T_7685; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7687 = _T_7686 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7689 = _T_7687 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7699 = _T_4469 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7702 = _T_7156 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7703 = _T_7699 | _T_7702; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7704 = _T_7703 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7706 = _T_7704 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7716 = _T_4470 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7719 = _T_7173 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7720 = _T_7716 | _T_7719; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7721 = _T_7720 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7723 = _T_7721 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7733 = _T_4471 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7736 = _T_7190 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7737 = _T_7733 | _T_7736; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7738 = _T_7737 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7740 = _T_7738 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7750 = _T_4472 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7753 = _T_7207 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7754 = _T_7750 | _T_7753; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7755 = _T_7754 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7757 = _T_7755 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7767 = _T_4473 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7770 = _T_7224 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7771 = _T_7767 | _T_7770; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7772 = _T_7771 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7774 = _T_7772 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7784 = _T_4474 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7787 = _T_7241 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7788 = _T_7784 | _T_7787; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7789 = _T_7788 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7791 = _T_7789 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7801 = _T_4475 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7804 = _T_7258 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7805 = _T_7801 | _T_7804; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7806 = _T_7805 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7808 = _T_7806 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7818 = _T_4476 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7821 = _T_7275 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7822 = _T_7818 | _T_7821; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7823 = _T_7822 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7825 = _T_7823 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7835 = _T_4477 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7838 = _T_7292 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7839 = _T_7835 | _T_7838; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7840 = _T_7839 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7842 = _T_7840 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7852 = _T_4478 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7855 = _T_7309 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7856 = _T_7852 | _T_7855; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7857 = _T_7856 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7859 = _T_7857 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7869 = _T_4479 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7872 = _T_7326 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7873 = _T_7869 | _T_7872; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7874 = _T_7873 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7876 = _T_7874 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7886 = _T_4480 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7889 = _T_7343 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7890 = _T_7886 | _T_7889; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7891 = _T_7890 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7893 = _T_7891 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7903 = _T_4481 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7906 = _T_7360 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7907 = _T_7903 | _T_7906; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7908 = _T_7907 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7910 = _T_7908 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7920 = _T_4482 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7923 = _T_7377 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7924 = _T_7920 | _T_7923; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7925 = _T_7924 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7927 = _T_7925 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7937 = _T_4483 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7940 = _T_7394 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7941 = _T_7937 | _T_7940; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7942 = _T_7941 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7944 = _T_7942 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7954 = _T_4484 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7957 = _T_7411 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7958 = _T_7954 | _T_7957; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7959 = _T_7958 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7961 = _T_7959 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7971 = _T_4485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7974 = _T_7428 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7975 = _T_7971 | _T_7974; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7976 = _T_7975 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7978 = _T_7976 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_7988 = _T_4486 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_7991 = _T_7445 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_7992 = _T_7988 | _T_7991; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_7993 = _T_7992 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_7995 = _T_7993 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8005 = _T_4487 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8008 = _T_7462 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8009 = _T_8005 | _T_8008; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8010 = _T_8009 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8012 = _T_8010 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8022 = _T_4488 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8025 = _T_7479 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8026 = _T_8022 | _T_8025; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8027 = _T_8026 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8029 = _T_8027 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8039 = _T_4489 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8042 = _T_7496 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8043 = _T_8039 | _T_8042; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8044 = _T_8043 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8046 = _T_8044 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8056 = _T_4490 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8059 = _T_7513 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8060 = _T_8056 | _T_8059; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8061 = _T_8060 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8063 = _T_8061 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8073 = _T_4491 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8076 = _T_7530 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8077 = _T_8073 | _T_8076; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8078 = _T_8077 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8080 = _T_8078 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8090 = _T_4492 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8093 = _T_7547 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8094 = _T_8090 | _T_8093; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8095 = _T_8094 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8097 = _T_8095 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8107 = _T_4493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8110 = _T_7564 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8111 = _T_8107 | _T_8110; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8112 = _T_8111 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8114 = _T_8112 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8124 = _T_4494 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8127 = _T_7581 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8128 = _T_8124 | _T_8127; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8129 = _T_8128 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8131 = _T_8129 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8141 = _T_4495 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8142 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8144 = _T_8142 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8145 = _T_8141 | _T_8144; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8146 = _T_8145 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8148 = _T_8146 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8158 = _T_4496 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8159 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8161 = _T_8159 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8162 = _T_8158 | _T_8161; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8163 = _T_8162 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8165 = _T_8163 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8175 = _T_4497 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8176 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8178 = _T_8176 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8179 = _T_8175 | _T_8178; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8180 = _T_8179 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8182 = _T_8180 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8192 = _T_4498 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8193 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8195 = _T_8193 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8196 = _T_8192 | _T_8195; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8197 = _T_8196 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8199 = _T_8197 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8209 = _T_4499 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8210 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8212 = _T_8210 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8213 = _T_8209 | _T_8212; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8214 = _T_8213 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8216 = _T_8214 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8226 = _T_4500 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8227 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8229 = _T_8227 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8230 = _T_8226 | _T_8229; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8231 = _T_8230 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8233 = _T_8231 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8243 = _T_4501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8244 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8246 = _T_8244 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8247 = _T_8243 | _T_8246; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8248 = _T_8247 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8250 = _T_8248 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8260 = _T_4502 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8261 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8263 = _T_8261 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8264 = _T_8260 | _T_8263; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8265 = _T_8264 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8267 = _T_8265 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8277 = _T_4503 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8278 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8280 = _T_8278 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8281 = _T_8277 | _T_8280; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8282 = _T_8281 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8284 = _T_8282 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8294 = _T_4504 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8295 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8297 = _T_8295 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8298 = _T_8294 | _T_8297; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8299 = _T_8298 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8301 = _T_8299 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8311 = _T_4505 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8312 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8314 = _T_8312 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8315 = _T_8311 | _T_8314; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8316 = _T_8315 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8318 = _T_8316 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8328 = _T_4506 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8329 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8331 = _T_8329 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8332 = _T_8328 | _T_8331; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8333 = _T_8332 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8335 = _T_8333 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8345 = _T_4507 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8346 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8348 = _T_8346 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8349 = _T_8345 | _T_8348; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8350 = _T_8349 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8352 = _T_8350 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8362 = _T_4508 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8363 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8365 = _T_8363 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8366 = _T_8362 | _T_8365; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8367 = _T_8366 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8369 = _T_8367 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8379 = _T_4509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8380 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8382 = _T_8380 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8383 = _T_8379 | _T_8382; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8384 = _T_8383 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8386 = _T_8384 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8396 = _T_4510 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8397 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8399 = _T_8397 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8400 = _T_8396 | _T_8399; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8401 = _T_8400 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8403 = _T_8401 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8413 = _T_4511 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8414 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8416 = _T_8414 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8417 = _T_8413 | _T_8416; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8418 = _T_8417 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8420 = _T_8418 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8430 = _T_4512 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8431 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8433 = _T_8431 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8434 = _T_8430 | _T_8433; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8435 = _T_8434 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8437 = _T_8435 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8447 = _T_4513 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8448 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8450 = _T_8448 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8451 = _T_8447 | _T_8450; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8452 = _T_8451 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8454 = _T_8452 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8464 = _T_4514 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8465 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8467 = _T_8465 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8468 = _T_8464 | _T_8467; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8469 = _T_8468 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8471 = _T_8469 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8481 = _T_4515 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8482 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8484 = _T_8482 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8485 = _T_8481 | _T_8484; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8486 = _T_8485 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8488 = _T_8486 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8498 = _T_4516 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8499 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8501 = _T_8499 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8502 = _T_8498 | _T_8501; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8503 = _T_8502 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8505 = _T_8503 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8515 = _T_4517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8516 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8518 = _T_8516 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8519 = _T_8515 | _T_8518; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8520 = _T_8519 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8522 = _T_8520 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8532 = _T_4518 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8533 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8535 = _T_8533 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8536 = _T_8532 | _T_8535; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8537 = _T_8536 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8539 = _T_8537 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8549 = _T_4519 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8550 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8552 = _T_8550 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8553 = _T_8549 | _T_8552; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8554 = _T_8553 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8556 = _T_8554 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8566 = _T_4520 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8567 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8569 = _T_8567 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8570 = _T_8566 | _T_8569; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8571 = _T_8570 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8573 = _T_8571 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8583 = _T_4521 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8584 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8586 = _T_8584 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8587 = _T_8583 | _T_8586; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8588 = _T_8587 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8590 = _T_8588 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8600 = _T_4522 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8601 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8603 = _T_8601 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8604 = _T_8600 | _T_8603; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8605 = _T_8604 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8607 = _T_8605 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8617 = _T_4523 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8618 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8620 = _T_8618 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8621 = _T_8617 | _T_8620; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8622 = _T_8621 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8624 = _T_8622 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8634 = _T_4524 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8635 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8637 = _T_8635 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8638 = _T_8634 | _T_8637; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8639 = _T_8638 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8641 = _T_8639 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8651 = _T_4525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8652 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8654 = _T_8652 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8655 = _T_8651 | _T_8654; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8656 = _T_8655 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8658 = _T_8656 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8668 = _T_4526 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8669 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 760:102]
  wire  _T_8671 = _T_8669 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8672 = _T_8668 | _T_8671; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8673 = _T_8672 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8675 = _T_8673 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8685 = _T_4495 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8688 = _T_8142 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8689 = _T_8685 | _T_8688; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8690 = _T_8689 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8692 = _T_8690 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8702 = _T_4496 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8705 = _T_8159 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8706 = _T_8702 | _T_8705; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8707 = _T_8706 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8709 = _T_8707 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8719 = _T_4497 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8722 = _T_8176 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8723 = _T_8719 | _T_8722; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8724 = _T_8723 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8726 = _T_8724 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8736 = _T_4498 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8739 = _T_8193 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8740 = _T_8736 | _T_8739; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8741 = _T_8740 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8743 = _T_8741 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8753 = _T_4499 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8756 = _T_8210 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8757 = _T_8753 | _T_8756; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8758 = _T_8757 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8760 = _T_8758 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8770 = _T_4500 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8773 = _T_8227 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8774 = _T_8770 | _T_8773; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8775 = _T_8774 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8777 = _T_8775 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8787 = _T_4501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8790 = _T_8244 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8791 = _T_8787 | _T_8790; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8792 = _T_8791 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8794 = _T_8792 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8804 = _T_4502 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8807 = _T_8261 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8808 = _T_8804 | _T_8807; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8809 = _T_8808 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8811 = _T_8809 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8821 = _T_4503 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8824 = _T_8278 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8825 = _T_8821 | _T_8824; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8826 = _T_8825 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8828 = _T_8826 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8838 = _T_4504 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8841 = _T_8295 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8842 = _T_8838 | _T_8841; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8843 = _T_8842 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8845 = _T_8843 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8855 = _T_4505 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8858 = _T_8312 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8859 = _T_8855 | _T_8858; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8860 = _T_8859 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8862 = _T_8860 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8872 = _T_4506 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8875 = _T_8329 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8876 = _T_8872 | _T_8875; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8877 = _T_8876 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8879 = _T_8877 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8889 = _T_4507 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8892 = _T_8346 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8893 = _T_8889 | _T_8892; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8894 = _T_8893 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8896 = _T_8894 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8906 = _T_4508 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8909 = _T_8363 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8910 = _T_8906 | _T_8909; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8911 = _T_8910 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8913 = _T_8911 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8923 = _T_4509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8926 = _T_8380 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8927 = _T_8923 | _T_8926; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8928 = _T_8927 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8930 = _T_8928 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8940 = _T_4510 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8943 = _T_8397 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8944 = _T_8940 | _T_8943; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8945 = _T_8944 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8947 = _T_8945 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8957 = _T_4511 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8960 = _T_8414 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8961 = _T_8957 | _T_8960; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8962 = _T_8961 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8964 = _T_8962 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8974 = _T_4512 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8977 = _T_8431 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8978 = _T_8974 | _T_8977; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8979 = _T_8978 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8981 = _T_8979 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_8991 = _T_4513 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_8994 = _T_8448 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_8995 = _T_8991 | _T_8994; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_8996 = _T_8995 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_8998 = _T_8996 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9008 = _T_4514 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9011 = _T_8465 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9012 = _T_9008 | _T_9011; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9013 = _T_9012 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9015 = _T_9013 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9025 = _T_4515 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9028 = _T_8482 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9029 = _T_9025 | _T_9028; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9030 = _T_9029 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9032 = _T_9030 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9042 = _T_4516 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9045 = _T_8499 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9046 = _T_9042 | _T_9045; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9047 = _T_9046 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9049 = _T_9047 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9059 = _T_4517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9062 = _T_8516 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9063 = _T_9059 | _T_9062; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9064 = _T_9063 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9066 = _T_9064 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9076 = _T_4518 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9079 = _T_8533 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9080 = _T_9076 | _T_9079; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9081 = _T_9080 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9083 = _T_9081 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9093 = _T_4519 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9096 = _T_8550 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9097 = _T_9093 | _T_9096; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9098 = _T_9097 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9100 = _T_9098 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9110 = _T_4520 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9113 = _T_8567 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9114 = _T_9110 | _T_9113; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9115 = _T_9114 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9117 = _T_9115 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9127 = _T_4521 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9130 = _T_8584 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9131 = _T_9127 | _T_9130; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9132 = _T_9131 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9134 = _T_9132 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9144 = _T_4522 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9147 = _T_8601 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9148 = _T_9144 | _T_9147; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9149 = _T_9148 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9151 = _T_9149 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9161 = _T_4523 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9164 = _T_8618 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9165 = _T_9161 | _T_9164; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9166 = _T_9165 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9168 = _T_9166 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9178 = _T_4524 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9181 = _T_8635 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9182 = _T_9178 | _T_9181; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9183 = _T_9182 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9185 = _T_9183 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9195 = _T_4525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9198 = _T_8652 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9199 = _T_9195 | _T_9198; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9200 = _T_9199 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9202 = _T_9200 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_9212 = _T_4526 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 760:59]
  wire  _T_9215 = _T_8669 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 760:124]
  wire  _T_9216 = _T_9212 | _T_9215; // @[el2_ifu_mem_ctl.scala 760:81]
  wire  _T_9217 = _T_9216 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 760:147]
  wire  _T_9219 = _T_9217 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 760:165]
  wire  _T_10021 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 815:63]
  wire  _T_10022 = _T_10021 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 815:85]
  wire [1:0] _T_10024 = _T_10022 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10031; // @[el2_ifu_mem_ctl.scala 820:57]
  reg  _T_10032; // @[el2_ifu_mem_ctl.scala 821:56]
  reg  _T_10033; // @[el2_ifu_mem_ctl.scala 822:59]
  wire  _T_10034 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 823:80]
  wire  _T_10035 = ifu_bus_arvalid_ff & _T_10034; // @[el2_ifu_mem_ctl.scala 823:78]
  wire  _T_10036 = _T_10035 & miss_pending; // @[el2_ifu_mem_ctl.scala 823:100]
  reg  _T_10037; // @[el2_ifu_mem_ctl.scala 823:58]
  reg  _T_10038; // @[el2_ifu_mem_ctl.scala 824:58]
  wire  _T_10041 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 831:71]
  wire  _T_10043 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 831:124]
  wire  _T_10045 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 832:50]
  wire  _T_10047 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 832:103]
  wire [3:0] _T_10050 = {_T_10041,_T_10043,_T_10045,_T_10047}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 834:53]
  reg  _T_10061; // @[Reg.scala 27:20]
  rvecc_encode m1 ( // @[el2_ifu_mem_ctl.scala 635:18]
    .io_din(m1_io_din),
    .io_ecc_out(m1_io_ecc_out)
  );
  rvecc_encode m2 ( // @[el2_ifu_mem_ctl.scala 637:18]
    .io_din(m2_io_din),
    .io_ecc_out(m2_io_ecc_out)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 327:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 326:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 191:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3588; // @[el2_ifu_mem_ctl.scala 701:21]
  assign io_ifu_pmu_ic_miss = _T_10031; // @[el2_ifu_mem_ctl.scala 820:22]
  assign io_ifu_pmu_ic_hit = _T_10032; // @[el2_ifu_mem_ctl.scala 821:21]
  assign io_ifu_pmu_bus_error = _T_10033; // @[el2_ifu_mem_ctl.scala 822:24]
  assign io_ifu_pmu_bus_busy = _T_10037; // @[el2_ifu_mem_ctl.scala 823:23]
  assign io_ifu_pmu_bus_trxn = _T_10038; // @[el2_ifu_mem_ctl.scala 824:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 141:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 140:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 135:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 139:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 150:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 145:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 143:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 136:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 132:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 133:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 142:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 151:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 559:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2572; // @[el2_ifu_mem_ctl.scala 560:19]
  assign io_ifu_axi_araddr = _T_2574 & _T_2576; // @[el2_ifu_mem_ctl.scala 561:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 564:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 147:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 562:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 565:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 563:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 566:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 660:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 658:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 662:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 653:20]
  assign io_iccm_ready = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 629:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 336:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3574; // @[el2_ifu_mem_ctl.scala 700:15]
  assign io_ic_rd_en = _T_3566 | _T_3571; // @[el2_ifu_mem_ctl.scala 691:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 343:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 343:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 344:23]
  assign io_ifu_ic_debug_rd_data = _T_1209; // @[el2_ifu_mem_ctl.scala 352:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 827:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 829:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 830:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 828:25]
  assign io_ic_debug_way = _T_10050[1:0]; // @[el2_ifu_mem_ctl.scala 831:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10024; // @[el2_ifu_mem_ctl.scala 815:19]
  assign io_iccm_rw_addr = _T_2720[14:0]; // @[el2_ifu_mem_ctl.scala 664:19]
  assign io_iccm_wren = _T_2679 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 631:16]
  assign io_iccm_rden = _T_2683 | _T_2684; // @[el2_ifu_mem_ctl.scala 632:16]
  assign io_iccm_wr_data = _T_2695 ? _T_2696 : _T_2703; // @[el2_ifu_mem_ctl.scala 641:19]
  assign io_iccm_wr_size = _T_2689 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 634:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 288:15]
  assign io_ic_access_fault_f = _T_2457 & _T_317; // @[el2_ifu_mem_ctl.scala 384:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1271; // @[el2_ifu_mem_ctl.scala 385:29]
  assign io_iccm_rd_ecc_single_err = _T_3511 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 677:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 678:29]
  assign io_ic_error_start = _T_1197 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 346:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 190:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 189:24]
  assign io_ic_fetch_val_f = {_T_1279,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 388:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 381:16]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[el2_ifu_mem_ctl.scala 378:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 379:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10061; // @[el2_ifu_mem_ctl.scala 838:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2462; // @[el2_ifu_mem_ctl.scala 478:27]
  assign io_iccm_correction_state = _T_2490 ? 1'h0 : _GEN_60; // @[el2_ifu_mem_ctl.scala 513:28 el2_ifu_mem_ctl.scala 526:32 el2_ifu_mem_ctl.scala 533:32 el2_ifu_mem_ctl.scala 540:32]
  assign m1_io_din = io_dma_mem_wdata[31:0]; // @[el2_ifu_mem_ctl.scala 636:13]
  assign m2_io_din = io_dma_mem_wdata[63:32]; // @[el2_ifu_mem_ctl.scala 638:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1209 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_443[6:0];
  _RAND_444 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_446[2:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_449[0:0];
  _RAND_450 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_450[38:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_453[2:0];
  _RAND_454 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_454[0:0];
  _RAND_455 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_455[63:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_456[13:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_458[13:0];
  _RAND_459 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_459[6:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way_status_new_ff = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  ic_valid_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10031 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10032 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10033 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10037 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10038 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_10061 = _RAND_469[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_3622) begin
      way_status_out_0 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_3627) begin
      way_status_out_1 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_3632) begin
      way_status_out_2 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_3637) begin
      way_status_out_3 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_3642) begin
      way_status_out_4 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_3647) begin
      way_status_out_5 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_3652) begin
      way_status_out_6 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_3657) begin
      way_status_out_7 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_3662) begin
      way_status_out_8 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_3667) begin
      way_status_out_9 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_3672) begin
      way_status_out_10 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_3677) begin
      way_status_out_11 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_3682) begin
      way_status_out_12 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_3687) begin
      way_status_out_13 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_3692) begin
      way_status_out_14 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_3697) begin
      way_status_out_15 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_3702) begin
      way_status_out_16 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_3707) begin
      way_status_out_17 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_3712) begin
      way_status_out_18 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_3717) begin
      way_status_out_19 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_3722) begin
      way_status_out_20 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_3727) begin
      way_status_out_21 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_3732) begin
      way_status_out_22 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_3737) begin
      way_status_out_23 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_3742) begin
      way_status_out_24 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_3747) begin
      way_status_out_25 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_3752) begin
      way_status_out_26 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_3757) begin
      way_status_out_27 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_3762) begin
      way_status_out_28 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_3767) begin
      way_status_out_29 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_3772) begin
      way_status_out_30 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_3777) begin
      way_status_out_31 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_3782) begin
      way_status_out_32 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_3787) begin
      way_status_out_33 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_3792) begin
      way_status_out_34 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_3797) begin
      way_status_out_35 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_3802) begin
      way_status_out_36 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_3807) begin
      way_status_out_37 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_3812) begin
      way_status_out_38 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_3817) begin
      way_status_out_39 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_3822) begin
      way_status_out_40 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_3827) begin
      way_status_out_41 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_3832) begin
      way_status_out_42 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_3837) begin
      way_status_out_43 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_3842) begin
      way_status_out_44 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_3847) begin
      way_status_out_45 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_3852) begin
      way_status_out_46 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_3857) begin
      way_status_out_47 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_3862) begin
      way_status_out_48 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_3867) begin
      way_status_out_49 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_3872) begin
      way_status_out_50 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_3877) begin
      way_status_out_51 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_3882) begin
      way_status_out_52 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_3887) begin
      way_status_out_53 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_3892) begin
      way_status_out_54 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_3897) begin
      way_status_out_55 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_3902) begin
      way_status_out_56 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_3907) begin
      way_status_out_57 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_3912) begin
      way_status_out_58 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_3917) begin
      way_status_out_59 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_3922) begin
      way_status_out_60 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_3927) begin
      way_status_out_61 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_3932) begin
      way_status_out_62 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_3937) begin
      way_status_out_63 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_3942) begin
      way_status_out_64 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_3947) begin
      way_status_out_65 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_3952) begin
      way_status_out_66 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_3957) begin
      way_status_out_67 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_3962) begin
      way_status_out_68 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_3967) begin
      way_status_out_69 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_3972) begin
      way_status_out_70 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_3977) begin
      way_status_out_71 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_3982) begin
      way_status_out_72 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_3987) begin
      way_status_out_73 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_3992) begin
      way_status_out_74 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_3997) begin
      way_status_out_75 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4002) begin
      way_status_out_76 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4007) begin
      way_status_out_77 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4012) begin
      way_status_out_78 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4017) begin
      way_status_out_79 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4022) begin
      way_status_out_80 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4027) begin
      way_status_out_81 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_82 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_83 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4042) begin
      way_status_out_84 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4047) begin
      way_status_out_85 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4052) begin
      way_status_out_86 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4057) begin
      way_status_out_87 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4062) begin
      way_status_out_88 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4067) begin
      way_status_out_89 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4072) begin
      way_status_out_90 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4077) begin
      way_status_out_91 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4082) begin
      way_status_out_92 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4087) begin
      way_status_out_93 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4092) begin
      way_status_out_94 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4097) begin
      way_status_out_95 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4102) begin
      way_status_out_96 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4107) begin
      way_status_out_97 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4112) begin
      way_status_out_98 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4117) begin
      way_status_out_99 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4122) begin
      way_status_out_100 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4127) begin
      way_status_out_101 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4132) begin
      way_status_out_102 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4137) begin
      way_status_out_103 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4142) begin
      way_status_out_104 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4147) begin
      way_status_out_105 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4152) begin
      way_status_out_106 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4157) begin
      way_status_out_107 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4162) begin
      way_status_out_108 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4167) begin
      way_status_out_109 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4172) begin
      way_status_out_110 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4177) begin
      way_status_out_111 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4182) begin
      way_status_out_112 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4187) begin
      way_status_out_113 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4192) begin
      way_status_out_114 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4197) begin
      way_status_out_115 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4202) begin
      way_status_out_116 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4207) begin
      way_status_out_117 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4212) begin
      way_status_out_118 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4217) begin
      way_status_out_119 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4222) begin
      way_status_out_120 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4227) begin
      way_status_out_121 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4232) begin
      way_status_out_122 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4237) begin
      way_status_out_123 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4242) begin
      way_status_out_124 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4247) begin
      way_status_out_125 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4252) begin
      way_status_out_126 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4257) begin
      way_status_out_127 <= way_status_new_ff;
    end
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2615) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2611;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5428) begin
      ic_tag_valid_out_1_0 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5445) begin
      ic_tag_valid_out_1_1 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5462) begin
      ic_tag_valid_out_1_2 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5479) begin
      ic_tag_valid_out_1_3 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5496) begin
      ic_tag_valid_out_1_4 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5513) begin
      ic_tag_valid_out_1_5 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5530) begin
      ic_tag_valid_out_1_6 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5547) begin
      ic_tag_valid_out_1_7 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5564) begin
      ic_tag_valid_out_1_8 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5581) begin
      ic_tag_valid_out_1_9 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5598) begin
      ic_tag_valid_out_1_10 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5615) begin
      ic_tag_valid_out_1_11 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5632) begin
      ic_tag_valid_out_1_12 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5649) begin
      ic_tag_valid_out_1_13 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5666) begin
      ic_tag_valid_out_1_14 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5683) begin
      ic_tag_valid_out_1_15 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5700) begin
      ic_tag_valid_out_1_16 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5717) begin
      ic_tag_valid_out_1_17 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5734) begin
      ic_tag_valid_out_1_18 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5751) begin
      ic_tag_valid_out_1_19 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5768) begin
      ic_tag_valid_out_1_20 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5785) begin
      ic_tag_valid_out_1_21 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5802) begin
      ic_tag_valid_out_1_22 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5819) begin
      ic_tag_valid_out_1_23 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5836) begin
      ic_tag_valid_out_1_24 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5853) begin
      ic_tag_valid_out_1_25 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5870) begin
      ic_tag_valid_out_1_26 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5887) begin
      ic_tag_valid_out_1_27 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_5904) begin
      ic_tag_valid_out_1_28 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_5921) begin
      ic_tag_valid_out_1_29 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_5938) begin
      ic_tag_valid_out_1_30 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_5955) begin
      ic_tag_valid_out_1_31 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6516) begin
      ic_tag_valid_out_1_32 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6533) begin
      ic_tag_valid_out_1_33 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6550) begin
      ic_tag_valid_out_1_34 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6567) begin
      ic_tag_valid_out_1_35 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6584) begin
      ic_tag_valid_out_1_36 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6601) begin
      ic_tag_valid_out_1_37 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6618) begin
      ic_tag_valid_out_1_38 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6635) begin
      ic_tag_valid_out_1_39 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6652) begin
      ic_tag_valid_out_1_40 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6669) begin
      ic_tag_valid_out_1_41 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6686) begin
      ic_tag_valid_out_1_42 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6703) begin
      ic_tag_valid_out_1_43 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6720) begin
      ic_tag_valid_out_1_44 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6737) begin
      ic_tag_valid_out_1_45 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6754) begin
      ic_tag_valid_out_1_46 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6771) begin
      ic_tag_valid_out_1_47 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6788) begin
      ic_tag_valid_out_1_48 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6805) begin
      ic_tag_valid_out_1_49 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6822) begin
      ic_tag_valid_out_1_50 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6839) begin
      ic_tag_valid_out_1_51 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6856) begin
      ic_tag_valid_out_1_52 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6873) begin
      ic_tag_valid_out_1_53 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6890) begin
      ic_tag_valid_out_1_54 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6907) begin
      ic_tag_valid_out_1_55 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6924) begin
      ic_tag_valid_out_1_56 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6941) begin
      ic_tag_valid_out_1_57 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6958) begin
      ic_tag_valid_out_1_58 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6975) begin
      ic_tag_valid_out_1_59 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6992) begin
      ic_tag_valid_out_1_60 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7009) begin
      ic_tag_valid_out_1_61 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7026) begin
      ic_tag_valid_out_1_62 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7043) begin
      ic_tag_valid_out_1_63 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7604) begin
      ic_tag_valid_out_1_64 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7621) begin
      ic_tag_valid_out_1_65 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7638) begin
      ic_tag_valid_out_1_66 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7655) begin
      ic_tag_valid_out_1_67 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7672) begin
      ic_tag_valid_out_1_68 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7689) begin
      ic_tag_valid_out_1_69 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7706) begin
      ic_tag_valid_out_1_70 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7723) begin
      ic_tag_valid_out_1_71 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7740) begin
      ic_tag_valid_out_1_72 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7757) begin
      ic_tag_valid_out_1_73 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7774) begin
      ic_tag_valid_out_1_74 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7791) begin
      ic_tag_valid_out_1_75 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7808) begin
      ic_tag_valid_out_1_76 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7825) begin
      ic_tag_valid_out_1_77 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7842) begin
      ic_tag_valid_out_1_78 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7859) begin
      ic_tag_valid_out_1_79 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7876) begin
      ic_tag_valid_out_1_80 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7893) begin
      ic_tag_valid_out_1_81 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7910) begin
      ic_tag_valid_out_1_82 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7927) begin
      ic_tag_valid_out_1_83 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7944) begin
      ic_tag_valid_out_1_84 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7961) begin
      ic_tag_valid_out_1_85 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7978) begin
      ic_tag_valid_out_1_86 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7995) begin
      ic_tag_valid_out_1_87 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8012) begin
      ic_tag_valid_out_1_88 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8029) begin
      ic_tag_valid_out_1_89 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8046) begin
      ic_tag_valid_out_1_90 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8063) begin
      ic_tag_valid_out_1_91 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8080) begin
      ic_tag_valid_out_1_92 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8097) begin
      ic_tag_valid_out_1_93 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8114) begin
      ic_tag_valid_out_1_94 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8131) begin
      ic_tag_valid_out_1_95 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8692) begin
      ic_tag_valid_out_1_96 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8709) begin
      ic_tag_valid_out_1_97 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8726) begin
      ic_tag_valid_out_1_98 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8743) begin
      ic_tag_valid_out_1_99 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8760) begin
      ic_tag_valid_out_1_100 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8777) begin
      ic_tag_valid_out_1_101 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8794) begin
      ic_tag_valid_out_1_102 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8811) begin
      ic_tag_valid_out_1_103 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8828) begin
      ic_tag_valid_out_1_104 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8845) begin
      ic_tag_valid_out_1_105 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8862) begin
      ic_tag_valid_out_1_106 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8879) begin
      ic_tag_valid_out_1_107 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8896) begin
      ic_tag_valid_out_1_108 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8913) begin
      ic_tag_valid_out_1_109 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8930) begin
      ic_tag_valid_out_1_110 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8947) begin
      ic_tag_valid_out_1_111 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8964) begin
      ic_tag_valid_out_1_112 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8981) begin
      ic_tag_valid_out_1_113 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8998) begin
      ic_tag_valid_out_1_114 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9015) begin
      ic_tag_valid_out_1_115 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9032) begin
      ic_tag_valid_out_1_116 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9049) begin
      ic_tag_valid_out_1_117 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9066) begin
      ic_tag_valid_out_1_118 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9083) begin
      ic_tag_valid_out_1_119 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9100) begin
      ic_tag_valid_out_1_120 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9117) begin
      ic_tag_valid_out_1_121 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9134) begin
      ic_tag_valid_out_1_122 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9151) begin
      ic_tag_valid_out_1_123 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9168) begin
      ic_tag_valid_out_1_124 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9185) begin
      ic_tag_valid_out_1_125 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9202) begin
      ic_tag_valid_out_1_126 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9219) begin
      ic_tag_valid_out_1_127 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_4884) begin
      ic_tag_valid_out_0_0 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_4901) begin
      ic_tag_valid_out_0_1 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_4918) begin
      ic_tag_valid_out_0_2 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_4935) begin
      ic_tag_valid_out_0_3 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_4952) begin
      ic_tag_valid_out_0_4 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_4969) begin
      ic_tag_valid_out_0_5 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_4986) begin
      ic_tag_valid_out_0_6 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5003) begin
      ic_tag_valid_out_0_7 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5020) begin
      ic_tag_valid_out_0_8 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5037) begin
      ic_tag_valid_out_0_9 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5054) begin
      ic_tag_valid_out_0_10 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5071) begin
      ic_tag_valid_out_0_11 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5088) begin
      ic_tag_valid_out_0_12 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5105) begin
      ic_tag_valid_out_0_13 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5122) begin
      ic_tag_valid_out_0_14 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5139) begin
      ic_tag_valid_out_0_15 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5156) begin
      ic_tag_valid_out_0_16 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5173) begin
      ic_tag_valid_out_0_17 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5190) begin
      ic_tag_valid_out_0_18 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5207) begin
      ic_tag_valid_out_0_19 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5224) begin
      ic_tag_valid_out_0_20 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5241) begin
      ic_tag_valid_out_0_21 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5258) begin
      ic_tag_valid_out_0_22 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5275) begin
      ic_tag_valid_out_0_23 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5292) begin
      ic_tag_valid_out_0_24 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5309) begin
      ic_tag_valid_out_0_25 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5326) begin
      ic_tag_valid_out_0_26 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5343) begin
      ic_tag_valid_out_0_27 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5360) begin
      ic_tag_valid_out_0_28 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5377) begin
      ic_tag_valid_out_0_29 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5394) begin
      ic_tag_valid_out_0_30 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5411) begin
      ic_tag_valid_out_0_31 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_5972) begin
      ic_tag_valid_out_0_32 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_5989) begin
      ic_tag_valid_out_0_33 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6006) begin
      ic_tag_valid_out_0_34 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6023) begin
      ic_tag_valid_out_0_35 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6040) begin
      ic_tag_valid_out_0_36 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6057) begin
      ic_tag_valid_out_0_37 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6074) begin
      ic_tag_valid_out_0_38 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6091) begin
      ic_tag_valid_out_0_39 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6108) begin
      ic_tag_valid_out_0_40 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6125) begin
      ic_tag_valid_out_0_41 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6142) begin
      ic_tag_valid_out_0_42 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6159) begin
      ic_tag_valid_out_0_43 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6176) begin
      ic_tag_valid_out_0_44 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6193) begin
      ic_tag_valid_out_0_45 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6210) begin
      ic_tag_valid_out_0_46 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6227) begin
      ic_tag_valid_out_0_47 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6244) begin
      ic_tag_valid_out_0_48 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6261) begin
      ic_tag_valid_out_0_49 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6278) begin
      ic_tag_valid_out_0_50 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6295) begin
      ic_tag_valid_out_0_51 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6312) begin
      ic_tag_valid_out_0_52 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6329) begin
      ic_tag_valid_out_0_53 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6346) begin
      ic_tag_valid_out_0_54 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6363) begin
      ic_tag_valid_out_0_55 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6380) begin
      ic_tag_valid_out_0_56 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6397) begin
      ic_tag_valid_out_0_57 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6414) begin
      ic_tag_valid_out_0_58 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6431) begin
      ic_tag_valid_out_0_59 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6448) begin
      ic_tag_valid_out_0_60 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6465) begin
      ic_tag_valid_out_0_61 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6482) begin
      ic_tag_valid_out_0_62 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6499) begin
      ic_tag_valid_out_0_63 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7060) begin
      ic_tag_valid_out_0_64 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7077) begin
      ic_tag_valid_out_0_65 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7094) begin
      ic_tag_valid_out_0_66 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7111) begin
      ic_tag_valid_out_0_67 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7128) begin
      ic_tag_valid_out_0_68 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7145) begin
      ic_tag_valid_out_0_69 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7162) begin
      ic_tag_valid_out_0_70 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7179) begin
      ic_tag_valid_out_0_71 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7196) begin
      ic_tag_valid_out_0_72 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7213) begin
      ic_tag_valid_out_0_73 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7230) begin
      ic_tag_valid_out_0_74 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7247) begin
      ic_tag_valid_out_0_75 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7264) begin
      ic_tag_valid_out_0_76 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7281) begin
      ic_tag_valid_out_0_77 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7298) begin
      ic_tag_valid_out_0_78 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7315) begin
      ic_tag_valid_out_0_79 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7332) begin
      ic_tag_valid_out_0_80 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7349) begin
      ic_tag_valid_out_0_81 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7366) begin
      ic_tag_valid_out_0_82 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7383) begin
      ic_tag_valid_out_0_83 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7400) begin
      ic_tag_valid_out_0_84 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7417) begin
      ic_tag_valid_out_0_85 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7434) begin
      ic_tag_valid_out_0_86 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7451) begin
      ic_tag_valid_out_0_87 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7468) begin
      ic_tag_valid_out_0_88 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7485) begin
      ic_tag_valid_out_0_89 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7502) begin
      ic_tag_valid_out_0_90 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7519) begin
      ic_tag_valid_out_0_91 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7536) begin
      ic_tag_valid_out_0_92 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7553) begin
      ic_tag_valid_out_0_93 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7570) begin
      ic_tag_valid_out_0_94 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7587) begin
      ic_tag_valid_out_0_95 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8148) begin
      ic_tag_valid_out_0_96 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8165) begin
      ic_tag_valid_out_0_97 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8182) begin
      ic_tag_valid_out_0_98 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8199) begin
      ic_tag_valid_out_0_99 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8216) begin
      ic_tag_valid_out_0_100 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8233) begin
      ic_tag_valid_out_0_101 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8250) begin
      ic_tag_valid_out_0_102 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8267) begin
      ic_tag_valid_out_0_103 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8284) begin
      ic_tag_valid_out_0_104 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8301) begin
      ic_tag_valid_out_0_105 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8318) begin
      ic_tag_valid_out_0_106 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8335) begin
      ic_tag_valid_out_0_107 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8352) begin
      ic_tag_valid_out_0_108 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8369) begin
      ic_tag_valid_out_0_109 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8386) begin
      ic_tag_valid_out_0_110 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8403) begin
      ic_tag_valid_out_0_111 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8420) begin
      ic_tag_valid_out_0_112 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8437) begin
      ic_tag_valid_out_0_113 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8454) begin
      ic_tag_valid_out_0_114 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8471) begin
      ic_tag_valid_out_0_115 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8488) begin
      ic_tag_valid_out_0_116 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8505) begin
      ic_tag_valid_out_0_117 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8522) begin
      ic_tag_valid_out_0_118 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8539) begin
      ic_tag_valid_out_0_119 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8556) begin
      ic_tag_valid_out_0_120 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8573) begin
      ic_tag_valid_out_0_121 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8590) begin
      ic_tag_valid_out_0_122 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8607) begin
      ic_tag_valid_out_0_123 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8624) begin
      ic_tag_valid_out_0_124 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8641) begin
      ic_tag_valid_out_0_125 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8658) begin
      ic_tag_valid_out_0_126 <= _T_4874;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8675) begin
      ic_tag_valid_out_0_127 <= _T_4874;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1209 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_1209 <= {{5'd0}, _T_1208};
      end else begin
        _T_1209 <= io_ic_debug_rd_data;
      end
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2564) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2639) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2683;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2465) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2467) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2477) begin
        perr_state <= 3'h0;
      end else if (_T_2480) begin
        if (_T_2482) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2486) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2490) begin
        err_stop_state <= 2'h1;
      end else if (_T_2495) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (_T_2518) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2522) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2539) begin
        if (_T_2543) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1368;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3597) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1408;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3532;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_2707;
    end else begin
      iccm_dma_rdata_temp <= _T_2708;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3528;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3597) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_3600) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_10009) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3600) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10061 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10061 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10031 <= 1'h0;
    end else begin
      _T_10031 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10032 <= 1'h0;
    end else begin
      _T_10032 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10033 <= 1'h0;
    end else begin
      _T_10033 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10037 <= 1'h0;
    end else begin
      _T_10037 <= _T_10036;
    end
    if (reset) begin
      _T_10038 <= 1'h0;
    end else begin
      _T_10038 <= bus_cmd_sent;
    end
  end
endmodule
