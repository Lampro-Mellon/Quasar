module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[el2_lib.scala 408:26]
  wire  clkhdr_CK; // @[el2_lib.scala 408:26]
  wire  clkhdr_EN; // @[el2_lib.scala 408:26]
  wire  clkhdr_SE; // @[el2_lib.scala 408:26]
  TEC_RV_ICG clkhdr ( // @[el2_lib.scala 408:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[el2_lib.scala 409:14]
  assign clkhdr_CK = io_clk; // @[el2_lib.scala 410:18]
  assign clkhdr_EN = io_en; // @[el2_lib.scala 411:18]
  assign clkhdr_SE = io_scan_mode; // @[el2_lib.scala 412:18]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  input         io_ifu_axi_arready,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  input         io_ifu_axi_rvalid,
  output        io_ifu_axi_rready,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [95:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [63:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_scan_mode; // @[el2_lib.scala 417:22]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 178:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 311:36]
  wire  _T_309 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 312:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_309; // @[el2_ifu_mem_ctl.scala 312:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 179:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 244:30]
  wire  _T_1 = _T | miss_pending; // @[el2_ifu_mem_ctl.scala 179:71]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 180:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 299:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 652:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 652:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_309}; // @[el2_ifu_mem_ctl.scala 655:91]
  wire [1:0] _T_3064 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 655:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 313:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 266:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 655:113]
  wire [1:0] _T_3065 = _T_3064 & _GEN_465; // @[el2_ifu_mem_ctl.scala 655:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 641:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 655:130]
  wire [1:0] _T_3066 = _T_3065 | _GEN_466; // @[el2_ifu_mem_ctl.scala 655:130]
  wire  _T_3067 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 655:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_3067}; // @[el2_ifu_mem_ctl.scala 655:152]
  wire [1:0] _T_3068 = _T_3066 & _GEN_467; // @[el2_ifu_mem_ctl.scala 655:152]
  wire [1:0] _T_3057 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 655:91]
  wire [1:0] _T_3058 = _T_3057 & _GEN_465; // @[el2_ifu_mem_ctl.scala 655:113]
  wire [1:0] _T_3059 = _T_3058 | _GEN_466; // @[el2_ifu_mem_ctl.scala 655:130]
  wire [1:0] _T_3061 = _T_3059 & _GEN_467; // @[el2_ifu_mem_ctl.scala 655:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3068,_T_3061}; // @[Cat.scala 29:58]
  wire  _T_3168 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3169 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3170 = _T_3168 ^ _T_3169; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3178 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3179 = ^_T_3178; // @[el2_lib.scala 301:83]
  wire  _T_3180 = io_iccm_rd_data_ecc[37] ^ _T_3179; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3187 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3195 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3187}; // @[el2_lib.scala 301:103]
  wire  _T_3196 = ^_T_3195; // @[el2_lib.scala 301:110]
  wire  _T_3197 = io_iccm_rd_data_ecc[36] ^ _T_3196; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3204 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3212 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3204}; // @[el2_lib.scala 301:130]
  wire  _T_3213 = ^_T_3212; // @[el2_lib.scala 301:137]
  wire  _T_3214 = io_iccm_rd_data_ecc[35] ^ _T_3213; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3223 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3232 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3223}; // @[el2_lib.scala 301:157]
  wire  _T_3233 = ^_T_3232; // @[el2_lib.scala 301:164]
  wire  _T_3234 = io_iccm_rd_data_ecc[34] ^ _T_3233; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3243 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3252 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3243}; // @[el2_lib.scala 301:184]
  wire  _T_3253 = ^_T_3252; // @[el2_lib.scala 301:191]
  wire  _T_3254 = io_iccm_rd_data_ecc[33] ^ _T_3253; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3263 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3272 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3263}; // @[el2_lib.scala 301:211]
  wire  _T_3273 = ^_T_3272; // @[el2_lib.scala 301:218]
  wire  _T_3274 = io_iccm_rd_data_ecc[32] ^ _T_3273; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3280 = {_T_3170,_T_3180,_T_3197,_T_3214,_T_3234,_T_3254,_T_3274}; // @[Cat.scala 29:58]
  wire  _T_3281 = _T_3280 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3282 = iccm_ecc_word_enable[0] & _T_3281; // @[el2_lib.scala 302:32]
  wire  _T_3284 = _T_3282 & _T_3280[6]; // @[el2_lib.scala 302:53]
  wire  _T_3553 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3554 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3555 = _T_3553 ^ _T_3554; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3563 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3564 = ^_T_3563; // @[el2_lib.scala 301:83]
  wire  _T_3565 = io_iccm_rd_data_ecc[76] ^ _T_3564; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3572 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3580 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3572}; // @[el2_lib.scala 301:103]
  wire  _T_3581 = ^_T_3580; // @[el2_lib.scala 301:110]
  wire  _T_3582 = io_iccm_rd_data_ecc[75] ^ _T_3581; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3589 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3597 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3589}; // @[el2_lib.scala 301:130]
  wire  _T_3598 = ^_T_3597; // @[el2_lib.scala 301:137]
  wire  _T_3599 = io_iccm_rd_data_ecc[74] ^ _T_3598; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3608 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3617 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3608}; // @[el2_lib.scala 301:157]
  wire  _T_3618 = ^_T_3617; // @[el2_lib.scala 301:164]
  wire  _T_3619 = io_iccm_rd_data_ecc[73] ^ _T_3618; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3628 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3637 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3628}; // @[el2_lib.scala 301:184]
  wire  _T_3638 = ^_T_3637; // @[el2_lib.scala 301:191]
  wire  _T_3639 = io_iccm_rd_data_ecc[72] ^ _T_3638; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3648 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3657 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3648}; // @[el2_lib.scala 301:211]
  wire  _T_3658 = ^_T_3657; // @[el2_lib.scala 301:218]
  wire  _T_3659 = io_iccm_rd_data_ecc[71] ^ _T_3658; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3665 = {_T_3555,_T_3565,_T_3582,_T_3599,_T_3619,_T_3639,_T_3659}; // @[Cat.scala 29:58]
  wire  _T_3666 = _T_3665 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3667 = iccm_ecc_word_enable[1] & _T_3666; // @[el2_lib.scala 302:32]
  wire  _T_3669 = _T_3667 & _T_3665[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3284,_T_3669}; // @[Cat.scala 29:58]
  wire  _T_4 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 183:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 619:51]
  wire  _T_7 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 184:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_8 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 185:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 465:34]
  wire  _T_9 = iccm_correct_ecc | _T_8; // @[el2_ifu_mem_ctl.scala 185:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_10 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 185:90]
  wire  _T_11 = _T_9 | _T_10; // @[el2_ifu_mem_ctl.scala 185:72]
  wire  _T_2435 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2440 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2460 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 515:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 381:42]
  wire  _T_2462 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 515:79]
  wire  _T_2463 = _T_2460 | _T_2462; // @[el2_ifu_mem_ctl.scala 515:56]
  wire  _T_2464 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 515:122]
  wire  _T_2465 = ~_T_2464; // @[el2_ifu_mem_ctl.scala 515:101]
  wire  _T_2466 = _T_2463 & _T_2465; // @[el2_ifu_mem_ctl.scala 515:99]
  wire  _T_2467 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2481 = io_ifu_fetch_val[0] & _T_309; // @[el2_ifu_mem_ctl.scala 522:45]
  wire  _T_2482 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 522:69]
  wire  _T_2483 = _T_2481 & _T_2482; // @[el2_ifu_mem_ctl.scala 522:67]
  wire  _T_2484 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_2467 ? _T_2483 : _T_2484; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2440 ? _T_2466 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2435 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_12 = _T_11 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 185:112]
  wire  _T_14 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 186:44]
  wire  _T_15 = _T_14 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 186:65]
  wire  _T_219 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 274:37]
  wire  _T_220 = ~_T_219; // @[el2_ifu_mem_ctl.scala 274:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 687:53]
  wire  _T_221 = _T_220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 274:41]
  wire  _T_199 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 265:48]
  wire  _T_200 = ifc_fetch_req_f & _T_199; // @[el2_ifu_mem_ctl.scala 265:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 315:42]
  wire  _T_201 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 265:69]
  wire  fetch_req_icache_f = _T_200 & _T_201; // @[el2_ifu_mem_ctl.scala 265:67]
  wire  _T_222 = _T_221 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 274:59]
  wire  _T_223 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 274:82]
  wire  _T_224 = _T_222 & _T_223; // @[el2_ifu_mem_ctl.scala 274:80]
  wire  ic_act_miss_f = _T_224 & _T_201; // @[el2_ifu_mem_ctl.scala 274:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 535:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 576:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 603:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 301:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 584:56]
  wire  _T_2584 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 601:69]
  wire  _T_2585 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 601:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2584 : _T_2585; // @[el2_ifu_mem_ctl.scala 601:28]
  wire  _T_2531 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 580:68]
  wire  _T_2532 = ic_act_miss_f | _T_2531; // @[el2_ifu_mem_ctl.scala 580:48]
  wire  bus_reset_data_beat_cnt = _T_2532 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 580:91]
  wire  _T_2528 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 579:50]
  wire  _T_2529 = bus_ifu_wr_en_ff & _T_2528; // @[el2_ifu_mem_ctl.scala 579:48]
  wire  _T_2530 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 579:72]
  wire  bus_inc_data_beat_cnt = _T_2529 & _T_2530; // @[el2_ifu_mem_ctl.scala 579:70]
  wire [2:0] _T_2536 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 583:115]
  wire [2:0] _T_2538 = bus_inc_data_beat_cnt ? _T_2536 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2533 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 581:32]
  wire  _T_2534 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 581:57]
  wire  bus_hold_data_beat_cnt = _T_2533 & _T_2534; // @[el2_ifu_mem_ctl.scala 581:55]
  wire [2:0] _T_2539 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2538 | _T_2539; // @[Mux.scala 27:72]
  wire  _T_16 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 186:111]
  wire  _T_17 = _T_15 & _T_16; // @[el2_ifu_mem_ctl.scala 186:85]
  wire  _T_18 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 187:39]
  wire  _T_26 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_28 = ic_act_miss_f & _T_309; // @[el2_ifu_mem_ctl.scala 193:43]
  wire [2:0] _T_30 = _T_28 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 193:27]
  wire  _T_33 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 417:45]
  wire  _T_2100 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 438:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 394:60]
  wire  _T_2131 = _T_2100 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2104 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2132 = _T_2104 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2139 = _T_2131 | _T_2132; // @[Mux.scala 27:72]
  wire  _T_2108 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2133 = _T_2108 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2140 = _T_2139 | _T_2133; // @[Mux.scala 27:72]
  wire  _T_2112 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2134 = _T_2112 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2141 = _T_2140 | _T_2134; // @[Mux.scala 27:72]
  wire  _T_2116 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2135 = _T_2116 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2142 = _T_2141 | _T_2135; // @[Mux.scala 27:72]
  wire  _T_2120 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2136 = _T_2120 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2143 = _T_2142 | _T_2136; // @[Mux.scala 27:72]
  wire  _T_2124 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2137 = _T_2124 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2144 = _T_2143 | _T_2137; // @[Mux.scala 27:72]
  wire  _T_2128 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2138 = _T_2128 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2144 | _T_2138; // @[Mux.scala 27:72]
  wire  _T_2186 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 440:69]
  wire  _T_2187 = ic_miss_buff_data_valid_bypass_index & _T_2186; // @[el2_ifu_mem_ctl.scala 440:67]
  wire  _T_2189 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 440:91]
  wire  _T_2190 = _T_2187 & _T_2189; // @[el2_ifu_mem_ctl.scala 440:89]
  wire  _T_2195 = _T_2187 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 441:65]
  wire  _T_2196 = _T_2190 | _T_2195; // @[el2_ifu_mem_ctl.scala 440:112]
  wire  _T_2198 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 442:43]
  wire  _T_2201 = _T_2198 & _T_2189; // @[el2_ifu_mem_ctl.scala 442:65]
  wire  _T_2202 = _T_2196 | _T_2201; // @[el2_ifu_mem_ctl.scala 441:88]
  wire  _T_2206 = _T_2198 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 443:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 420:75]
  wire  _T_2146 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2170 = _T_2146 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2149 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2171 = _T_2149 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2178 = _T_2170 | _T_2171; // @[Mux.scala 27:72]
  wire  _T_2152 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2172 = _T_2152 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2179 = _T_2178 | _T_2172; // @[Mux.scala 27:72]
  wire  _T_2155 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2173 = _T_2155 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2180 = _T_2179 | _T_2173; // @[Mux.scala 27:72]
  wire  _T_2158 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2174 = _T_2158 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2181 = _T_2180 | _T_2174; // @[Mux.scala 27:72]
  wire  _T_2161 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2175 = _T_2161 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2182 = _T_2181 | _T_2175; // @[Mux.scala 27:72]
  wire  _T_2164 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2176 = _T_2164 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2183 = _T_2182 | _T_2176; // @[Mux.scala 27:72]
  wire  _T_2167 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2177 = _T_2167 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2183 | _T_2177; // @[Mux.scala 27:72]
  wire  _T_2207 = _T_2206 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 443:87]
  wire  _T_2208 = _T_2202 | _T_2207; // @[el2_ifu_mem_ctl.scala 442:88]
  wire  _T_2218 = _T_2190 & _T_2128; // @[el2_ifu_mem_ctl.scala 444:87]
  wire  miss_buff_hit_unq_f = _T_2208 | _T_2218; // @[el2_ifu_mem_ctl.scala 443:131]
  wire  _T_2233 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 449:55]
  wire  _T_2234 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 449:87]
  wire  _T_2235 = _T_2233 | _T_2234; // @[el2_ifu_mem_ctl.scala 449:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2235; // @[el2_ifu_mem_ctl.scala 449:41]
  wire  _T_2219 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 446:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 302:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 437:51]
  wire  _T_2220 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 446:68]
  wire  _T_2221 = miss_buff_hit_unq_f & _T_2220; // @[el2_ifu_mem_ctl.scala 446:66]
  wire  stream_hit_f = _T_2219 & _T_2221; // @[el2_ifu_mem_ctl.scala 446:43]
  wire  _T_207 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 269:35]
  wire  _T_208 = _T_207 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 269:52]
  wire  ic_byp_hit_f = _T_208 & miss_pending; // @[el2_ifu_mem_ctl.scala 269:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 586:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 613:35]
  wire  _T_34 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 196:112]
  wire  _T_35 = last_data_recieved_ff | _T_34; // @[el2_ifu_mem_ctl.scala 196:92]
  wire  _T_36 = ic_byp_hit_f & _T_35; // @[el2_ifu_mem_ctl.scala 196:66]
  wire  _T_37 = _T_36 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 196:126]
  wire  _T_38 = io_dec_tlu_force_halt | _T_37; // @[el2_ifu_mem_ctl.scala 196:51]
  wire  _T_40 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 197:30]
  wire  _T_41 = ic_byp_hit_f & _T_40; // @[el2_ifu_mem_ctl.scala 197:27]
  wire  _T_42 = _T_41 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 197:53]
  wire  _T_44 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 198:16]
  wire  _T_46 = _T_44 & _T_309; // @[el2_ifu_mem_ctl.scala 198:30]
  wire  _T_48 = _T_46 & _T_34; // @[el2_ifu_mem_ctl.scala 198:52]
  wire  _T_49 = _T_48 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 198:85]
  wire  _T_52 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 199:51]
  wire  _T_53 = _T_34 & _T_52; // @[el2_ifu_mem_ctl.scala 199:49]
  wire  _T_55 = ic_byp_hit_f | bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 200:34]
  wire  _T_57 = _T_55 & _T_309; // @[el2_ifu_mem_ctl.scala 200:54]
  wire  _T_59 = ~_T_34; // @[el2_ifu_mem_ctl.scala 200:78]
  wire  _T_60 = _T_57 & _T_59; // @[el2_ifu_mem_ctl.scala 200:76]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 189:52]
  wire  _T_61 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 200:112]
  wire  _T_62 = _T_60 & _T_61; // @[el2_ifu_mem_ctl.scala 200:110]
  wire  _T_64 = _T_62 & _T_52; // @[el2_ifu_mem_ctl.scala 200:134]
  wire  _T_72 = _T_48 & _T_52; // @[el2_ifu_mem_ctl.scala 201:100]
  wire  _T_74 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 202:44]
  wire  _T_77 = _T_74 & _T_59; // @[el2_ifu_mem_ctl.scala 202:68]
  wire [2:0] _T_79 = _T_77 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 202:22]
  wire [2:0] _T_80 = _T_72 ? 3'h0 : _T_79; // @[el2_ifu_mem_ctl.scala 201:20]
  wire [2:0] _T_81 = _T_64 ? 3'h6 : _T_80; // @[el2_ifu_mem_ctl.scala 200:18]
  wire [2:0] _T_82 = _T_53 ? 3'h0 : _T_81; // @[el2_ifu_mem_ctl.scala 199:16]
  wire [2:0] _T_83 = _T_49 ? 3'h1 : _T_82; // @[el2_ifu_mem_ctl.scala 198:14]
  wire [2:0] _T_84 = _T_42 ? 3'h3 : _T_83; // @[el2_ifu_mem_ctl.scala 197:12]
  wire [2:0] _T_85 = _T_38 ? 3'h0 : _T_84; // @[el2_ifu_mem_ctl.scala 196:27]
  wire  _T_94 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_98 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2230 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 448:60]
  wire  _T_2231 = _T_2230 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 448:92]
  wire  stream_eol_f = _T_2231 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_100 = _T_74 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 210:72]
  wire  _T_103 = _T_100 & _T_59; // @[el2_ifu_mem_ctl.scala 210:87]
  wire  _T_105 = _T_103 & _T_2530; // @[el2_ifu_mem_ctl.scala 210:122]
  wire [2:0] _T_107 = _T_105 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 210:27]
  wire  _T_113 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_116 = io_exu_flush_final & _T_59; // @[el2_ifu_mem_ctl.scala 214:48]
  wire  _T_118 = _T_116 & _T_2530; // @[el2_ifu_mem_ctl.scala 214:82]
  wire [2:0] _T_120 = _T_118 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 214:27]
  wire  _T_124 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_228 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 275:28]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 275:42]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 275:60]
  wire  _T_231 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 275:94]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 275:81]
  wire  _T_235 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 276:39]
  wire  _T_236 = _T_232 & _T_235; // @[el2_ifu_mem_ctl.scala 275:111]
  wire  _T_238 = _T_236 & _T_52; // @[el2_ifu_mem_ctl.scala 276:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 329:51]
  wire  _T_239 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 276:116]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 276:114]
  wire  ic_miss_under_miss_f = _T_240 & _T_201; // @[el2_ifu_mem_ctl.scala 276:132]
  wire  _T_127 = ic_miss_under_miss_f & _T_59; // @[el2_ifu_mem_ctl.scala 218:50]
  wire  _T_129 = _T_127 & _T_2530; // @[el2_ifu_mem_ctl.scala 218:84]
  wire  _T_248 = _T_222 & _T_231; // @[el2_ifu_mem_ctl.scala 277:85]
  wire  _T_251 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 278:39]
  wire  _T_252 = _T_251 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 278:91]
  wire  ic_ignore_2nd_miss_f = _T_248 & _T_252; // @[el2_ifu_mem_ctl.scala 277:117]
  wire  _T_133 = ic_ignore_2nd_miss_f & _T_59; // @[el2_ifu_mem_ctl.scala 219:35]
  wire  _T_135 = _T_133 & _T_2530; // @[el2_ifu_mem_ctl.scala 219:69]
  wire [2:0] _T_137 = _T_135 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 219:12]
  wire [2:0] _T_138 = _T_129 ? 3'h5 : _T_137; // @[el2_ifu_mem_ctl.scala 218:27]
  wire  _T_143 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_146 = _T_34 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 224:12]
  wire [2:0] _T_147 = io_exu_flush_final ? _T_146 : 3'h1; // @[el2_ifu_mem_ctl.scala 223:62]
  wire [2:0] _T_148 = io_dec_tlu_force_halt ? 3'h0 : _T_147; // @[el2_ifu_mem_ctl.scala 223:27]
  wire  _T_152 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_156 = io_exu_flush_final ? _T_146 : 3'h0; // @[el2_ifu_mem_ctl.scala 228:62]
  wire [2:0] _T_157 = io_dec_tlu_force_halt ? 3'h0 : _T_156; // @[el2_ifu_mem_ctl.scala 228:27]
  wire [2:0] _GEN_0 = _T_152 ? _T_157 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_143 ? _T_148 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_124 ? _T_138 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_113 ? _T_120 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_98 ? _T_107 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_94 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_33 ? _T_85 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_26 ? _T_30 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_19 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 187:71]
  wire  _T_20 = _T_18 | _T_19; // @[el2_ifu_mem_ctl.scala 187:55]
  wire  _T_21 = uncacheable_miss_ff >> _T_20; // @[el2_ifu_mem_ctl.scala 187:26]
  wire  _T_23 = ~_T_21; // @[el2_ifu_mem_ctl.scala 187:5]
  wire  _T_24 = _T_17 & _T_23; // @[el2_ifu_mem_ctl.scala 186:116]
  wire  scnd_miss_req_in = _T_24 & _T_309; // @[el2_ifu_mem_ctl.scala 187:89]
  wire  _T_32 = ic_act_miss_f & _T_2530; // @[el2_ifu_mem_ctl.scala 194:38]
  wire  _T_86 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 203:46]
  wire  _T_87 = _T_86 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 203:67]
  wire  _T_88 = _T_87 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 203:82]
  wire  _T_90 = _T_88 | _T_34; // @[el2_ifu_mem_ctl.scala 203:105]
  wire  _T_92 = bus_ifu_wr_en_ff & _T_52; // @[el2_ifu_mem_ctl.scala 203:158]
  wire  _T_93 = _T_90 | _T_92; // @[el2_ifu_mem_ctl.scala 203:138]
  wire  _T_95 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 207:43]
  wire  _T_96 = _T_95 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:59]
  wire  _T_97 = _T_96 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 207:74]
  wire  _T_111 = _T_100 | _T_34; // @[el2_ifu_mem_ctl.scala 211:84]
  wire  _T_112 = _T_111 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 211:118]
  wire  _T_122 = io_exu_flush_final | _T_34; // @[el2_ifu_mem_ctl.scala 215:43]
  wire  _T_123 = _T_122 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 215:76]
  wire  _T_140 = _T_34 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 220:55]
  wire  _T_141 = _T_140 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 220:78]
  wire  _T_142 = _T_141 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 220:101]
  wire  _T_150 = _T_34 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 225:55]
  wire  _T_151 = _T_150 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _GEN_1 = _T_152 & _T_151; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_143 ? _T_151 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_124 ? _T_142 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_113 ? _T_123 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_98 ? _T_112 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_94 ? _T_97 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_33 ? _T_93 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_26 ? _T_32 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_166 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 245:95]
  wire  _T_167 = _T_2233 & _T_166; // @[el2_ifu_mem_ctl.scala 245:93]
  wire  crit_wd_byp_ok_ff = _T_2234 | _T_167; // @[el2_ifu_mem_ctl.scala 245:58]
  wire  _T_170 = miss_pending & _T_59; // @[el2_ifu_mem_ctl.scala 246:36]
  wire  _T_172 = _T_2233 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 246:106]
  wire  _T_173 = ~_T_172; // @[el2_ifu_mem_ctl.scala 246:72]
  wire  _T_174 = _T_170 & _T_173; // @[el2_ifu_mem_ctl.scala 246:70]
  wire  _T_176 = _T_2233 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 247:57]
  wire  _T_177 = ~_T_176; // @[el2_ifu_mem_ctl.scala 247:23]
  wire  _T_178 = _T_174 & _T_177; // @[el2_ifu_mem_ctl.scala 246:128]
  wire  _T_179 = _T_178 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 247:77]
  wire  _T_180 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 248:36]
  wire  _T_181 = miss_pending & _T_180; // @[el2_ifu_mem_ctl.scala 248:19]
  wire  sel_hold_imb = _T_179 | _T_181; // @[el2_ifu_mem_ctl.scala 247:93]
  wire  _T_183 = _T_18 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 250:57]
  wire  sel_hold_imb_scnd = _T_183 & _T_166; // @[el2_ifu_mem_ctl.scala 250:81]
  reg [6:0] _T_4981; // @[el2_ifu_mem_ctl.scala 717:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_4981[5:0]; // @[el2_ifu_mem_ctl.scala 716:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 713:121]
  wire  _T_4846 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4848 = _T_4846 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4337; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_4337[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4849 = _T_4848 & _GEN_473; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4842 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4844 = _T_4842 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4334; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_4334[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4845 = _T_4844 & _GEN_475; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4838 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4840 = _T_4838 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4331; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_4331[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4841 = _T_4840 & _GEN_477; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4834 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4836 = _T_4834 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4328; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_4328[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4837 = _T_4836 & _GEN_479; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4830 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4832 = _T_4830 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4325; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_4325[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4833 = _T_4832 & _GEN_481; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4826 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4828 = _T_4826 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4322; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_4322[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4829 = _T_4828 & _GEN_483; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4822 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4824 = _T_4822 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4319; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_4319[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4825 = _T_4824 & _GEN_485; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4818 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4820 = _T_4818 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4316; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_4316[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4821 = _T_4820 & _GEN_487; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4814 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4816 = _T_4814 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4313; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_4313[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4817 = _T_4816 & _GEN_489; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4810 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4812 = _T_4810 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4310; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_4310[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4813 = _T_4812 & _GEN_491; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [59:0] _T_4858 = {_T_4849,_T_4845,_T_4841,_T_4837,_T_4833,_T_4829,_T_4825,_T_4821,_T_4817,_T_4813}; // @[Cat.scala 29:58]
  wire  _T_4806 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4808 = _T_4806 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4307; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_4307[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4809 = _T_4808 & _GEN_493; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4802 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4804 = _T_4802 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4304; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_4304[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4805 = _T_4804 & _GEN_495; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4798 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4800 = _T_4798 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4301; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_4301[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4801 = _T_4800 & _GEN_497; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4794 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4796 = _T_4794 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4298; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_4298[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4797 = _T_4796 & _GEN_499; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4790 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4792 = _T_4790 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4295; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_4295[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4793 = _T_4792 & _GEN_501; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4786 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4788 = _T_4786 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4292; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_4292[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4789 = _T_4788 & _GEN_503; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4782 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4784 = _T_4782 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4289; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_4289[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4785 = _T_4784 & _GEN_505; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4778 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4780 = _T_4778 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4286; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_4286[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4781 = _T_4780 & _GEN_507; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4774 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4776 = _T_4774 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4283; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_4283[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4777 = _T_4776 & _GEN_509; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [113:0] _T_4867 = {_T_4858,_T_4809,_T_4805,_T_4801,_T_4797,_T_4793,_T_4789,_T_4785,_T_4781,_T_4777}; // @[Cat.scala 29:58]
  wire  _T_4770 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4772 = _T_4770 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4280; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_4280[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4773 = _T_4772 & _GEN_511; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4766 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4768 = _T_4766 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4277; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_4277[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4769 = _T_4768 & _GEN_513; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4762 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4764 = _T_4762 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4274; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_4274[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4765 = _T_4764 & _GEN_515; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4758 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4760 = _T_4758 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4271; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_4271[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4761 = _T_4760 & _GEN_517; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4754 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4756 = _T_4754 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4268; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_4268[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4757 = _T_4756 & _GEN_519; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4750 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4752 = _T_4750 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4265; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_4265[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4753 = _T_4752 & _GEN_521; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4746 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4748 = _T_4746 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4262; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_4262[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4749 = _T_4748 & _GEN_523; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4742 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4744 = _T_4742 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4259; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_4259[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4745 = _T_4744 & _GEN_525; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4738 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4740 = _T_4738 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4256; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_4256[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4741 = _T_4740 & _GEN_527; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [167:0] _T_4876 = {_T_4867,_T_4773,_T_4769,_T_4765,_T_4761,_T_4757,_T_4753,_T_4749,_T_4745,_T_4741}; // @[Cat.scala 29:58]
  wire  _T_4734 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4736 = _T_4734 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4253; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_4253[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4737 = _T_4736 & _GEN_529; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4730 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4732 = _T_4730 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4250; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_4250[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4733 = _T_4732 & _GEN_531; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4726 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4728 = _T_4726 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4247; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_4247[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4729 = _T_4728 & _GEN_533; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4722 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4724 = _T_4722 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4244; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_4244[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4725 = _T_4724 & _GEN_535; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4718 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4720 = _T_4718 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4241; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_4241[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4721 = _T_4720 & _GEN_537; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4714 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4716 = _T_4714 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4238; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_4238[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4717 = _T_4716 & _GEN_539; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4710 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4712 = _T_4710 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4235; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_4235[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4713 = _T_4712 & _GEN_541; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4706 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4708 = _T_4706 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4232; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_4232[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4709 = _T_4708 & _GEN_543; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4702 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4704 = _T_4702 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4229; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_4229[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4705 = _T_4704 & _GEN_545; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [221:0] _T_4885 = {_T_4876,_T_4737,_T_4733,_T_4729,_T_4725,_T_4721,_T_4717,_T_4713,_T_4709,_T_4705}; // @[Cat.scala 29:58]
  wire  _T_4698 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4700 = _T_4698 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4226; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_4226[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4701 = _T_4700 & _GEN_547; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4694 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4696 = _T_4694 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4223; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_4223[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4697 = _T_4696 & _GEN_549; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4690 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4692 = _T_4690 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4220; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_4220[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4693 = _T_4692 & _GEN_551; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4686 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4688 = _T_4686 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4217; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_4217[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4689 = _T_4688 & _GEN_553; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4682 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4684 = _T_4682 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4214; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_4214[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4685 = _T_4684 & _GEN_555; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4678 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4680 = _T_4678 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4211; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_4211[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4681 = _T_4680 & _GEN_557; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4674 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4676 = _T_4674 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4208; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_4208[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4677 = _T_4676 & _GEN_559; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4670 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4672 = _T_4670 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4205; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_4205[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4673 = _T_4672 & _GEN_561; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4666 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4668 = _T_4666 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4202; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_4202[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4669 = _T_4668 & _GEN_563; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [275:0] _T_4894 = {_T_4885,_T_4701,_T_4697,_T_4693,_T_4689,_T_4685,_T_4681,_T_4677,_T_4673,_T_4669}; // @[Cat.scala 29:58]
  wire  _T_4662 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4664 = _T_4662 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4199; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_4199[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4665 = _T_4664 & _GEN_565; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4658 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4660 = _T_4658 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4196; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_4196[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4661 = _T_4660 & _GEN_567; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4654 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4656 = _T_4654 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4193; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_4193[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4657 = _T_4656 & _GEN_569; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4650 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4652 = _T_4650 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4190; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_4190[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4653 = _T_4652 & _GEN_571; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4646 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4648 = _T_4646 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4187; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_4187[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4649 = _T_4648 & _GEN_573; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4642 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4644 = _T_4642 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4184; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_4184[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4645 = _T_4644 & _GEN_575; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4638 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4640 = _T_4638 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4181; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_4181[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4641 = _T_4640 & _GEN_577; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4634 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4636 = _T_4634 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4178; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_4178[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4637 = _T_4636 & _GEN_579; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4630 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4632 = _T_4630 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4175; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_4175[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4633 = _T_4632 & _GEN_581; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [329:0] _T_4903 = {_T_4894,_T_4665,_T_4661,_T_4657,_T_4653,_T_4649,_T_4645,_T_4641,_T_4637,_T_4633}; // @[Cat.scala 29:58]
  wire  _T_4626 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4628 = _T_4626 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4172; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_4172[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4629 = _T_4628 & _GEN_583; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4622 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4624 = _T_4622 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4169; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_4169[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4625 = _T_4624 & _GEN_585; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4618 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4620 = _T_4618 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4166; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_4166[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4621 = _T_4620 & _GEN_587; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4614 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4616 = _T_4614 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4163; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_4163[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4617 = _T_4616 & _GEN_589; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4610 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4612 = _T_4610 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4160; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_4160[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4613 = _T_4612 & _GEN_591; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4606 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4608 = _T_4606 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4157; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_4157[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4609 = _T_4608 & _GEN_593; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4602 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4604 = _T_4602 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4154; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_4154[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4605 = _T_4604 & _GEN_595; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4598 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4600 = _T_4598 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4151; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_4151[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4601 = _T_4600 & _GEN_597; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4594 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4596 = _T_4594 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4148; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_4148[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4597 = _T_4596 & _GEN_599; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [383:0] _T_4912 = {_T_4903,_T_4629,_T_4625,_T_4621,_T_4617,_T_4613,_T_4609,_T_4605,_T_4601,_T_4597}; // @[Cat.scala 29:58]
  wire  _T_4590 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4592 = _T_4590 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4145; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_4145[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4593 = _T_4592 & _GEN_600; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4586 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4588 = _T_4586 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4142; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_4142[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4589 = _T_4588 & _GEN_601; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4582 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4584 = _T_4582 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4139; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_4139[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4585 = _T_4584 & _GEN_602; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4578 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4580 = _T_4578 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4136; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_4136[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4581 = _T_4580 & _GEN_603; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4574 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4576 = _T_4574 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4133; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_4133[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4577 = _T_4576 & _GEN_604; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4570 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4572 = _T_4570 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4130; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_4130[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4573 = _T_4572 & _GEN_605; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4566 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4568 = _T_4566 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4127; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_4127[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4569 = _T_4568 & _GEN_606; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4562 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4564 = _T_4562 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4124; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_4124[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4565 = _T_4564 & _GEN_607; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4558 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4560 = _T_4558 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4121; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_4121[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4561 = _T_4560 & _GEN_608; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [437:0] _T_4921 = {_T_4912,_T_4593,_T_4589,_T_4585,_T_4581,_T_4577,_T_4573,_T_4569,_T_4565,_T_4561}; // @[Cat.scala 29:58]
  wire  _T_4554 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4556 = _T_4554 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4118; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_4118[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4557 = _T_4556 & _GEN_609; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4550 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4552 = _T_4550 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4115; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_4115[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4553 = _T_4552 & _GEN_610; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4546 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4548 = _T_4546 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4112; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_4112[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4549 = _T_4548 & _GEN_611; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4542 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4544 = _T_4542 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4109; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_4109[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4545 = _T_4544 & _GEN_612; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4538 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4540 = _T_4538 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4106; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_4106[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4541 = _T_4540 & _GEN_613; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4534 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4536 = _T_4534 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4103; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_4103[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4537 = _T_4536 & _GEN_614; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4530 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4532 = _T_4530 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4100; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_4100[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4533 = _T_4532 & _GEN_615; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4526 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4528 = _T_4526 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4097; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_4097[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4529 = _T_4528 & _GEN_616; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4522 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4524 = _T_4522 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4094; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_4094[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4525 = _T_4524 & _GEN_617; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [491:0] _T_4930 = {_T_4921,_T_4557,_T_4553,_T_4549,_T_4545,_T_4541,_T_4537,_T_4533,_T_4529,_T_4525}; // @[Cat.scala 29:58]
  wire  _T_4518 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4520 = _T_4518 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4091; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_4091[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4521 = _T_4520 & _GEN_618; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4514 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4516 = _T_4514 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4088; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_4088[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4517 = _T_4516 & _GEN_619; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4510 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4512 = _T_4510 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4085; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_4085[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4513 = _T_4512 & _GEN_620; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4506 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4508 = _T_4506 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4082; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_4082[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4509 = _T_4508 & _GEN_621; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4502 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4504 = _T_4502 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4079; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_4079[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4505 = _T_4504 & _GEN_622; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4498 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4500 = _T_4498 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4076; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_4076[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4501 = _T_4500 & _GEN_623; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4494 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4496 = _T_4494 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4073; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_4073[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4497 = _T_4496 & _GEN_624; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4490 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4492 = _T_4490 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4070; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_4070[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4493 = _T_4492 & _GEN_625; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4486 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4488 = _T_4486 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4067; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_4067[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4489 = _T_4488 & _GEN_626; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [545:0] _T_4939 = {_T_4930,_T_4521,_T_4517,_T_4513,_T_4509,_T_4505,_T_4501,_T_4497,_T_4493,_T_4489}; // @[Cat.scala 29:58]
  wire  _T_4482 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4484 = _T_4482 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4064; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_4064[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4485 = _T_4484 & _GEN_627; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4478 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4480 = _T_4478 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4061; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_4061[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4481 = _T_4480 & _GEN_628; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4474 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4476 = _T_4474 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4058; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_4058[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4477 = _T_4476 & _GEN_629; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4470 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4472 = _T_4470 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4055; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_4055[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4473 = _T_4472 & _GEN_630; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4466 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4468 = _T_4466 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4052; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_4052[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4469 = _T_4468 & _GEN_631; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4462 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4464 = _T_4462 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4049; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_4049[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4465 = _T_4464 & _GEN_632; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4458 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4460 = _T_4458 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4046; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_4046[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4461 = _T_4460 & _GEN_633; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4454 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4456 = _T_4454 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4043; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_4043[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4457 = _T_4456 & _GEN_634; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4450 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4452 = _T_4450 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4040; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_4040[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4453 = _T_4452 & _GEN_635; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [599:0] _T_4948 = {_T_4939,_T_4485,_T_4481,_T_4477,_T_4473,_T_4469,_T_4465,_T_4461,_T_4457,_T_4453}; // @[Cat.scala 29:58]
  wire  _T_4446 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4448 = _T_4446 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4037; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_4037[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4449 = _T_4448 & _GEN_636; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4442 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4444 = _T_4442 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4034; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_4034[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4445 = _T_4444 & _GEN_637; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4438 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4440 = _T_4438 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4031; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_4031[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4441 = _T_4440 & _GEN_638; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4434 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4436 = _T_4434 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4028; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_4028[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4437 = _T_4436 & _GEN_639; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4430 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4432 = _T_4430 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4025; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_4025[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4433 = _T_4432 & _GEN_640; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4426 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4428 = _T_4426 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4022; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_4022[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4429 = _T_4428 & _GEN_641; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4422 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4424 = _T_4422 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4019; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_4019[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4425 = _T_4424 & _GEN_642; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4418 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4420 = _T_4418 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4016; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_4016[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4421 = _T_4420 & _GEN_643; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4414 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4416 = _T_4414 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4013; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_4013[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4417 = _T_4416 & _GEN_644; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [653:0] _T_4957 = {_T_4948,_T_4449,_T_4445,_T_4441,_T_4437,_T_4433,_T_4429,_T_4425,_T_4421,_T_4417}; // @[Cat.scala 29:58]
  wire  _T_4410 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4412 = _T_4410 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4010; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_4010[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4413 = _T_4412 & _GEN_645; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4406 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4408 = _T_4406 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4007; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_4007[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4409 = _T_4408 & _GEN_646; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4402 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4404 = _T_4402 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4004; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_4004[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4405 = _T_4404 & _GEN_647; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4398 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4400 = _T_4398 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4001; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_4001[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4401 = _T_4400 & _GEN_648; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4394 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4396 = _T_4394 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3998; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_3998[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4397 = _T_4396 & _GEN_649; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4390 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4392 = _T_4390 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3995; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_3995[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4393 = _T_4392 & _GEN_650; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4386 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4388 = _T_4386 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3992; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_3992[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4389 = _T_4388 & _GEN_651; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4382 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4384 = _T_4382 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3989; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_3989[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4385 = _T_4384 & _GEN_652; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4378 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4380 = _T_4378 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3986; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_3986[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4381 = _T_4380 & _GEN_653; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [707:0] _T_4966 = {_T_4957,_T_4413,_T_4409,_T_4405,_T_4401,_T_4397,_T_4393,_T_4389,_T_4385,_T_4381}; // @[Cat.scala 29:58]
  wire  _T_4374 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4376 = _T_4374 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3983; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3983[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4377 = _T_4376 & _GEN_654; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4370 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4372 = _T_4370 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3980; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3980[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4373 = _T_4372 & _GEN_655; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4366 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4368 = _T_4366 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3977; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3977[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4369 = _T_4368 & _GEN_656; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4362 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4364 = _T_4362 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3974; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3974[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4365 = _T_4364 & _GEN_657; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4358 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4360 = _T_4358 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3971; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3971[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4361 = _T_4360 & _GEN_658; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4354 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4356 = _T_4354 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3968; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3968[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4357 = _T_4356 & _GEN_659; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4350 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4352 = _T_4350 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3965; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3965[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4353 = _T_4352 & _GEN_660; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4346 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4348 = _T_4346 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3962; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3962[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4349 = _T_4348 & _GEN_661; // @[el2_ifu_mem_ctl.scala 713:130]
  wire  _T_4342 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4344 = _T_4342 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3959; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3959[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4345 = _T_4344 & _GEN_662; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [761:0] _T_4975 = {_T_4966,_T_4377,_T_4373,_T_4369,_T_4365,_T_4361,_T_4357,_T_4353,_T_4349,_T_4345}; // @[Cat.scala 29:58]
  wire  _T_4338 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 713:121]
  wire [5:0] _T_4340 = _T_4338 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3956; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3956[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [5:0] _T_4341 = _T_4340 & _GEN_663; // @[el2_ifu_mem_ctl.scala 713:130]
  wire [767:0] _T_4976 = {_T_4975,_T_4341}; // @[Cat.scala 29:58]
  wire  way_status = _T_4976[0]; // @[el2_ifu_mem_ctl.scala 713:16]
  wire  _T_187 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 253:96]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 257:25]
  wire [2:0] _T_198 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_198; // @[el2_ifu_mem_ctl.scala 262:45]
  wire  _T_204 = _T_223 | _T_231; // @[el2_ifu_mem_ctl.scala 267:59]
  wire  _T_206 = _T_204 | _T_2219; // @[el2_ifu_mem_ctl.scala 267:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_206; // @[el2_ifu_mem_ctl.scala 267:41]
  wire  _T_211 = _T_219 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 273:39]
  wire  _T_213 = _T_211 & _T_187; // @[el2_ifu_mem_ctl.scala 273:60]
  wire  _T_217 = _T_213 & _T_204; // @[el2_ifu_mem_ctl.scala 273:78]
  wire  ic_act_hit_f = _T_217 & _T_239; // @[el2_ifu_mem_ctl.scala 273:126]
  wire  _T_254 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 280:31]
  wire  _T_255 = _T_254 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 280:46]
  wire  _T_256 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 280:94]
  wire  uncacheable_miss_in = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 281:84]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2605 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 609:48]
  wire  _T_2606 = _T_2605 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 609:52]
  wire  bus_ifu_wr_data_error_ff = _T_2606 & miss_pending; // @[el2_ifu_mem_ctl.scala 609:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 356:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 355:55]
  wire  _T_268 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 284:145]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 536:52]
  wire  _T_289 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 296:36]
  wire  _T_290 = miss_pending & _T_289; // @[el2_ifu_mem_ctl.scala 296:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 297:25]
  wire  _T_291 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 296:72]
  wire  reset_ic_in = _T_290 & _T_291; // @[el2_ifu_mem_ctl.scala 296:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 298:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 306:23]
  wire  _T_305 = _T_2233 & flush_final_f; // @[el2_ifu_mem_ctl.scala 310:87]
  wire  _T_306 = ~_T_305; // @[el2_ifu_mem_ctl.scala 310:55]
  wire  _T_307 = io_ifc_fetch_req_bf & _T_306; // @[el2_ifu_mem_ctl.scala 310:53]
  wire  stream_miss_f = stream_hit_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 447:83]
  wire  _T_308 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 310:106]
  wire  ifc_fetch_req_qual_bf = _T_307 & _T_308; // @[el2_ifu_mem_ctl.scala 310:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 316:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_315 = _T_231 | _T_2219; // @[el2_ifu_mem_ctl.scala 318:55]
  wire  _T_318 = _T_315 & _T_59; // @[el2_ifu_mem_ctl.scala 318:82]
  wire  _T_2239 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 452:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2239}; // @[Cat.scala 29:58]
  wire  _T_2240 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2264 = _T_2240 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2243 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2265 = _T_2243 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2272 = _T_2264 | _T_2265; // @[Mux.scala 27:72]
  wire  _T_2246 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2266 = _T_2246 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2273 = _T_2272 | _T_2266; // @[Mux.scala 27:72]
  wire  _T_2249 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2267 = _T_2249 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2274 = _T_2273 | _T_2267; // @[Mux.scala 27:72]
  wire  _T_2252 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2268 = _T_2252 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2275 = _T_2274 | _T_2268; // @[Mux.scala 27:72]
  wire  _T_2255 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2269 = _T_2255 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2276 = _T_2275 | _T_2269; // @[Mux.scala 27:72]
  wire  _T_2258 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2270 = _T_2258 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2277 = _T_2276 | _T_2270; // @[Mux.scala 27:72]
  wire  _T_2261 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2271 = _T_2261 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2277 | _T_2271; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 454:46]
  wire  _T_322 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 322:35]
  wire  _T_324 = _T_322 & _T_52; // @[el2_ifu_mem_ctl.scala 322:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 606:61]
  wire  _T_2599 = ic_act_miss_f_delayed & _T_2234; // @[el2_ifu_mem_ctl.scala 607:53]
  wire  reset_tag_valid_for_miss = _T_2599 & _T_52; // @[el2_ifu_mem_ctl.scala 607:84]
  wire  sel_mb_addr = _T_324 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 322:79]
  wire [30:0] _T_329 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_331 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 324:37]
  wire [30:0] _T_332 = sel_mb_addr ? _T_329 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_333 = _T_331 ? ifu_fetch_addr_int_f : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_332 | _T_333; // @[Mux.scala 27:72]
  wire  _T_338 = _T_324 & last_beat; // @[el2_ifu_mem_ctl.scala 326:84]
  wire  _T_2593 = ~_T_2605; // @[el2_ifu_mem_ctl.scala 604:84]
  wire  _T_2594 = _T_92 & _T_2593; // @[el2_ifu_mem_ctl.scala 604:82]
  wire  bus_ifu_wr_en_ff_q = _T_2594 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 604:108]
  wire  sel_mb_status_addr = _T_338 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 326:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_329 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 327:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [7:0] _T_562 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_571 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_562}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_579 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_588 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_579}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_589 = {_T_588,_T_571}; // @[el2_lib.scala 348:27]
  wire  _T_590 = ^_T_589; // @[el2_lib.scala 348:34]
  wire [7:0] _T_597 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_606 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_597}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_614 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_623 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_614}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_624 = {_T_623,_T_606}; // @[el2_lib.scala 348:44]
  wire  _T_625 = ^_T_624; // @[el2_lib.scala 348:51]
  wire [7:0] _T_632 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_641 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_632}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_649 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_658 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_649}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_659 = {_T_658,_T_641}; // @[el2_lib.scala 348:61]
  wire  _T_660 = ^_T_659; // @[el2_lib.scala 348:68]
  wire [6:0] _T_666 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_674 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_666}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_681 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_690 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_681,_T_674}; // @[el2_lib.scala 348:78]
  wire  _T_691 = ^_T_690; // @[el2_lib.scala 348:85]
  wire [6:0] _T_697 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_705 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_697}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_712 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_721 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_712,_T_705}; // @[el2_lib.scala 348:95]
  wire  _T_722 = ^_T_721; // @[el2_lib.scala 348:102]
  wire [6:0] _T_728 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_736 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_728}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_752 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_712,_T_736}; // @[el2_lib.scala 348:112]
  wire  _T_753 = ^_T_752; // @[el2_lib.scala 348:119]
  wire [6:0] _T_759 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 348:129]
  wire  _T_760 = ^_T_759; // @[el2_lib.scala 348:136]
  wire [3:0] _T_2280 = {ifu_bus_rid_ff[2:1],_T_2239,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2281 = _T_2280 == 4'h0; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1287; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_0 = _T_1287[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2328 = _T_2281 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2284 = _T_2280 == 4'h1; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1289; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_1 = _T_1289[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2329 = _T_2284 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2344 = _T_2328 | _T_2329; // @[Mux.scala 27:72]
  wire  _T_2287 = _T_2280 == 4'h2; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1291; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_2 = _T_1291[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2330 = _T_2287 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2345 = _T_2344 | _T_2330; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2280 == 4'h3; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1293; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_3 = _T_1293[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2331 = _T_2290 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2346 = _T_2345 | _T_2331; // @[Mux.scala 27:72]
  wire  _T_2293 = _T_2280 == 4'h4; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1295; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_4 = _T_1295[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2332 = _T_2293 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2347 = _T_2346 | _T_2332; // @[Mux.scala 27:72]
  wire  _T_2296 = _T_2280 == 4'h5; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1297; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_5 = _T_1297[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2333 = _T_2296 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2348 = _T_2347 | _T_2333; // @[Mux.scala 27:72]
  wire  _T_2299 = _T_2280 == 4'h6; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1299; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_6 = _T_1299[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2334 = _T_2299 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2349 = _T_2348 | _T_2334; // @[Mux.scala 27:72]
  wire  _T_2302 = _T_2280 == 4'h7; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1301; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_7 = _T_1301[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2335 = _T_2302 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2350 = _T_2349 | _T_2335; // @[Mux.scala 27:72]
  wire  _T_2305 = _T_2280 == 4'h8; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1303; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_8 = _T_1303[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2336 = _T_2305 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2351 = _T_2350 | _T_2336; // @[Mux.scala 27:72]
  wire  _T_2308 = _T_2280 == 4'h9; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1305; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_9 = _T_1305[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2337 = _T_2308 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2352 = _T_2351 | _T_2337; // @[Mux.scala 27:72]
  wire  _T_2311 = _T_2280 == 4'ha; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1307; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_10 = _T_1307[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2338 = _T_2311 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2353 = _T_2352 | _T_2338; // @[Mux.scala 27:72]
  wire  _T_2314 = _T_2280 == 4'hb; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1309; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_11 = _T_1309[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2339 = _T_2314 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2354 = _T_2353 | _T_2339; // @[Mux.scala 27:72]
  wire  _T_2317 = _T_2280 == 4'hc; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1311; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_12 = _T_1311[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2340 = _T_2317 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2355 = _T_2354 | _T_2340; // @[Mux.scala 27:72]
  wire  _T_2320 = _T_2280 == 4'hd; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1313; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_13 = _T_1313[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2341 = _T_2320 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2356 = _T_2355 | _T_2341; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2280 == 4'he; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1315; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_14 = _T_1315[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2342 = _T_2323 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2357 = _T_2356 | _T_2342; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2280 == 4'hf; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1317; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_15 = _T_1317[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2343 = _T_2326 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2358 = _T_2357 | _T_2343; // @[Mux.scala 27:72]
  wire [3:0] _T_2360 = {ifu_bus_rid_ff[2:1],_T_2239,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2361 = _T_2360 == 4'h0; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2384 = _T_2361 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2364 = _T_2360 == 4'h1; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2385 = _T_2364 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2392 = _T_2384 | _T_2385; // @[Mux.scala 27:72]
  wire  _T_2367 = _T_2360 == 4'h2; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2386 = _T_2367 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2393 = _T_2392 | _T_2386; // @[Mux.scala 27:72]
  wire  _T_2370 = _T_2360 == 4'h3; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2387 = _T_2370 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2394 = _T_2393 | _T_2387; // @[Mux.scala 27:72]
  wire  _T_2373 = _T_2360 == 4'h4; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2388 = _T_2373 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2395 = _T_2394 | _T_2388; // @[Mux.scala 27:72]
  wire  _T_2376 = _T_2360 == 4'h5; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2389 = _T_2376 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2396 = _T_2395 | _T_2389; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2360 == 4'h6; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2390 = _T_2379 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2397 = _T_2396 | _T_2390; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2360 == 4'h7; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2391 = _T_2382 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2398 = _T_2397 | _T_2391; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2358,_T_2398}; // @[Cat.scala 29:58]
  wire [7:0] _T_984 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_993 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_984}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_1001 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_1010 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1001}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_1011 = {_T_1010,_T_993}; // @[el2_lib.scala 348:27]
  wire  _T_1012 = ^_T_1011; // @[el2_lib.scala 348:34]
  wire [7:0] _T_1019 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_1028 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1019}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_1036 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_1045 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1036}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_1046 = {_T_1045,_T_1028}; // @[el2_lib.scala 348:44]
  wire  _T_1047 = ^_T_1046; // @[el2_lib.scala 348:51]
  wire [7:0] _T_1054 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_1063 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1054}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_1071 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_1080 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1071}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_1081 = {_T_1080,_T_1063}; // @[el2_lib.scala 348:61]
  wire  _T_1082 = ^_T_1081; // @[el2_lib.scala 348:68]
  wire [6:0] _T_1088 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_1096 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1088}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_1103 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_1112 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1103,_T_1096}; // @[el2_lib.scala 348:78]
  wire  _T_1113 = ^_T_1112; // @[el2_lib.scala 348:85]
  wire [6:0] _T_1119 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_1127 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1119}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_1134 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_1143 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1134,_T_1127}; // @[el2_lib.scala 348:95]
  wire  _T_1144 = ^_T_1143; // @[el2_lib.scala 348:102]
  wire [6:0] _T_1150 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_1158 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_1150}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_1174 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1134,_T_1158}; // @[el2_lib.scala 348:112]
  wire  _T_1175 = ^_T_1174; // @[el2_lib.scala 348:119]
  wire [6:0] _T_1181 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 348:129]
  wire  _T_1182 = ^_T_1181; // @[el2_lib.scala 348:136]
  wire [70:0] _T_1229 = {_T_590,_T_625,_T_660,_T_691,_T_722,_T_753,_T_760,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1228 = {_T_1012,_T_1047,_T_1082,_T_1113,_T_1144,_T_1175,_T_1182,_T_2358,_T_2398}; // @[Cat.scala 29:58]
  wire [141:0] _T_1230 = {_T_590,_T_625,_T_660,_T_691,_T_722,_T_753,_T_760,ifu_bus_rdata_ff,_T_1228}; // @[Cat.scala 29:58]
  wire [141:0] _T_1233 = {_T_1012,_T_1047,_T_1082,_T_1113,_T_1144,_T_1175,_T_1182,_T_2358,_T_2398,_T_1229}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1230 : _T_1233; // @[el2_ifu_mem_ctl.scala 348:28]
  wire  _T_1190 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 338:56]
  wire  _T_1191 = _T_1190 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 338:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 402:28]
  wire  _T_1393 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  bus_ifu_wr_en = _T_14 & miss_pending; // @[el2_ifu_mem_ctl.scala 602:35]
  wire  _T_1278 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1278; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1319 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 393:118]
  wire  _T_1320 = ic_miss_buff_data_valid[0] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1320; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1416 = _T_1393 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1396 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1279 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1279; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1323 = ic_miss_buff_data_valid[1] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1323; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1417 = _T_1396 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1424 = _T_1416 | _T_1417; // @[Mux.scala 27:72]
  wire  _T_1399 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1280 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1280; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1326 = ic_miss_buff_data_valid[2] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1326; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1418 = _T_1399 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1425 = _T_1424 | _T_1418; // @[Mux.scala 27:72]
  wire  _T_1402 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1281 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1281; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1329 = ic_miss_buff_data_valid[3] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1329; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1419 = _T_1402 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1426 = _T_1425 | _T_1419; // @[Mux.scala 27:72]
  wire  _T_1405 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1282 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1332 = ic_miss_buff_data_valid[4] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1332; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1420 = _T_1405 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1427 = _T_1426 | _T_1420; // @[Mux.scala 27:72]
  wire  _T_1408 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1335 = ic_miss_buff_data_valid[5] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1335; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1421 = _T_1408 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1428 = _T_1427 | _T_1421; // @[Mux.scala 27:72]
  wire  _T_1411 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1284 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1338 = ic_miss_buff_data_valid[6] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1338; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1422 = _T_1411 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1429 = _T_1428 | _T_1422; // @[Mux.scala 27:72]
  wire  _T_1414 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1341 = ic_miss_buff_data_valid[7] & _T_1319; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1341; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1423 = _T_1414 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1429 | _T_1423; // @[Mux.scala 27:72]
  wire  _T_1432 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 405:58]
  wire  _T_1433 = bypass_valid_value_check & _T_1432; // @[el2_ifu_mem_ctl.scala 405:56]
  wire  _T_1435 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 405:77]
  wire  _T_1436 = _T_1433 & _T_1435; // @[el2_ifu_mem_ctl.scala 405:75]
  wire  _T_1441 = _T_1433 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 406:75]
  wire  _T_1442 = _T_1436 | _T_1441; // @[el2_ifu_mem_ctl.scala 405:95]
  wire  _T_1444 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 407:56]
  wire  _T_1447 = _T_1444 & _T_1435; // @[el2_ifu_mem_ctl.scala 407:74]
  wire  _T_1448 = _T_1442 | _T_1447; // @[el2_ifu_mem_ctl.scala 406:94]
  wire  _T_1452 = _T_1444 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 408:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 403:70]
  wire  _T_1453 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1469 = _T_1453 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1455 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1470 = _T_1455 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1477 = _T_1469 | _T_1470; // @[Mux.scala 27:72]
  wire  _T_1457 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1471 = _T_1457 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1478 = _T_1477 | _T_1471; // @[Mux.scala 27:72]
  wire  _T_1459 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1472 = _T_1459 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1479 = _T_1478 | _T_1472; // @[Mux.scala 27:72]
  wire  _T_1461 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1473 = _T_1461 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1480 = _T_1479 | _T_1473; // @[Mux.scala 27:72]
  wire  _T_1463 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1474 = _T_1463 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1481 = _T_1480 | _T_1474; // @[Mux.scala 27:72]
  wire  _T_1465 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1475 = _T_1465 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1482 = _T_1481 | _T_1475; // @[Mux.scala 27:72]
  wire  _T_1467 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1476 = _T_1467 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1483 = _T_1482 | _T_1476; // @[Mux.scala 27:72]
  wire  _T_1485 = _T_1452 & _T_1483; // @[el2_ifu_mem_ctl.scala 408:69]
  wire  _T_1486 = _T_1448 | _T_1485; // @[el2_ifu_mem_ctl.scala 407:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 409:95]
  wire  _T_1489 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 409:95]
  wire  _T_1490 = bypass_valid_value_check & _T_1489; // @[el2_ifu_mem_ctl.scala 409:56]
  wire  bypass_data_ready_in = _T_1486 | _T_1490; // @[el2_ifu_mem_ctl.scala 408:181]
  wire  _T_1491 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 413:53]
  wire  _T_1492 = _T_1491 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 413:73]
  wire  _T_1494 = _T_1492 & _T_309; // @[el2_ifu_mem_ctl.scala 413:96]
  wire  _T_1496 = _T_1494 & _T_61; // @[el2_ifu_mem_ctl.scala 413:118]
  wire  _T_1498 = crit_wd_byp_ok_ff & _T_52; // @[el2_ifu_mem_ctl.scala 414:73]
  wire  _T_1500 = _T_1498 & _T_309; // @[el2_ifu_mem_ctl.scala 414:96]
  wire  _T_1502 = _T_1500 & _T_61; // @[el2_ifu_mem_ctl.scala 414:118]
  wire  _T_1503 = _T_1496 | _T_1502; // @[el2_ifu_mem_ctl.scala 413:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 416:58]
  wire  _T_1504 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 415:54]
  wire  _T_1505 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 415:76]
  wire  _T_1506 = _T_1504 & _T_1505; // @[el2_ifu_mem_ctl.scala 415:74]
  wire  _T_1508 = _T_1506 & _T_309; // @[el2_ifu_mem_ctl.scala 415:96]
  wire  ic_crit_wd_rdy_new_in = _T_1503 | _T_1508; // @[el2_ifu_mem_ctl.scala 414:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 612:43]
  wire  _T_1245 = ic_crit_wd_rdy | _T_2219; // @[el2_ifu_mem_ctl.scala 360:38]
  wire  _T_1247 = _T_1245 | _T_2234; // @[el2_ifu_mem_ctl.scala 360:64]
  wire  _T_1248 = ~_T_1247; // @[el2_ifu_mem_ctl.scala 360:21]
  wire  _T_1249 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 360:98]
  wire  sel_ic_data = _T_1248 & _T_1249; // @[el2_ifu_mem_ctl.scala 360:96]
  wire  _T_2401 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 458:44]
  wire  _T_1602 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 427:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 399:60]
  wire  _T_1546 = _T_1393 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1547 = _T_1396 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1554 = _T_1546 | _T_1547; // @[Mux.scala 27:72]
  wire  _T_1548 = _T_1399 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1554 | _T_1548; // @[Mux.scala 27:72]
  wire  _T_1549 = _T_1402 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1555 | _T_1549; // @[Mux.scala 27:72]
  wire  _T_1550 = _T_1405 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1556 | _T_1550; // @[Mux.scala 27:72]
  wire  _T_1551 = _T_1408 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1558 = _T_1557 | _T_1551; // @[Mux.scala 27:72]
  wire  _T_1552 = _T_1411 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1559 = _T_1558 | _T_1552; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1414 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1559 | _T_1553; // @[Mux.scala 27:72]
  wire  _T_1585 = _T_2146 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1586 = _T_2149 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1593 = _T_1585 | _T_1586; // @[Mux.scala 27:72]
  wire  _T_1587 = _T_2152 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1594 = _T_1593 | _T_1587; // @[Mux.scala 27:72]
  wire  _T_1588 = _T_2155 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1595 = _T_1594 | _T_1588; // @[Mux.scala 27:72]
  wire  _T_1589 = _T_2158 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1596 = _T_1595 | _T_1589; // @[Mux.scala 27:72]
  wire  _T_1590 = _T_2161 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1597 = _T_1596 | _T_1590; // @[Mux.scala 27:72]
  wire  _T_1591 = _T_2164 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1598 = _T_1597 | _T_1591; // @[Mux.scala 27:72]
  wire  _T_1592 = _T_2167 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1598 | _T_1592; // @[Mux.scala 27:72]
  wire  _T_1603 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 429:70]
  wire  ifu_byp_data_err_new = _T_1602 ? ic_miss_buff_data_error_bypass : _T_1603; // @[el2_ifu_mem_ctl.scala 427:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 371:42]
  wire  _T_2402 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 458:91]
  wire  _T_2403 = ~_T_2402; // @[el2_ifu_mem_ctl.scala 458:60]
  wire  ic_rd_parity_final_err = _T_2401 & _T_2403; // @[el2_ifu_mem_ctl.scala 458:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9040 = _T_4338 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 743:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9042 = _T_4342 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9295 = _T_9040 | _T_9042; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9044 = _T_4346 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9296 = _T_9295 | _T_9044; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9046 = _T_4350 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9297 = _T_9296 | _T_9046; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9048 = _T_4354 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9298 = _T_9297 | _T_9048; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9050 = _T_4358 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9299 = _T_9298 | _T_9050; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9052 = _T_4362 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9300 = _T_9299 | _T_9052; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9054 = _T_4366 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9301 = _T_9300 | _T_9054; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9056 = _T_4370 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9302 = _T_9301 | _T_9056; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9058 = _T_4374 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9303 = _T_9302 | _T_9058; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9060 = _T_4378 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9304 = _T_9303 | _T_9060; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9062 = _T_4382 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9305 = _T_9304 | _T_9062; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9064 = _T_4386 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9306 = _T_9305 | _T_9064; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9066 = _T_4390 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9307 = _T_9306 | _T_9066; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9068 = _T_4394 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9308 = _T_9307 | _T_9068; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9070 = _T_4398 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9309 = _T_9308 | _T_9070; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9072 = _T_4402 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9310 = _T_9309 | _T_9072; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9074 = _T_4406 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9311 = _T_9310 | _T_9074; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9076 = _T_4410 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9312 = _T_9311 | _T_9076; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9078 = _T_4414 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9313 = _T_9312 | _T_9078; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9080 = _T_4418 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9314 = _T_9313 | _T_9080; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9082 = _T_4422 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9315 = _T_9314 | _T_9082; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9084 = _T_4426 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9316 = _T_9315 | _T_9084; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9086 = _T_4430 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9317 = _T_9316 | _T_9086; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9088 = _T_4434 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9318 = _T_9317 | _T_9088; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9090 = _T_4438 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9319 = _T_9318 | _T_9090; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9092 = _T_4442 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9320 = _T_9319 | _T_9092; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9094 = _T_4446 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9321 = _T_9320 | _T_9094; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9096 = _T_4450 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9322 = _T_9321 | _T_9096; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9098 = _T_4454 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9323 = _T_9322 | _T_9098; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9100 = _T_4458 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9324 = _T_9323 | _T_9100; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9102 = _T_4462 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9325 = _T_9324 | _T_9102; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9104 = _T_4466 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9326 = _T_9325 | _T_9104; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9106 = _T_4470 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9327 = _T_9326 | _T_9106; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9108 = _T_4474 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9328 = _T_9327 | _T_9108; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9110 = _T_4478 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9329 = _T_9328 | _T_9110; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9112 = _T_4482 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9330 = _T_9329 | _T_9112; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9114 = _T_4486 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9331 = _T_9330 | _T_9114; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9116 = _T_4490 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9332 = _T_9331 | _T_9116; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9118 = _T_4494 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9333 = _T_9332 | _T_9118; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9120 = _T_4498 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9334 = _T_9333 | _T_9120; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9122 = _T_4502 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9335 = _T_9334 | _T_9122; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9124 = _T_4506 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9336 = _T_9335 | _T_9124; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9126 = _T_4510 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9337 = _T_9336 | _T_9126; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9128 = _T_4514 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9338 = _T_9337 | _T_9128; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9130 = _T_4518 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9339 = _T_9338 | _T_9130; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9132 = _T_4522 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9340 = _T_9339 | _T_9132; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9134 = _T_4526 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9341 = _T_9340 | _T_9134; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9136 = _T_4530 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9342 = _T_9341 | _T_9136; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9138 = _T_4534 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9343 = _T_9342 | _T_9138; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9140 = _T_4538 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9344 = _T_9343 | _T_9140; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9142 = _T_4542 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9345 = _T_9344 | _T_9142; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9144 = _T_4546 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9346 = _T_9345 | _T_9144; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9146 = _T_4550 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9347 = _T_9346 | _T_9146; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9148 = _T_4554 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9348 = _T_9347 | _T_9148; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9150 = _T_4558 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9349 = _T_9348 | _T_9150; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9152 = _T_4562 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9350 = _T_9349 | _T_9152; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9154 = _T_4566 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9351 = _T_9350 | _T_9154; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9156 = _T_4570 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9352 = _T_9351 | _T_9156; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9158 = _T_4574 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9353 = _T_9352 | _T_9158; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9160 = _T_4578 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9354 = _T_9353 | _T_9160; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9162 = _T_4582 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9355 = _T_9354 | _T_9162; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9164 = _T_4586 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9356 = _T_9355 | _T_9164; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9166 = _T_4590 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9357 = _T_9356 | _T_9166; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9168 = _T_4594 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9358 = _T_9357 | _T_9168; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9170 = _T_4598 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9359 = _T_9358 | _T_9170; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9172 = _T_4602 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9360 = _T_9359 | _T_9172; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9174 = _T_4606 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9361 = _T_9360 | _T_9174; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9176 = _T_4610 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9362 = _T_9361 | _T_9176; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9178 = _T_4614 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9363 = _T_9362 | _T_9178; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9180 = _T_4618 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9364 = _T_9363 | _T_9180; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9182 = _T_4622 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9365 = _T_9364 | _T_9182; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9184 = _T_4626 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9366 = _T_9365 | _T_9184; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9186 = _T_4630 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9367 = _T_9366 | _T_9186; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9188 = _T_4634 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9368 = _T_9367 | _T_9188; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9190 = _T_4638 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9369 = _T_9368 | _T_9190; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9192 = _T_4642 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9370 = _T_9369 | _T_9192; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9194 = _T_4646 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9371 = _T_9370 | _T_9194; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9196 = _T_4650 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9372 = _T_9371 | _T_9196; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9198 = _T_4654 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9373 = _T_9372 | _T_9198; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9200 = _T_4658 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9374 = _T_9373 | _T_9200; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9202 = _T_4662 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9375 = _T_9374 | _T_9202; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9204 = _T_4666 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9376 = _T_9375 | _T_9204; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9206 = _T_4670 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9377 = _T_9376 | _T_9206; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9208 = _T_4674 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9378 = _T_9377 | _T_9208; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9210 = _T_4678 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9379 = _T_9378 | _T_9210; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9212 = _T_4682 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9380 = _T_9379 | _T_9212; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9214 = _T_4686 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9381 = _T_9380 | _T_9214; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9216 = _T_4690 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9382 = _T_9381 | _T_9216; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9218 = _T_4694 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9383 = _T_9382 | _T_9218; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9220 = _T_4698 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9384 = _T_9383 | _T_9220; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9222 = _T_4702 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9385 = _T_9384 | _T_9222; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9224 = _T_4706 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9386 = _T_9385 | _T_9224; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9226 = _T_4710 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9387 = _T_9386 | _T_9226; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9228 = _T_4714 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9388 = _T_9387 | _T_9228; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9230 = _T_4718 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9389 = _T_9388 | _T_9230; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9232 = _T_4722 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9390 = _T_9389 | _T_9232; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9234 = _T_4726 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9391 = _T_9390 | _T_9234; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9236 = _T_4730 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9392 = _T_9391 | _T_9236; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9238 = _T_4734 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9393 = _T_9392 | _T_9238; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9240 = _T_4738 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9394 = _T_9393 | _T_9240; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9242 = _T_4742 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9395 = _T_9394 | _T_9242; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9244 = _T_4746 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9396 = _T_9395 | _T_9244; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9246 = _T_4750 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9397 = _T_9396 | _T_9246; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9248 = _T_4754 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9398 = _T_9397 | _T_9248; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9250 = _T_4758 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9399 = _T_9398 | _T_9250; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9252 = _T_4762 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9400 = _T_9399 | _T_9252; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9254 = _T_4766 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9401 = _T_9400 | _T_9254; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9256 = _T_4770 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9402 = _T_9401 | _T_9256; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9258 = _T_4774 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9403 = _T_9402 | _T_9258; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9260 = _T_4778 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9404 = _T_9403 | _T_9260; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9262 = _T_4782 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9405 = _T_9404 | _T_9262; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9264 = _T_4786 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9406 = _T_9405 | _T_9264; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9266 = _T_4790 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9407 = _T_9406 | _T_9266; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9268 = _T_4794 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9408 = _T_9407 | _T_9268; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9270 = _T_4798 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9409 = _T_9408 | _T_9270; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9272 = _T_4802 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9410 = _T_9409 | _T_9272; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9274 = _T_4806 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9411 = _T_9410 | _T_9274; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9276 = _T_4810 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9412 = _T_9411 | _T_9276; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9278 = _T_4814 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9413 = _T_9412 | _T_9278; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9280 = _T_4818 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9414 = _T_9413 | _T_9280; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9282 = _T_4822 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9415 = _T_9414 | _T_9282; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9284 = _T_4826 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9416 = _T_9415 | _T_9284; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9286 = _T_4830 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9417 = _T_9416 | _T_9286; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9288 = _T_4834 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9418 = _T_9417 | _T_9288; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9290 = _T_4838 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9419 = _T_9418 | _T_9290; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9292 = _T_4842 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9420 = _T_9419 | _T_9292; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9294 = _T_4846 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9421 = _T_9420 | _T_9294; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8657 = _T_4338 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 743:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8659 = _T_4342 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8912 = _T_8657 | _T_8659; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8661 = _T_4346 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8913 = _T_8912 | _T_8661; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8663 = _T_4350 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8914 = _T_8913 | _T_8663; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8665 = _T_4354 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8915 = _T_8914 | _T_8665; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8667 = _T_4358 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8916 = _T_8915 | _T_8667; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8669 = _T_4362 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8917 = _T_8916 | _T_8669; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8671 = _T_4366 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8918 = _T_8917 | _T_8671; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8673 = _T_4370 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8919 = _T_8918 | _T_8673; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8675 = _T_4374 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8920 = _T_8919 | _T_8675; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8677 = _T_4378 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8921 = _T_8920 | _T_8677; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8679 = _T_4382 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8922 = _T_8921 | _T_8679; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8681 = _T_4386 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8923 = _T_8922 | _T_8681; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8683 = _T_4390 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8924 = _T_8923 | _T_8683; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8685 = _T_4394 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8925 = _T_8924 | _T_8685; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8687 = _T_4398 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8926 = _T_8925 | _T_8687; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8689 = _T_4402 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8927 = _T_8926 | _T_8689; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8691 = _T_4406 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8928 = _T_8927 | _T_8691; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8693 = _T_4410 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8929 = _T_8928 | _T_8693; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8695 = _T_4414 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8930 = _T_8929 | _T_8695; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8697 = _T_4418 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8931 = _T_8930 | _T_8697; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8699 = _T_4422 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8932 = _T_8931 | _T_8699; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8701 = _T_4426 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8933 = _T_8932 | _T_8701; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8703 = _T_4430 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8934 = _T_8933 | _T_8703; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8705 = _T_4434 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8935 = _T_8934 | _T_8705; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8707 = _T_4438 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8936 = _T_8935 | _T_8707; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8709 = _T_4442 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8937 = _T_8936 | _T_8709; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8711 = _T_4446 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8938 = _T_8937 | _T_8711; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8713 = _T_4450 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8939 = _T_8938 | _T_8713; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8715 = _T_4454 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8940 = _T_8939 | _T_8715; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_8717 = _T_4458 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8941 = _T_8940 | _T_8717; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_8719 = _T_4462 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8942 = _T_8941 | _T_8719; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_8721 = _T_4466 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8943 = _T_8942 | _T_8721; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_8723 = _T_4470 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8944 = _T_8943 | _T_8723; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_8725 = _T_4474 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8945 = _T_8944 | _T_8725; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_8727 = _T_4478 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8946 = _T_8945 | _T_8727; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_8729 = _T_4482 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8947 = _T_8946 | _T_8729; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_8731 = _T_4486 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8948 = _T_8947 | _T_8731; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_8733 = _T_4490 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8949 = _T_8948 | _T_8733; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_8735 = _T_4494 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8950 = _T_8949 | _T_8735; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_8737 = _T_4498 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8951 = _T_8950 | _T_8737; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_8739 = _T_4502 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8952 = _T_8951 | _T_8739; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_8741 = _T_4506 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8953 = _T_8952 | _T_8741; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_8743 = _T_4510 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8954 = _T_8953 | _T_8743; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_8745 = _T_4514 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8955 = _T_8954 | _T_8745; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_8747 = _T_4518 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8956 = _T_8955 | _T_8747; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_8749 = _T_4522 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8957 = _T_8956 | _T_8749; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_8751 = _T_4526 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8958 = _T_8957 | _T_8751; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_8753 = _T_4530 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8959 = _T_8958 | _T_8753; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_8755 = _T_4534 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8960 = _T_8959 | _T_8755; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_8757 = _T_4538 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8961 = _T_8960 | _T_8757; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_8759 = _T_4542 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8962 = _T_8961 | _T_8759; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_8761 = _T_4546 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8963 = _T_8962 | _T_8761; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_8763 = _T_4550 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8964 = _T_8963 | _T_8763; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_8765 = _T_4554 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8965 = _T_8964 | _T_8765; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_8767 = _T_4558 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8966 = _T_8965 | _T_8767; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_8769 = _T_4562 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8967 = _T_8966 | _T_8769; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_8771 = _T_4566 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8968 = _T_8967 | _T_8771; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_8773 = _T_4570 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8969 = _T_8968 | _T_8773; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_8775 = _T_4574 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8970 = _T_8969 | _T_8775; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_8777 = _T_4578 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8971 = _T_8970 | _T_8777; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_8779 = _T_4582 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8972 = _T_8971 | _T_8779; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_8781 = _T_4586 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8973 = _T_8972 | _T_8781; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_8783 = _T_4590 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8974 = _T_8973 | _T_8783; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_8785 = _T_4594 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8975 = _T_8974 | _T_8785; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_8787 = _T_4598 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8976 = _T_8975 | _T_8787; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_8789 = _T_4602 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8977 = _T_8976 | _T_8789; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_8791 = _T_4606 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8978 = _T_8977 | _T_8791; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_8793 = _T_4610 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8979 = _T_8978 | _T_8793; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_8795 = _T_4614 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8980 = _T_8979 | _T_8795; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_8797 = _T_4618 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8981 = _T_8980 | _T_8797; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_8799 = _T_4622 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8982 = _T_8981 | _T_8799; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_8801 = _T_4626 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8983 = _T_8982 | _T_8801; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_8803 = _T_4630 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8984 = _T_8983 | _T_8803; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_8805 = _T_4634 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8985 = _T_8984 | _T_8805; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_8807 = _T_4638 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8986 = _T_8985 | _T_8807; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_8809 = _T_4642 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8987 = _T_8986 | _T_8809; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_8811 = _T_4646 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8988 = _T_8987 | _T_8811; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_8813 = _T_4650 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8989 = _T_8988 | _T_8813; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_8815 = _T_4654 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8990 = _T_8989 | _T_8815; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_8817 = _T_4658 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8991 = _T_8990 | _T_8817; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_8819 = _T_4662 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8992 = _T_8991 | _T_8819; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_8821 = _T_4666 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8993 = _T_8992 | _T_8821; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_8823 = _T_4670 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8994 = _T_8993 | _T_8823; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_8825 = _T_4674 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8995 = _T_8994 | _T_8825; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_8827 = _T_4678 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8996 = _T_8995 | _T_8827; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_8829 = _T_4682 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8997 = _T_8996 | _T_8829; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_8831 = _T_4686 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8998 = _T_8997 | _T_8831; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_8833 = _T_4690 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_8999 = _T_8998 | _T_8833; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_8835 = _T_4694 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9000 = _T_8999 | _T_8835; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_8837 = _T_4698 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9001 = _T_9000 | _T_8837; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_8839 = _T_4702 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9002 = _T_9001 | _T_8839; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_8841 = _T_4706 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9003 = _T_9002 | _T_8841; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_8843 = _T_4710 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9004 = _T_9003 | _T_8843; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_8845 = _T_4714 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9005 = _T_9004 | _T_8845; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_8847 = _T_4718 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9006 = _T_9005 | _T_8847; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_8849 = _T_4722 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9007 = _T_9006 | _T_8849; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_8851 = _T_4726 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9008 = _T_9007 | _T_8851; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_8853 = _T_4730 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9009 = _T_9008 | _T_8853; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_8855 = _T_4734 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9010 = _T_9009 | _T_8855; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_8857 = _T_4738 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9011 = _T_9010 | _T_8857; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_8859 = _T_4742 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9012 = _T_9011 | _T_8859; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_8861 = _T_4746 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9013 = _T_9012 | _T_8861; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_8863 = _T_4750 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9014 = _T_9013 | _T_8863; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_8865 = _T_4754 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9015 = _T_9014 | _T_8865; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_8867 = _T_4758 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9016 = _T_9015 | _T_8867; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_8869 = _T_4762 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9017 = _T_9016 | _T_8869; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_8871 = _T_4766 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9018 = _T_9017 | _T_8871; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_8873 = _T_4770 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9019 = _T_9018 | _T_8873; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_8875 = _T_4774 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9020 = _T_9019 | _T_8875; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_8877 = _T_4778 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9021 = _T_9020 | _T_8877; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_8879 = _T_4782 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9022 = _T_9021 | _T_8879; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_8881 = _T_4786 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9023 = _T_9022 | _T_8881; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_8883 = _T_4790 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9024 = _T_9023 | _T_8883; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_8885 = _T_4794 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9025 = _T_9024 | _T_8885; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_8887 = _T_4798 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9026 = _T_9025 | _T_8887; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_8889 = _T_4802 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9027 = _T_9026 | _T_8889; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_8891 = _T_4806 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9028 = _T_9027 | _T_8891; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_8893 = _T_4810 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9029 = _T_9028 | _T_8893; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_8895 = _T_4814 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9030 = _T_9029 | _T_8895; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_8897 = _T_4818 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9031 = _T_9030 | _T_8897; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_8899 = _T_4822 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9032 = _T_9031 | _T_8899; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_8901 = _T_4826 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9033 = _T_9032 | _T_8901; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_8903 = _T_4830 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9034 = _T_9033 | _T_8903; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_8905 = _T_4834 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9035 = _T_9034 | _T_8905; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_8907 = _T_4838 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9036 = _T_9035 | _T_8907; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_8909 = _T_4842 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9037 = _T_9036 | _T_8909; // @[el2_ifu_mem_ctl.scala 743:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_8911 = _T_4846 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 743:10]
  wire  _T_9038 = _T_9037 | _T_8911; // @[el2_ifu_mem_ctl.scala 743:91]
  wire [1:0] ic_tag_valid_unq = {_T_9421,_T_9038}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 814:54]
  wire [1:0] _T_9460 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9461 = ic_debug_way_ff & _T_9460; // @[el2_ifu_mem_ctl.scala 797:67]
  wire [1:0] _T_9462 = ic_tag_valid_unq & _T_9461; // @[el2_ifu_mem_ctl.scala 797:48]
  wire  ic_debug_tag_val_rd_out = |_T_9462; // @[el2_ifu_mem_ctl.scala 797:115]
  wire [65:0] _T_1202 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1203; // @[el2_ifu_mem_ctl.scala 344:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2534; // @[el2_ifu_mem_ctl.scala 354:80]
  wire  _T_1243 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 359:98]
  wire  sel_byp_data = _T_1247 & _T_1243; // @[el2_ifu_mem_ctl.scala 359:96]
  wire [63:0] _T_1254 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1255 = _T_1254 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 366:64]
  wire [63:0] _T_1257 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2093 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 435:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1607 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1655 = _T_1607 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1610 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1656 = _T_1610 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1671 = _T_1655 | _T_1656; // @[Mux.scala 27:72]
  wire  _T_1613 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1657 = _T_1613 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1672 = _T_1671 | _T_1657; // @[Mux.scala 27:72]
  wire  _T_1616 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1658 = _T_1616 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1673 = _T_1672 | _T_1658; // @[Mux.scala 27:72]
  wire  _T_1619 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1659 = _T_1619 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1674 = _T_1673 | _T_1659; // @[Mux.scala 27:72]
  wire  _T_1622 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1660 = _T_1622 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1675 = _T_1674 | _T_1660; // @[Mux.scala 27:72]
  wire  _T_1625 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1661 = _T_1625 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1676 = _T_1675 | _T_1661; // @[Mux.scala 27:72]
  wire  _T_1628 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1662 = _T_1628 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1677 = _T_1676 | _T_1662; // @[Mux.scala 27:72]
  wire  _T_1631 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1663 = _T_1631 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1678 = _T_1677 | _T_1663; // @[Mux.scala 27:72]
  wire  _T_1634 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1664 = _T_1634 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1679 = _T_1678 | _T_1664; // @[Mux.scala 27:72]
  wire  _T_1637 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1665 = _T_1637 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1680 = _T_1679 | _T_1665; // @[Mux.scala 27:72]
  wire  _T_1640 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1666 = _T_1640 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1681 = _T_1680 | _T_1666; // @[Mux.scala 27:72]
  wire  _T_1643 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1667 = _T_1643 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1682 = _T_1681 | _T_1667; // @[Mux.scala 27:72]
  wire  _T_1646 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1668 = _T_1646 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1683 = _T_1682 | _T_1668; // @[Mux.scala 27:72]
  wire  _T_1649 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1669 = _T_1649 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1684 = _T_1683 | _T_1669; // @[Mux.scala 27:72]
  wire  _T_1652 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1670 = _T_1652 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1685 = _T_1684 | _T_1670; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1687 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1735 = _T_1687 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1690 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1736 = _T_1690 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1751 = _T_1735 | _T_1736; // @[Mux.scala 27:72]
  wire  _T_1693 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1737 = _T_1693 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1752 = _T_1751 | _T_1737; // @[Mux.scala 27:72]
  wire  _T_1696 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1738 = _T_1696 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1753 = _T_1752 | _T_1738; // @[Mux.scala 27:72]
  wire  _T_1699 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1739 = _T_1699 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1754 = _T_1753 | _T_1739; // @[Mux.scala 27:72]
  wire  _T_1702 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1740 = _T_1702 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1755 = _T_1754 | _T_1740; // @[Mux.scala 27:72]
  wire  _T_1705 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1741 = _T_1705 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1756 = _T_1755 | _T_1741; // @[Mux.scala 27:72]
  wire  _T_1708 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1742 = _T_1708 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1757 = _T_1756 | _T_1742; // @[Mux.scala 27:72]
  wire  _T_1711 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1743 = _T_1711 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1758 = _T_1757 | _T_1743; // @[Mux.scala 27:72]
  wire  _T_1714 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1744 = _T_1714 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1759 = _T_1758 | _T_1744; // @[Mux.scala 27:72]
  wire  _T_1717 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1745 = _T_1717 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1760 = _T_1759 | _T_1745; // @[Mux.scala 27:72]
  wire  _T_1720 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1746 = _T_1720 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1761 = _T_1760 | _T_1746; // @[Mux.scala 27:72]
  wire  _T_1723 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1747 = _T_1723 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1762 = _T_1761 | _T_1747; // @[Mux.scala 27:72]
  wire  _T_1726 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1748 = _T_1726 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1763 = _T_1762 | _T_1748; // @[Mux.scala 27:72]
  wire  _T_1729 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1749 = _T_1729 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1764 = _T_1763 | _T_1749; // @[Mux.scala 27:72]
  wire  _T_1732 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1750 = _T_1732 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1765 = _T_1764 | _T_1750; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1767 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1815 = _T_1767 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1770 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1816 = _T_1770 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1831 = _T_1815 | _T_1816; // @[Mux.scala 27:72]
  wire  _T_1773 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1817 = _T_1773 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1832 = _T_1831 | _T_1817; // @[Mux.scala 27:72]
  wire  _T_1776 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1818 = _T_1776 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1833 = _T_1832 | _T_1818; // @[Mux.scala 27:72]
  wire  _T_1779 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1819 = _T_1779 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1834 = _T_1833 | _T_1819; // @[Mux.scala 27:72]
  wire  _T_1782 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1820 = _T_1782 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1835 = _T_1834 | _T_1820; // @[Mux.scala 27:72]
  wire  _T_1785 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1821 = _T_1785 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1836 = _T_1835 | _T_1821; // @[Mux.scala 27:72]
  wire  _T_1788 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1822 = _T_1788 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1837 = _T_1836 | _T_1822; // @[Mux.scala 27:72]
  wire  _T_1791 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1823 = _T_1791 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1838 = _T_1837 | _T_1823; // @[Mux.scala 27:72]
  wire  _T_1794 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1824 = _T_1794 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1839 = _T_1838 | _T_1824; // @[Mux.scala 27:72]
  wire  _T_1797 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1825 = _T_1797 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1840 = _T_1839 | _T_1825; // @[Mux.scala 27:72]
  wire  _T_1800 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1826 = _T_1800 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1841 = _T_1840 | _T_1826; // @[Mux.scala 27:72]
  wire  _T_1803 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1827 = _T_1803 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1842 = _T_1841 | _T_1827; // @[Mux.scala 27:72]
  wire  _T_1806 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1828 = _T_1806 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1843 = _T_1842 | _T_1828; // @[Mux.scala 27:72]
  wire  _T_1809 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1829 = _T_1809 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1844 = _T_1843 | _T_1829; // @[Mux.scala 27:72]
  wire  _T_1812 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1830 = _T_1812 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1845 = _T_1844 | _T_1830; // @[Mux.scala 27:72]
  wire [79:0] _T_1848 = {_T_1685,_T_1765,_T_1845}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1849 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1897 = _T_1849 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1852 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1898 = _T_1852 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1913 = _T_1897 | _T_1898; // @[Mux.scala 27:72]
  wire  _T_1855 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1899 = _T_1855 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1914 = _T_1913 | _T_1899; // @[Mux.scala 27:72]
  wire  _T_1858 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1900 = _T_1858 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1915 = _T_1914 | _T_1900; // @[Mux.scala 27:72]
  wire  _T_1861 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1901 = _T_1861 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1916 = _T_1915 | _T_1901; // @[Mux.scala 27:72]
  wire  _T_1864 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1902 = _T_1864 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1917 = _T_1916 | _T_1902; // @[Mux.scala 27:72]
  wire  _T_1867 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1903 = _T_1867 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1918 = _T_1917 | _T_1903; // @[Mux.scala 27:72]
  wire  _T_1870 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1904 = _T_1870 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1919 = _T_1918 | _T_1904; // @[Mux.scala 27:72]
  wire  _T_1873 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1905 = _T_1873 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1920 = _T_1919 | _T_1905; // @[Mux.scala 27:72]
  wire  _T_1876 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1906 = _T_1876 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1921 = _T_1920 | _T_1906; // @[Mux.scala 27:72]
  wire  _T_1879 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1907 = _T_1879 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1922 = _T_1921 | _T_1907; // @[Mux.scala 27:72]
  wire  _T_1882 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1908 = _T_1882 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1923 = _T_1922 | _T_1908; // @[Mux.scala 27:72]
  wire  _T_1885 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1909 = _T_1885 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1924 = _T_1923 | _T_1909; // @[Mux.scala 27:72]
  wire  _T_1888 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1910 = _T_1888 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1925 = _T_1924 | _T_1910; // @[Mux.scala 27:72]
  wire  _T_1891 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1911 = _T_1891 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1926 = _T_1925 | _T_1911; // @[Mux.scala 27:72]
  wire  _T_1894 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1912 = _T_1894 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1927 = _T_1926 | _T_1912; // @[Mux.scala 27:72]
  wire [31:0] _T_1977 = _T_1607 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1978 = _T_1610 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1993 = _T_1977 | _T_1978; // @[Mux.scala 27:72]
  wire [31:0] _T_1979 = _T_1613 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1994 = _T_1993 | _T_1979; // @[Mux.scala 27:72]
  wire [31:0] _T_1980 = _T_1616 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1995 = _T_1994 | _T_1980; // @[Mux.scala 27:72]
  wire [31:0] _T_1981 = _T_1619 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1996 = _T_1995 | _T_1981; // @[Mux.scala 27:72]
  wire [31:0] _T_1982 = _T_1622 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1996 | _T_1982; // @[Mux.scala 27:72]
  wire [31:0] _T_1983 = _T_1625 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1997 | _T_1983; // @[Mux.scala 27:72]
  wire [31:0] _T_1984 = _T_1628 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1998 | _T_1984; // @[Mux.scala 27:72]
  wire [31:0] _T_1985 = _T_1631 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1999 | _T_1985; // @[Mux.scala 27:72]
  wire [31:0] _T_1986 = _T_1634 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_2000 | _T_1986; // @[Mux.scala 27:72]
  wire [31:0] _T_1987 = _T_1637 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_2001 | _T_1987; // @[Mux.scala 27:72]
  wire [31:0] _T_1988 = _T_1640 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_2002 | _T_1988; // @[Mux.scala 27:72]
  wire [31:0] _T_1989 = _T_1643 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_2003 | _T_1989; // @[Mux.scala 27:72]
  wire [31:0] _T_1990 = _T_1646 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_2004 | _T_1990; // @[Mux.scala 27:72]
  wire [31:0] _T_1991 = _T_1649 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_2005 | _T_1991; // @[Mux.scala 27:72]
  wire [31:0] _T_1992 = _T_1652 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_2006 | _T_1992; // @[Mux.scala 27:72]
  wire [79:0] _T_2090 = {_T_1927,_T_2007,_T_1765}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_2093 ? _T_1848 : _T_2090; // @[el2_ifu_mem_ctl.scala 431:37]
  wire [79:0] _T_2095 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2093 ? ic_byp_data_only_pre_new : _T_2095; // @[el2_ifu_mem_ctl.scala 435:30]
  wire [79:0] _GEN_793 = {{16'd0}, _T_1257}; // @[el2_ifu_mem_ctl.scala 366:109]
  wire [79:0] _T_1258 = _GEN_793 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 366:109]
  wire [79:0] _GEN_794 = {{16'd0}, _T_1255}; // @[el2_ifu_mem_ctl.scala 366:83]
  wire [79:0] ic_premux_data = _GEN_794 | _T_1258; // @[el2_ifu_mem_ctl.scala 366:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_309; // @[el2_ifu_mem_ctl.scala 373:38]
  wire [1:0] _T_1267 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 377:8]
  wire [7:0] _T_1348 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1353 = ic_miss_buff_data_error[0] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  _T_2602 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 608:47]
  wire  _T_2603 = _T_2602 & _T_14; // @[el2_ifu_mem_ctl.scala 608:50]
  wire  bus_ifu_wr_data_error = _T_2603 & miss_pending; // @[el2_ifu_mem_ctl.scala 608:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1353; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1357 = ic_miss_buff_data_error[1] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1357; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1361 = ic_miss_buff_data_error[2] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1361; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1365 = ic_miss_buff_data_error[3] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1365; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1369 = ic_miss_buff_data_error[4] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1369; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1373 = ic_miss_buff_data_error[5] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1373; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1377 = ic_miss_buff_data_error[6] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1377; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1381 = ic_miss_buff_data_error[7] & _T_1319; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1381; // @[el2_ifu_mem_ctl.scala 397:72]
  wire [7:0] _T_1388 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2410 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2418 = _T_7 & _T_309; // @[el2_ifu_mem_ctl.scala 478:65]
  wire  _T_2419 = _T_2418 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 478:88]
  wire  _T_2421 = _T_2419 & _T_2530; // @[el2_ifu_mem_ctl.scala 478:112]
  wire  _T_2422 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2423 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 483:50]
  wire  _T_2425 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2431 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2433 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2431 | _T_2433; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2425 ? _T_2423 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2422 ? _T_2423 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2410 ? _T_2421 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2410 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2424 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 484:56]
  wire  _GEN_43 = _T_2422 & _T_2424; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2410 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 469:58]
  wire  _T_2407 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 468:49]
  wire  _T_2412 = io_ic_error_start & _T_309; // @[el2_ifu_mem_ctl.scala 477:87]
  wire  _T_2426 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 487:54]
  wire  _T_2427 = _T_2426 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 487:84]
  wire  _T_2436 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 508:66]
  wire  _T_2437 = io_dec_tlu_flush_err_wb & _T_2436; // @[el2_ifu_mem_ctl.scala 508:52]
  wire  _T_2439 = _T_2437 & _T_2530; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2441 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 511:59]
  wire  _T_2442 = _T_2441 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 511:86]
  wire  _T_2456 = _T_2441 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 514:81]
  wire  _T_2457 = _T_2456 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 514:103]
  wire  _T_2458 = _T_2457 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 514:126]
  wire  _T_2478 = _T_2456 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 521:103]
  wire  _T_2485 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 526:62]
  wire  _T_2486 = io_dec_tlu_flush_lower_wb & _T_2485; // @[el2_ifu_mem_ctl.scala 526:60]
  wire  _T_2487 = _T_2486 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 526:88]
  wire  _T_2488 = _T_2487 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 526:115]
  wire  _GEN_50 = _T_2484 & _T_2442; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_2467 ? _T_2478 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_2467 | _T_2484; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_2440 ? _T_2458 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2440 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2435 ? _T_2439 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2498 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 542:64]
  wire  _T_2500 = _T_2498 & _T_2530; // @[el2_ifu_mem_ctl.scala 542:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2502 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 542:133]
  wire  _T_2503 = _T_2502 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 542:164]
  wire  _T_2504 = _T_2503 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 542:184]
  wire  _T_2505 = _T_2504 & miss_pending; // @[el2_ifu_mem_ctl.scala 542:204]
  wire  _T_2506 = ~_T_2505; // @[el2_ifu_mem_ctl.scala 542:112]
  wire  ifc_bus_ic_req_ff_in = _T_2500 & _T_2506; // @[el2_ifu_mem_ctl.scala 542:110]
  wire  _T_2507 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 543:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 574:45]
  wire  _T_2524 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 577:35]
  wire  _T_2525 = _T_2524 & miss_pending; // @[el2_ifu_mem_ctl.scala 577:53]
  wire  bus_cmd_sent = _T_2525 & _T_2530; // @[el2_ifu_mem_ctl.scala 577:68]
  wire [2:0] _T_2515 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2517 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2519 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 575:51]
  wire  _T_2548 = last_data_recieved_ff & _T_1319; // @[el2_ifu_mem_ctl.scala 585:114]
  wire  last_data_recieved_in = _T_2531 | _T_2548; // @[el2_ifu_mem_ctl.scala 585:89]
  wire [2:0] _T_2554 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 590:45]
  wire  _T_2557 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 591:81]
  wire  _T_2558 = _T_2557 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 591:97]
  wire  _T_2560 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 593:48]
  wire  _T_2561 = _T_2560 & miss_pending; // @[el2_ifu_mem_ctl.scala 593:68]
  wire  bus_inc_cmd_beat_cnt = _T_2561 & _T_2530; // @[el2_ifu_mem_ctl.scala 593:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 595:57]
  wire  _T_2565 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 596:31]
  wire  _T_2567 = ic_act_miss_f | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 596:87]
  wire  _T_2568 = ~_T_2567; // @[el2_ifu_mem_ctl.scala 596:55]
  wire  bus_hold_cmd_beat_cnt = _T_2565 & _T_2568; // @[el2_ifu_mem_ctl.scala 596:53]
  wire  _T_2569 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 597:46]
  wire  bus_cmd_beat_en = _T_2569 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 597:62]
  wire [2:0] _T_2572 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 599:46]
  wire [2:0] _T_2574 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2575 = bus_inc_cmd_beat_cnt ? _T_2572 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2576 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2578 = _T_2574 | _T_2575; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2578 | _T_2576; // @[Mux.scala 27:72]
  wire  _T_2582 = _T_2558 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 600:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 611:62]
  wire  _T_2610 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 616:50]
  wire  _T_2611 = io_ifc_dma_access_ok & _T_2610; // @[el2_ifu_mem_ctl.scala 616:47]
  wire  _T_2612 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 616:70]
  wire  ifc_dma_access_ok_d = _T_2611 & _T_2612; // @[el2_ifu_mem_ctl.scala 616:68]
  wire  _T_2616 = _T_2611 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 617:72]
  wire  _T_2617 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 617:111]
  wire  _T_2618 = _T_2616 & _T_2617; // @[el2_ifu_mem_ctl.scala 617:97]
  wire  ifc_dma_access_q_ok = _T_2618 & _T_2612; // @[el2_ifu_mem_ctl.scala 617:127]
  wire  _T_2621 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 620:40]
  wire  _T_2622 = _T_2621 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 620:58]
  wire  _T_2625 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 621:60]
  wire  _T_2626 = _T_2621 & _T_2625; // @[el2_ifu_mem_ctl.scala 621:58]
  wire  _T_2627 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 621:104]
  wire [2:0] _T_2632 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2738 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2747 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2738}; // @[el2_lib.scala 268:22]
  wire  _T_2748 = ^_T_2747; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2756 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2765 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2756}; // @[el2_lib.scala 268:39]
  wire  _T_2766 = ^_T_2765; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2774 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2783 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2774}; // @[el2_lib.scala 268:56]
  wire  _T_2784 = ^_T_2783; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2790 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2798 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2790}; // @[el2_lib.scala 268:73]
  wire  _T_2799 = ^_T_2798; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2813 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2790}; // @[el2_lib.scala 268:90]
  wire  _T_2814 = ^_T_2813; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2819 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2820 = ^_T_2819; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2825 = {_T_2748,_T_2766,_T_2784,_T_2799,_T_2814,_T_2820}; // @[Cat.scala 29:58]
  wire  _T_2826 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2827 = ^_T_2825; // @[el2_lib.scala 269:23]
  wire  _T_2828 = _T_2826 ^ _T_2827; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2934 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2943 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2934}; // @[el2_lib.scala 268:22]
  wire  _T_2944 = ^_T_2943; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2952 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2961 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2952}; // @[el2_lib.scala 268:39]
  wire  _T_2962 = ^_T_2961; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2970 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2979 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2970}; // @[el2_lib.scala 268:56]
  wire  _T_2980 = ^_T_2979; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2986 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2994 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2986}; // @[el2_lib.scala 268:73]
  wire  _T_2995 = ^_T_2994; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3009 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2986}; // @[el2_lib.scala 268:90]
  wire  _T_3010 = ^_T_3009; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3015 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3016 = ^_T_3015; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3021 = {_T_2944,_T_2962,_T_2980,_T_2995,_T_3010,_T_3016}; // @[Cat.scala 29:58]
  wire  _T_3022 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3023 = ^_T_3021; // @[el2_lib.scala 269:23]
  wire  _T_3024 = _T_3022 ^ _T_3023; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3025 = {_T_3024,_T_2944,_T_2962,_T_2980,_T_2995,_T_3010,_T_3016}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2828,_T_2748,_T_2766,_T_2784,_T_2799,_T_2814,_T_2820,_T_3025}; // @[Cat.scala 29:58]
  wire  _T_3027 = ~_T_2621; // @[el2_ifu_mem_ctl.scala 626:45]
  wire  _T_3028 = iccm_correct_ecc & _T_3027; // @[el2_ifu_mem_ctl.scala 626:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3029 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3036 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 640:53]
  wire  _T_3368 = _T_3280[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3366 = _T_3280[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3364 = _T_3280[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3362 = _T_3280[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3360 = _T_3280[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3358 = _T_3280[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3356 = _T_3280[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3354 = _T_3280[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3352 = _T_3280[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3350 = _T_3280[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3426 = {_T_3368,_T_3366,_T_3364,_T_3362,_T_3360,_T_3358,_T_3356,_T_3354,_T_3352,_T_3350}; // @[el2_lib.scala 310:69]
  wire  _T_3348 = _T_3280[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3346 = _T_3280[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3344 = _T_3280[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3342 = _T_3280[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3340 = _T_3280[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3338 = _T_3280[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3336 = _T_3280[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3334 = _T_3280[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3332 = _T_3280[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3330 = _T_3280[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3417 = {_T_3348,_T_3346,_T_3344,_T_3342,_T_3340,_T_3338,_T_3336,_T_3334,_T_3332,_T_3330}; // @[el2_lib.scala 310:69]
  wire  _T_3328 = _T_3280[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3326 = _T_3280[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3324 = _T_3280[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3322 = _T_3280[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3320 = _T_3280[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3318 = _T_3280[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3316 = _T_3280[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3314 = _T_3280[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3312 = _T_3280[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3310 = _T_3280[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3407 = {_T_3328,_T_3326,_T_3324,_T_3322,_T_3320,_T_3318,_T_3316,_T_3314,_T_3312,_T_3310}; // @[el2_lib.scala 310:69]
  wire  _T_3308 = _T_3280[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3306 = _T_3280[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3304 = _T_3280[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3302 = _T_3280[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3300 = _T_3280[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3298 = _T_3280[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3296 = _T_3280[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3294 = _T_3280[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3292 = _T_3280[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3408 = {_T_3407,_T_3308,_T_3306,_T_3304,_T_3302,_T_3300,_T_3298,_T_3296,_T_3294,_T_3292}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3428 = {_T_3426,_T_3417,_T_3408}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3383 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3389 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3383}; // @[Cat.scala 29:58]
  wire [38:0] _T_3429 = _T_3428 ^ _T_3389; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3430 = _T_3284 ? _T_3429 : _T_3389; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3430[37:32],_T_3430[30:16],_T_3430[14:8],_T_3430[6:4],_T_3430[2]}; // @[Cat.scala 29:58]
  wire  _T_3753 = _T_3665[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3751 = _T_3665[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3749 = _T_3665[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3747 = _T_3665[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3745 = _T_3665[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3743 = _T_3665[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3741 = _T_3665[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3739 = _T_3665[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3737 = _T_3665[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3735 = _T_3665[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3811 = {_T_3753,_T_3751,_T_3749,_T_3747,_T_3745,_T_3743,_T_3741,_T_3739,_T_3737,_T_3735}; // @[el2_lib.scala 310:69]
  wire  _T_3733 = _T_3665[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3731 = _T_3665[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3729 = _T_3665[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3727 = _T_3665[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3725 = _T_3665[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3723 = _T_3665[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3721 = _T_3665[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3719 = _T_3665[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3717 = _T_3665[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3715 = _T_3665[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3802 = {_T_3733,_T_3731,_T_3729,_T_3727,_T_3725,_T_3723,_T_3721,_T_3719,_T_3717,_T_3715}; // @[el2_lib.scala 310:69]
  wire  _T_3713 = _T_3665[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3711 = _T_3665[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3709 = _T_3665[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3707 = _T_3665[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3705 = _T_3665[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3703 = _T_3665[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3701 = _T_3665[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3699 = _T_3665[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3697 = _T_3665[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3695 = _T_3665[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3792 = {_T_3713,_T_3711,_T_3709,_T_3707,_T_3705,_T_3703,_T_3701,_T_3699,_T_3697,_T_3695}; // @[el2_lib.scala 310:69]
  wire  _T_3693 = _T_3665[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3691 = _T_3665[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3689 = _T_3665[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3687 = _T_3665[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3685 = _T_3665[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3683 = _T_3665[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3681 = _T_3665[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3679 = _T_3665[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3677 = _T_3665[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3793 = {_T_3792,_T_3693,_T_3691,_T_3689,_T_3687,_T_3685,_T_3683,_T_3681,_T_3679,_T_3677}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3813 = {_T_3811,_T_3802,_T_3793}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3768 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3774 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3768}; // @[Cat.scala 29:58]
  wire [38:0] _T_3814 = _T_3813 ^ _T_3774; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3815 = _T_3669 ? _T_3814 : _T_3774; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3815[37:32],_T_3815[30:16],_T_3815[14:8],_T_3815[6:4],_T_3815[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 632:35]
  wire  _T_3288 = ~_T_3280[6]; // @[el2_lib.scala 303:55]
  wire  _T_3289 = _T_3282 & _T_3288; // @[el2_lib.scala 303:53]
  wire  _T_3673 = ~_T_3665[6]; // @[el2_lib.scala 303:55]
  wire  _T_3674 = _T_3667 & _T_3673; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3289,_T_3674}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 634:53]
  wire [63:0] _T_3040 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3041 = {iccm_dma_rdata_1_muxed,_T_3430[37:32],_T_3430[30:16],_T_3430[14:8],_T_3430[6:4],_T_3430[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 636:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 637:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 642:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 646:70]
  wire  _T_3046 = _T_2621 & _T_2610; // @[el2_ifu_mem_ctl.scala 649:65]
  wire  _T_3049 = _T_3027 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 650:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3050 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3052 = _T_3049 ? {{1'd0}, _T_3050} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 650:8]
  wire [31:0] _T_3053 = _T_3046 ? io_dma_mem_addr : {{16'd0}, _T_3052}; // @[el2_ifu_mem_ctl.scala 649:25]
  wire  _T_3442 = _T_3280 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3443 = _T_3430[38] ^ _T_3442; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3443,_T_3430[31],_T_3430[15],_T_3430[7],_T_3430[3],_T_3430[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3827 = _T_3665 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3828 = _T_3815[38] ^ _T_3827; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3828,_T_3815[31],_T_3815[15],_T_3815[7],_T_3815[3],_T_3815[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3844 = _T_4 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 662:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 664:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 665:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 673:62]
  wire  _T_3852 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 667:76]
  wire  _T_3853 = io_iccm_rd_ecc_single_err & _T_3852; // @[el2_ifu_mem_ctl.scala 667:74]
  wire  _T_3855 = _T_3853 & _T_309; // @[el2_ifu_mem_ctl.scala 667:104]
  wire  iccm_ecc_write_status = _T_3855 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 667:127]
  wire  _T_3856 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 668:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3856 & _T_309; // @[el2_ifu_mem_ctl.scala 668:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 672:51]
  wire [13:0] _T_3861 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 671:102]
  wire [38:0] _T_3865 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3870 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 676:41]
  wire  _T_3871 = io_ifc_fetch_req_bf & _T_3870; // @[el2_ifu_mem_ctl.scala 676:39]
  wire  _T_3872 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 676:72]
  wire  _T_3873 = _T_3871 & _T_3872; // @[el2_ifu_mem_ctl.scala 676:70]
  wire  _T_3875 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 677:34]
  wire  _T_3876 = _T_2219 & _T_3875; // @[el2_ifu_mem_ctl.scala 677:32]
  wire  _T_3879 = _T_2234 & _T_3875; // @[el2_ifu_mem_ctl.scala 678:37]
  wire  _T_3880 = _T_3876 | _T_3879; // @[el2_ifu_mem_ctl.scala 677:88]
  wire  _T_3881 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 679:19]
  wire  _T_3883 = _T_3881 & _T_3875; // @[el2_ifu_mem_ctl.scala 679:41]
  wire  _T_3884 = _T_3880 | _T_3883; // @[el2_ifu_mem_ctl.scala 678:88]
  wire  _T_3885 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 680:19]
  wire  _T_3887 = _T_3885 & _T_3875; // @[el2_ifu_mem_ctl.scala 680:35]
  wire  _T_3888 = _T_3884 | _T_3887; // @[el2_ifu_mem_ctl.scala 679:88]
  wire  _T_3891 = _T_2233 & _T_3875; // @[el2_ifu_mem_ctl.scala 681:38]
  wire  _T_3892 = _T_3888 | _T_3891; // @[el2_ifu_mem_ctl.scala 680:88]
  wire  _T_3894 = _T_2234 & miss_state_en; // @[el2_ifu_mem_ctl.scala 682:37]
  wire  _T_3895 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 682:71]
  wire  _T_3896 = _T_3894 & _T_3895; // @[el2_ifu_mem_ctl.scala 682:54]
  wire  _T_3897 = _T_3892 | _T_3896; // @[el2_ifu_mem_ctl.scala 681:57]
  wire  _T_3898 = ~_T_3897; // @[el2_ifu_mem_ctl.scala 677:5]
  wire  _T_3899 = _T_3873 & _T_3898; // @[el2_ifu_mem_ctl.scala 676:96]
  wire  _T_3900 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 683:28]
  wire  _T_3902 = _T_3900 & _T_3870; // @[el2_ifu_mem_ctl.scala 683:50]
  wire  _T_3904 = _T_3902 & _T_3872; // @[el2_ifu_mem_ctl.scala 683:81]
  wire  _T_3913 = ~_T_100; // @[el2_ifu_mem_ctl.scala 686:106]
  wire  _T_3914 = _T_2219 & _T_3913; // @[el2_ifu_mem_ctl.scala 686:104]
  wire  _T_3915 = _T_2234 | _T_3914; // @[el2_ifu_mem_ctl.scala 686:77]
  wire  _T_3919 = ~_T_53; // @[el2_ifu_mem_ctl.scala 686:172]
  wire  _T_3920 = _T_3915 & _T_3919; // @[el2_ifu_mem_ctl.scala 686:170]
  wire  _T_3921 = ~_T_3920; // @[el2_ifu_mem_ctl.scala 686:44]
  wire  _T_3925 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 689:64]
  wire  _T_3926 = ~_T_3925; // @[el2_ifu_mem_ctl.scala 689:50]
  wire  _T_3927 = _T_268 & _T_3926; // @[el2_ifu_mem_ctl.scala 689:48]
  wire  _T_3928 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 689:81]
  wire  ic_valid = _T_3927 & _T_3928; // @[el2_ifu_mem_ctl.scala 689:79]
  wire  _T_3930 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 690:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 693:14]
  wire  _T_3933 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 696:74]
  wire  _T_9443 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 774:45]
  wire  way_status_wr_en = _T_9443 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 774:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3933; // @[el2_ifu_mem_ctl.scala 696:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 698:14]
  wire [2:0] _T_3937 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 702:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 770:41]
  wire  way_status_new = _T_9443 | way_status_hit_new; // @[el2_ifu_mem_ctl.scala 773:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 704:14]
  wire  _T_3954 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3955 = _T_3954 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_3957 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3958 = _T_3957 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_3960 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3961 = _T_3960 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_3963 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3964 = _T_3963 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_3966 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3967 = _T_3966 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_3969 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3970 = _T_3969 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_3972 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3973 = _T_3972 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_3975 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 711:65]
  wire  _T_3976 = _T_3975 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:73]
  wire  _T_9448 = _T_92 & miss_pending; // @[el2_ifu_mem_ctl.scala 777:108]
  wire  bus_wren_last_0 = _T_9448 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 777:123]
  wire  _T_9451 = bus_wren_last_0 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 779:73]
  wire [1:0] ifu_tag_wren = {1'h0,_T_9451}; // @[Cat.scala 29:58]
  wire [1:0] _T_9486 = _T_3933 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9486 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 810:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 721:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 723:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 727:14]
  wire  _T_4985 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 731:82]
  wire  _T_4987 = _T_4985 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_4989 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 732:74]
  wire  _T_4991 = _T_4989 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_4992 = _T_4987 | _T_4991; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_4993 = _T_4992 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire  _T_4997 = _T_4985 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_5001 = _T_4989 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_5002 = _T_4997 | _T_5001; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_5003 = _T_5002 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire [1:0] tag_valid_clken_0 = {_T_4993,_T_5003}; // @[Cat.scala 29:58]
  wire  _T_5005 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 731:82]
  wire  _T_5007 = _T_5005 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_5009 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 732:74]
  wire  _T_5011 = _T_5009 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_5012 = _T_5007 | _T_5011; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_5013 = _T_5012 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire  _T_5017 = _T_5005 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_5021 = _T_5009 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_5022 = _T_5017 | _T_5021; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_5023 = _T_5022 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire [1:0] tag_valid_clken_1 = {_T_5013,_T_5023}; // @[Cat.scala 29:58]
  wire  _T_5025 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 731:82]
  wire  _T_5027 = _T_5025 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_5029 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 732:74]
  wire  _T_5031 = _T_5029 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_5032 = _T_5027 | _T_5031; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_5033 = _T_5032 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire  _T_5037 = _T_5025 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_5041 = _T_5029 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_5042 = _T_5037 | _T_5041; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_5043 = _T_5042 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire [1:0] tag_valid_clken_2 = {_T_5033,_T_5043}; // @[Cat.scala 29:58]
  wire  _T_5045 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 731:82]
  wire  _T_5047 = _T_5045 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_5049 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 732:74]
  wire  _T_5051 = _T_5049 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_5052 = _T_5047 | _T_5051; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_5053 = _T_5052 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire  _T_5057 = _T_5045 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 731:91]
  wire  _T_5061 = _T_5049 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 732:83]
  wire  _T_5062 = _T_5057 | _T_5061; // @[el2_ifu_mem_ctl.scala 731:113]
  wire  _T_5063 = _T_5062 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 732:106]
  wire [1:0] tag_valid_clken_3 = {_T_5053,_T_5063}; // @[Cat.scala 29:58]
  wire  _T_5074 = ic_valid_ff & _T_187; // @[el2_ifu_mem_ctl.scala 738:31]
  wire  _T_5075 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 738:58]
  wire  _T_5076 = _T_5074 & _T_5075; // @[el2_ifu_mem_ctl.scala 738:56]
  wire  _T_5079 = _T_4338 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5080 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5082 = _T_5080 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5083 = _T_5079 | _T_5082; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5093 = _T_4342 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5094 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5096 = _T_5094 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5097 = _T_5093 | _T_5096; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5107 = _T_4346 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5108 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5110 = _T_5108 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5111 = _T_5107 | _T_5110; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5121 = _T_4350 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5122 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5124 = _T_5122 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5125 = _T_5121 | _T_5124; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5135 = _T_4354 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5136 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5138 = _T_5136 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5139 = _T_5135 | _T_5138; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5149 = _T_4358 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5150 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5152 = _T_5150 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5153 = _T_5149 | _T_5152; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5163 = _T_4362 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5164 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5166 = _T_5164 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5167 = _T_5163 | _T_5166; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5177 = _T_4366 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5178 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5180 = _T_5178 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5181 = _T_5177 | _T_5180; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5191 = _T_4370 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5192 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5194 = _T_5192 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5195 = _T_5191 | _T_5194; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5205 = _T_4374 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5206 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5208 = _T_5206 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5209 = _T_5205 | _T_5208; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5219 = _T_4378 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5220 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5222 = _T_5220 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5223 = _T_5219 | _T_5222; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5233 = _T_4382 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5234 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5236 = _T_5234 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5237 = _T_5233 | _T_5236; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5247 = _T_4386 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5248 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5250 = _T_5248 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5251 = _T_5247 | _T_5250; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5261 = _T_4390 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5262 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5264 = _T_5262 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5265 = _T_5261 | _T_5264; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5275 = _T_4394 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5276 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5278 = _T_5276 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5279 = _T_5275 | _T_5278; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5289 = _T_4398 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5290 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5292 = _T_5290 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5293 = _T_5289 | _T_5292; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5303 = _T_4402 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5304 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5306 = _T_5304 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5307 = _T_5303 | _T_5306; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5317 = _T_4406 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5318 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5320 = _T_5318 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5321 = _T_5317 | _T_5320; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5331 = _T_4410 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5332 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5334 = _T_5332 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5335 = _T_5331 | _T_5334; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5345 = _T_4414 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5346 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5348 = _T_5346 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5349 = _T_5345 | _T_5348; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5359 = _T_4418 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5360 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5362 = _T_5360 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5363 = _T_5359 | _T_5362; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5373 = _T_4422 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5374 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5376 = _T_5374 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5377 = _T_5373 | _T_5376; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5387 = _T_4426 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5388 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5390 = _T_5388 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5391 = _T_5387 | _T_5390; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5401 = _T_4430 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5402 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5404 = _T_5402 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5405 = _T_5401 | _T_5404; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5415 = _T_4434 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5416 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5418 = _T_5416 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5419 = _T_5415 | _T_5418; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5429 = _T_4438 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5430 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5432 = _T_5430 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5433 = _T_5429 | _T_5432; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5443 = _T_4442 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5444 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5446 = _T_5444 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5447 = _T_5443 | _T_5446; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5457 = _T_4446 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5458 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5460 = _T_5458 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5461 = _T_5457 | _T_5460; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5471 = _T_4450 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5472 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5474 = _T_5472 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5475 = _T_5471 | _T_5474; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5485 = _T_4454 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5486 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5488 = _T_5486 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5489 = _T_5485 | _T_5488; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5499 = _T_4458 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5500 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5502 = _T_5500 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5503 = _T_5499 | _T_5502; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5513 = _T_4462 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5514 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5516 = _T_5514 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5517 = _T_5513 | _T_5516; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5527 = _T_4338 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5530 = _T_5080 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5531 = _T_5527 | _T_5530; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5541 = _T_4342 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5544 = _T_5094 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5545 = _T_5541 | _T_5544; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5555 = _T_4346 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5558 = _T_5108 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5559 = _T_5555 | _T_5558; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5569 = _T_4350 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5572 = _T_5122 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5573 = _T_5569 | _T_5572; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5583 = _T_4354 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5586 = _T_5136 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5587 = _T_5583 | _T_5586; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5597 = _T_4358 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5600 = _T_5150 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5601 = _T_5597 | _T_5600; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5611 = _T_4362 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5614 = _T_5164 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5615 = _T_5611 | _T_5614; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5625 = _T_4366 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5628 = _T_5178 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5629 = _T_5625 | _T_5628; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5639 = _T_4370 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5642 = _T_5192 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5643 = _T_5639 | _T_5642; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5653 = _T_4374 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5656 = _T_5206 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5657 = _T_5653 | _T_5656; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5667 = _T_4378 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5670 = _T_5220 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5671 = _T_5667 | _T_5670; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5681 = _T_4382 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5684 = _T_5234 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5685 = _T_5681 | _T_5684; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5695 = _T_4386 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5698 = _T_5248 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5699 = _T_5695 | _T_5698; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5709 = _T_4390 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5712 = _T_5262 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5713 = _T_5709 | _T_5712; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5723 = _T_4394 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5726 = _T_5276 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5727 = _T_5723 | _T_5726; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5737 = _T_4398 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5740 = _T_5290 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5741 = _T_5737 | _T_5740; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5751 = _T_4402 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5754 = _T_5304 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5755 = _T_5751 | _T_5754; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5765 = _T_4406 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5768 = _T_5318 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5769 = _T_5765 | _T_5768; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5779 = _T_4410 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5782 = _T_5332 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5783 = _T_5779 | _T_5782; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5793 = _T_4414 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5796 = _T_5346 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5797 = _T_5793 | _T_5796; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5807 = _T_4418 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5810 = _T_5360 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5811 = _T_5807 | _T_5810; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5821 = _T_4422 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5824 = _T_5374 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5825 = _T_5821 | _T_5824; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5835 = _T_4426 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5838 = _T_5388 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5839 = _T_5835 | _T_5838; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5849 = _T_4430 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5852 = _T_5402 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5853 = _T_5849 | _T_5852; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5863 = _T_4434 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5866 = _T_5416 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5867 = _T_5863 | _T_5866; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5877 = _T_4438 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5880 = _T_5430 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5881 = _T_5877 | _T_5880; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5891 = _T_4442 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5894 = _T_5444 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5895 = _T_5891 | _T_5894; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5905 = _T_4446 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5908 = _T_5458 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5909 = _T_5905 | _T_5908; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5919 = _T_4450 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5922 = _T_5472 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5923 = _T_5919 | _T_5922; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5933 = _T_4454 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5936 = _T_5486 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5937 = _T_5933 | _T_5936; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5947 = _T_4458 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5950 = _T_5500 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5951 = _T_5947 | _T_5950; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5961 = _T_4462 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5964 = _T_5514 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5965 = _T_5961 | _T_5964; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5975 = _T_4466 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5976 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5978 = _T_5976 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5979 = _T_5975 | _T_5978; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_5989 = _T_4470 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_5990 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_5992 = _T_5990 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_5993 = _T_5989 | _T_5992; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6003 = _T_4474 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6004 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6006 = _T_6004 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6007 = _T_6003 | _T_6006; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6017 = _T_4478 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6018 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6020 = _T_6018 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6021 = _T_6017 | _T_6020; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6031 = _T_4482 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6032 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6034 = _T_6032 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6035 = _T_6031 | _T_6034; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6045 = _T_4486 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6046 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6048 = _T_6046 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6049 = _T_6045 | _T_6048; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6059 = _T_4490 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6060 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6062 = _T_6060 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6063 = _T_6059 | _T_6062; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6073 = _T_4494 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6074 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6076 = _T_6074 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6077 = _T_6073 | _T_6076; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6087 = _T_4498 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6088 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6090 = _T_6088 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6091 = _T_6087 | _T_6090; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6101 = _T_4502 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6102 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6104 = _T_6102 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6105 = _T_6101 | _T_6104; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6115 = _T_4506 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6116 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6118 = _T_6116 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6119 = _T_6115 | _T_6118; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6129 = _T_4510 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6130 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6132 = _T_6130 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6133 = _T_6129 | _T_6132; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6143 = _T_4514 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6144 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6146 = _T_6144 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6147 = _T_6143 | _T_6146; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6157 = _T_4518 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6158 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6160 = _T_6158 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6161 = _T_6157 | _T_6160; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6171 = _T_4522 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6172 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6174 = _T_6172 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6175 = _T_6171 | _T_6174; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6185 = _T_4526 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6186 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6188 = _T_6186 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6189 = _T_6185 | _T_6188; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6199 = _T_4530 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6200 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6202 = _T_6200 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6203 = _T_6199 | _T_6202; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6213 = _T_4534 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6214 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6216 = _T_6214 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6217 = _T_6213 | _T_6216; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6227 = _T_4538 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6228 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6230 = _T_6228 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6231 = _T_6227 | _T_6230; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6241 = _T_4542 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6242 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6244 = _T_6242 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6245 = _T_6241 | _T_6244; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6255 = _T_4546 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6256 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6258 = _T_6256 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6259 = _T_6255 | _T_6258; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6269 = _T_4550 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6270 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6272 = _T_6270 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6273 = _T_6269 | _T_6272; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6283 = _T_4554 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6284 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6286 = _T_6284 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6287 = _T_6283 | _T_6286; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6297 = _T_4558 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6298 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6300 = _T_6298 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6301 = _T_6297 | _T_6300; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6311 = _T_4562 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6312 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6314 = _T_6312 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6315 = _T_6311 | _T_6314; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6325 = _T_4566 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6326 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6328 = _T_6326 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6329 = _T_6325 | _T_6328; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6339 = _T_4570 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6340 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6342 = _T_6340 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6343 = _T_6339 | _T_6342; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6353 = _T_4574 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6354 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6356 = _T_6354 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6357 = _T_6353 | _T_6356; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6367 = _T_4578 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6368 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6370 = _T_6368 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6371 = _T_6367 | _T_6370; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6381 = _T_4582 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6382 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6384 = _T_6382 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6385 = _T_6381 | _T_6384; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6395 = _T_4586 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6396 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6398 = _T_6396 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6399 = _T_6395 | _T_6398; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6409 = _T_4590 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6410 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6412 = _T_6410 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6413 = _T_6409 | _T_6412; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6423 = _T_4466 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6426 = _T_5976 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6427 = _T_6423 | _T_6426; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6437 = _T_4470 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6440 = _T_5990 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6441 = _T_6437 | _T_6440; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6451 = _T_4474 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6454 = _T_6004 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6455 = _T_6451 | _T_6454; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6465 = _T_4478 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6468 = _T_6018 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6469 = _T_6465 | _T_6468; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6479 = _T_4482 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6482 = _T_6032 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6483 = _T_6479 | _T_6482; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6493 = _T_4486 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6496 = _T_6046 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6497 = _T_6493 | _T_6496; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6507 = _T_4490 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6510 = _T_6060 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6511 = _T_6507 | _T_6510; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6521 = _T_4494 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6524 = _T_6074 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6525 = _T_6521 | _T_6524; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6535 = _T_4498 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6538 = _T_6088 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6539 = _T_6535 | _T_6538; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6549 = _T_4502 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6552 = _T_6102 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6553 = _T_6549 | _T_6552; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6563 = _T_4506 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6566 = _T_6116 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6567 = _T_6563 | _T_6566; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6577 = _T_4510 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6580 = _T_6130 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6581 = _T_6577 | _T_6580; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6591 = _T_4514 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6594 = _T_6144 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6595 = _T_6591 | _T_6594; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6605 = _T_4518 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6608 = _T_6158 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6609 = _T_6605 | _T_6608; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6619 = _T_4522 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6622 = _T_6172 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6623 = _T_6619 | _T_6622; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6633 = _T_4526 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6636 = _T_6186 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6637 = _T_6633 | _T_6636; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6647 = _T_4530 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6650 = _T_6200 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6651 = _T_6647 | _T_6650; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6661 = _T_4534 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6664 = _T_6214 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6665 = _T_6661 | _T_6664; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6675 = _T_4538 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6678 = _T_6228 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6679 = _T_6675 | _T_6678; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6689 = _T_4542 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6692 = _T_6242 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6693 = _T_6689 | _T_6692; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6703 = _T_4546 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6706 = _T_6256 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6707 = _T_6703 | _T_6706; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6717 = _T_4550 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6720 = _T_6270 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6721 = _T_6717 | _T_6720; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6731 = _T_4554 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6734 = _T_6284 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6735 = _T_6731 | _T_6734; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6745 = _T_4558 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6748 = _T_6298 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6749 = _T_6745 | _T_6748; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6759 = _T_4562 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6762 = _T_6312 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6763 = _T_6759 | _T_6762; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6773 = _T_4566 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6776 = _T_6326 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6777 = _T_6773 | _T_6776; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6787 = _T_4570 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6790 = _T_6340 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6791 = _T_6787 | _T_6790; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6801 = _T_4574 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6804 = _T_6354 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6805 = _T_6801 | _T_6804; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6815 = _T_4578 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6818 = _T_6368 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6819 = _T_6815 | _T_6818; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6829 = _T_4582 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6832 = _T_6382 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6833 = _T_6829 | _T_6832; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6843 = _T_4586 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6846 = _T_6396 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6847 = _T_6843 | _T_6846; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6857 = _T_4590 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6860 = _T_6410 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6861 = _T_6857 | _T_6860; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6871 = _T_4594 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6872 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6874 = _T_6872 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6875 = _T_6871 | _T_6874; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6885 = _T_4598 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6886 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6888 = _T_6886 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6889 = _T_6885 | _T_6888; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6899 = _T_4602 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6900 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6902 = _T_6900 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6903 = _T_6899 | _T_6902; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6913 = _T_4606 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6914 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6916 = _T_6914 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6917 = _T_6913 | _T_6916; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6927 = _T_4610 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6928 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6930 = _T_6928 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6931 = _T_6927 | _T_6930; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6941 = _T_4614 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6942 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6944 = _T_6942 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6945 = _T_6941 | _T_6944; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6955 = _T_4618 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6956 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6958 = _T_6956 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6959 = _T_6955 | _T_6958; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6969 = _T_4622 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6970 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6972 = _T_6970 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6973 = _T_6969 | _T_6972; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6983 = _T_4626 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6984 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_6986 = _T_6984 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_6987 = _T_6983 | _T_6986; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_6997 = _T_4630 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_6998 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7000 = _T_6998 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7001 = _T_6997 | _T_7000; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7011 = _T_4634 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7012 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7014 = _T_7012 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7015 = _T_7011 | _T_7014; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7025 = _T_4638 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7026 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7028 = _T_7026 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7029 = _T_7025 | _T_7028; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7039 = _T_4642 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7040 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7042 = _T_7040 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7043 = _T_7039 | _T_7042; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7053 = _T_4646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7054 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7056 = _T_7054 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7057 = _T_7053 | _T_7056; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7067 = _T_4650 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7068 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7070 = _T_7068 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7071 = _T_7067 | _T_7070; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7081 = _T_4654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7082 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7084 = _T_7082 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7085 = _T_7081 | _T_7084; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7095 = _T_4658 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7096 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7098 = _T_7096 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7099 = _T_7095 | _T_7098; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7109 = _T_4662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7110 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7112 = _T_7110 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7113 = _T_7109 | _T_7112; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7123 = _T_4666 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7124 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7126 = _T_7124 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7127 = _T_7123 | _T_7126; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7137 = _T_4670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7138 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7140 = _T_7138 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7141 = _T_7137 | _T_7140; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7151 = _T_4674 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7152 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7154 = _T_7152 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7155 = _T_7151 | _T_7154; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7165 = _T_4678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7166 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7168 = _T_7166 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7169 = _T_7165 | _T_7168; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7179 = _T_4682 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7180 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7182 = _T_7180 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7183 = _T_7179 | _T_7182; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7193 = _T_4686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7194 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7196 = _T_7194 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7197 = _T_7193 | _T_7196; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7207 = _T_4690 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7208 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7210 = _T_7208 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7211 = _T_7207 | _T_7210; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7221 = _T_4694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7222 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7224 = _T_7222 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7225 = _T_7221 | _T_7224; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7235 = _T_4698 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7236 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7238 = _T_7236 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7239 = _T_7235 | _T_7238; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7249 = _T_4702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7250 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7252 = _T_7250 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7253 = _T_7249 | _T_7252; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7263 = _T_4706 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7264 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7266 = _T_7264 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7267 = _T_7263 | _T_7266; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7277 = _T_4710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7278 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7280 = _T_7278 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7281 = _T_7277 | _T_7280; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7291 = _T_4714 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7292 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7294 = _T_7292 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7295 = _T_7291 | _T_7294; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7305 = _T_4718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7306 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7308 = _T_7306 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7309 = _T_7305 | _T_7308; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7319 = _T_4594 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7322 = _T_6872 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7323 = _T_7319 | _T_7322; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7333 = _T_4598 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7336 = _T_6886 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7337 = _T_7333 | _T_7336; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7347 = _T_4602 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7350 = _T_6900 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7351 = _T_7347 | _T_7350; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7361 = _T_4606 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7364 = _T_6914 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7365 = _T_7361 | _T_7364; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7375 = _T_4610 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7378 = _T_6928 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7379 = _T_7375 | _T_7378; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7389 = _T_4614 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7392 = _T_6942 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7393 = _T_7389 | _T_7392; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7403 = _T_4618 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7406 = _T_6956 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7407 = _T_7403 | _T_7406; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7417 = _T_4622 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7420 = _T_6970 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7421 = _T_7417 | _T_7420; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7431 = _T_4626 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7434 = _T_6984 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7435 = _T_7431 | _T_7434; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7445 = _T_4630 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7448 = _T_6998 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7449 = _T_7445 | _T_7448; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7459 = _T_4634 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7462 = _T_7012 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7463 = _T_7459 | _T_7462; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7473 = _T_4638 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7476 = _T_7026 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7477 = _T_7473 | _T_7476; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7487 = _T_4642 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7490 = _T_7040 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7491 = _T_7487 | _T_7490; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7501 = _T_4646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7504 = _T_7054 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7505 = _T_7501 | _T_7504; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7515 = _T_4650 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7518 = _T_7068 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7519 = _T_7515 | _T_7518; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7529 = _T_4654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7532 = _T_7082 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7533 = _T_7529 | _T_7532; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7543 = _T_4658 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7546 = _T_7096 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7547 = _T_7543 | _T_7546; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7557 = _T_4662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7560 = _T_7110 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7561 = _T_7557 | _T_7560; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7571 = _T_4666 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7574 = _T_7124 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7575 = _T_7571 | _T_7574; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7585 = _T_4670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7588 = _T_7138 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7589 = _T_7585 | _T_7588; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7599 = _T_4674 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7602 = _T_7152 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7603 = _T_7599 | _T_7602; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7613 = _T_4678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7616 = _T_7166 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7617 = _T_7613 | _T_7616; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7627 = _T_4682 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7630 = _T_7180 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7631 = _T_7627 | _T_7630; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7641 = _T_4686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7644 = _T_7194 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7645 = _T_7641 | _T_7644; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7655 = _T_4690 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7658 = _T_7208 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7659 = _T_7655 | _T_7658; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7669 = _T_4694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7672 = _T_7222 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7673 = _T_7669 | _T_7672; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7683 = _T_4698 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7686 = _T_7236 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7687 = _T_7683 | _T_7686; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7697 = _T_4702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7700 = _T_7250 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7701 = _T_7697 | _T_7700; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7711 = _T_4706 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7714 = _T_7264 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7715 = _T_7711 | _T_7714; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7725 = _T_4710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7728 = _T_7278 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7729 = _T_7725 | _T_7728; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7739 = _T_4714 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7742 = _T_7292 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7743 = _T_7739 | _T_7742; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7753 = _T_4718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7756 = _T_7306 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7757 = _T_7753 | _T_7756; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7767 = _T_4722 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7768 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7770 = _T_7768 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7771 = _T_7767 | _T_7770; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7781 = _T_4726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7782 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7784 = _T_7782 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7785 = _T_7781 | _T_7784; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7795 = _T_4730 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7796 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7798 = _T_7796 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7799 = _T_7795 | _T_7798; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7809 = _T_4734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7810 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7812 = _T_7810 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7813 = _T_7809 | _T_7812; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7823 = _T_4738 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7824 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7826 = _T_7824 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7827 = _T_7823 | _T_7826; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7837 = _T_4742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7838 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7840 = _T_7838 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7841 = _T_7837 | _T_7840; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7851 = _T_4746 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7852 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7854 = _T_7852 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7855 = _T_7851 | _T_7854; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7865 = _T_4750 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7866 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7868 = _T_7866 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7869 = _T_7865 | _T_7868; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7879 = _T_4754 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7880 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7882 = _T_7880 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7883 = _T_7879 | _T_7882; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7893 = _T_4758 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7894 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7896 = _T_7894 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7897 = _T_7893 | _T_7896; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7907 = _T_4762 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7908 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7910 = _T_7908 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7911 = _T_7907 | _T_7910; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7921 = _T_4766 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7922 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7924 = _T_7922 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7925 = _T_7921 | _T_7924; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7935 = _T_4770 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7936 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7938 = _T_7936 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7939 = _T_7935 | _T_7938; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7949 = _T_4774 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7950 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7952 = _T_7950 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7953 = _T_7949 | _T_7952; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7963 = _T_4778 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7964 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7966 = _T_7964 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7967 = _T_7963 | _T_7966; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7977 = _T_4782 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7978 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7980 = _T_7978 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7981 = _T_7977 | _T_7980; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_7991 = _T_4786 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_7992 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_7994 = _T_7992 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_7995 = _T_7991 | _T_7994; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8005 = _T_4790 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8006 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8008 = _T_8006 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8009 = _T_8005 | _T_8008; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8019 = _T_4794 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8020 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8022 = _T_8020 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8023 = _T_8019 | _T_8022; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8033 = _T_4798 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8034 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8036 = _T_8034 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8037 = _T_8033 | _T_8036; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8047 = _T_4802 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8048 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8050 = _T_8048 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8051 = _T_8047 | _T_8050; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8061 = _T_4806 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8062 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8064 = _T_8062 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8065 = _T_8061 | _T_8064; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8075 = _T_4810 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8076 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8078 = _T_8076 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8079 = _T_8075 | _T_8078; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8089 = _T_4814 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8090 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8092 = _T_8090 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8093 = _T_8089 | _T_8092; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8103 = _T_4818 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8104 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8106 = _T_8104 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8107 = _T_8103 | _T_8106; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8117 = _T_4822 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8118 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8120 = _T_8118 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8121 = _T_8117 | _T_8120; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8131 = _T_4826 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8132 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8134 = _T_8132 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8135 = _T_8131 | _T_8134; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8145 = _T_4830 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8146 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8148 = _T_8146 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8149 = _T_8145 | _T_8148; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8159 = _T_4834 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8160 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8162 = _T_8160 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8163 = _T_8159 | _T_8162; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8173 = _T_4838 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8174 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8176 = _T_8174 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8177 = _T_8173 | _T_8176; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8187 = _T_4842 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8188 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8190 = _T_8188 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8191 = _T_8187 | _T_8190; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8201 = _T_4846 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8202 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 739:101]
  wire  _T_8204 = _T_8202 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8205 = _T_8201 | _T_8204; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8215 = _T_4722 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8218 = _T_7768 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8219 = _T_8215 | _T_8218; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8229 = _T_4726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8232 = _T_7782 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8233 = _T_8229 | _T_8232; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8243 = _T_4730 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8246 = _T_7796 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8247 = _T_8243 | _T_8246; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8257 = _T_4734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8260 = _T_7810 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8261 = _T_8257 | _T_8260; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8271 = _T_4738 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8274 = _T_7824 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8275 = _T_8271 | _T_8274; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8285 = _T_4742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8288 = _T_7838 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8289 = _T_8285 | _T_8288; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8299 = _T_4746 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8302 = _T_7852 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8303 = _T_8299 | _T_8302; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8313 = _T_4750 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8316 = _T_7866 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8317 = _T_8313 | _T_8316; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8327 = _T_4754 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8330 = _T_7880 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8331 = _T_8327 | _T_8330; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8341 = _T_4758 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8344 = _T_7894 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8345 = _T_8341 | _T_8344; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8355 = _T_4762 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8358 = _T_7908 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8359 = _T_8355 | _T_8358; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8369 = _T_4766 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8372 = _T_7922 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8373 = _T_8369 | _T_8372; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8383 = _T_4770 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8386 = _T_7936 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8387 = _T_8383 | _T_8386; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8397 = _T_4774 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8400 = _T_7950 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8401 = _T_8397 | _T_8400; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8411 = _T_4778 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8414 = _T_7964 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8415 = _T_8411 | _T_8414; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8425 = _T_4782 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8428 = _T_7978 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8429 = _T_8425 | _T_8428; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8439 = _T_4786 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8442 = _T_7992 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8443 = _T_8439 | _T_8442; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8453 = _T_4790 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8456 = _T_8006 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8457 = _T_8453 | _T_8456; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8467 = _T_4794 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8470 = _T_8020 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8471 = _T_8467 | _T_8470; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8481 = _T_4798 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8484 = _T_8034 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8485 = _T_8481 | _T_8484; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8495 = _T_4802 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8498 = _T_8048 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8499 = _T_8495 | _T_8498; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8509 = _T_4806 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8512 = _T_8062 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8513 = _T_8509 | _T_8512; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8523 = _T_4810 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8526 = _T_8076 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8527 = _T_8523 | _T_8526; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8537 = _T_4814 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8540 = _T_8090 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8541 = _T_8537 | _T_8540; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8551 = _T_4818 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8554 = _T_8104 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8555 = _T_8551 | _T_8554; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8565 = _T_4822 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8568 = _T_8118 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8569 = _T_8565 | _T_8568; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8579 = _T_4826 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8582 = _T_8132 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8583 = _T_8579 | _T_8582; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8593 = _T_4830 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8596 = _T_8146 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8597 = _T_8593 | _T_8596; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8607 = _T_4834 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8610 = _T_8160 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8611 = _T_8607 | _T_8610; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8621 = _T_4838 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8624 = _T_8174 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8625 = _T_8621 | _T_8624; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8635 = _T_4842 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8638 = _T_8188 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8639 = _T_8635 | _T_8638; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_8649 = _T_4846 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:58]
  wire  _T_8652 = _T_8202 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 739:123]
  wire  _T_8653 = _T_8649 | _T_8652; // @[el2_ifu_mem_ctl.scala 739:80]
  wire  _T_9454 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 794:63]
  wire  _T_9455 = _T_9454 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 794:85]
  wire [1:0] _T_9457 = _T_9455 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9464; // @[el2_ifu_mem_ctl.scala 799:58]
  reg  _T_9465; // @[el2_ifu_mem_ctl.scala 800:58]
  reg  _T_9466; // @[el2_ifu_mem_ctl.scala 801:59]
  wire  _T_9467 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 802:78]
  wire  _T_9468 = ifu_bus_arvalid_ff & _T_9467; // @[el2_ifu_mem_ctl.scala 802:76]
  wire  _T_9469 = _T_9468 & miss_pending; // @[el2_ifu_mem_ctl.scala 802:98]
  reg  _T_9470; // @[el2_ifu_mem_ctl.scala 802:56]
  reg  _T_9471; // @[el2_ifu_mem_ctl.scala 803:57]
  wire  _T_9474 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 808:71]
  wire  _T_9476 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 808:124]
  wire  _T_9478 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 809:50]
  wire  _T_9480 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 809:103]
  wire [3:0] _T_9483 = {_T_9474,_T_9476,_T_9478,_T_9480}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 811:53]
  reg  _T_9494; // @[Reg.scala 27:20]
  rvclkhdr rvclkhdr ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 319:26]
  assign io_ifu_ic_mb_empty = _T_318 | _T_223; // @[el2_ifu_mem_ctl.scala 318:22]
  assign io_ic_dma_active = _T_12 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 185:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3921; // @[el2_ifu_mem_ctl.scala 686:21]
  assign io_ifu_pmu_ic_miss = _T_9471; // @[el2_ifu_mem_ctl.scala 803:22]
  assign io_ifu_pmu_ic_hit = _T_9470; // @[el2_ifu_mem_ctl.scala 802:21]
  assign io_ifu_pmu_bus_error = _T_9466; // @[el2_ifu_mem_ctl.scala 801:24]
  assign io_ifu_pmu_bus_busy = _T_9465; // @[el2_ifu_mem_ctl.scala 800:23]
  assign io_ifu_pmu_bus_trxn = _T_9464; // @[el2_ifu_mem_ctl.scala 799:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 136:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 135:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 130:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 134:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 132:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 143:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 145:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 138:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 131:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 129:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 127:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 128:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 146:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 141:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 548:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2515; // @[el2_ifu_mem_ctl.scala 549:19]
  assign io_ifu_axi_araddr = _T_2517 & _T_2519; // @[el2_ifu_mem_ctl.scala 550:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 553:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 142:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 551:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 554:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 552:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 144:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 555:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 645:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 643:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 647:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 638:20]
  assign io_iccm_ready = _T_2618 & _T_2612; // @[el2_ifu_mem_ctl.scala 618:17]
  assign io_ic_rw_addr = _T_332 | _T_333; // @[el2_ifu_mem_ctl.scala 328:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 685:15]
  assign io_ic_rd_en = _T_3899 | _T_3904; // @[el2_ifu_mem_ctl.scala 676:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 335:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 335:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 336:23]
  assign io_ifu_ic_debug_rd_data = _T_1203; // @[el2_ifu_mem_ctl.scala 344:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 804:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 806:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 807:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 805:25]
  assign io_ic_debug_way = _T_9483[1:0]; // @[el2_ifu_mem_ctl.scala 808:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9457; // @[el2_ifu_mem_ctl.scala 794:19]
  assign io_iccm_rw_addr = _T_3053[14:0]; // @[el2_ifu_mem_ctl.scala 649:19]
  assign io_iccm_wren = _T_2622 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 620:16]
  assign io_iccm_rden = _T_2626 | _T_2627; // @[el2_ifu_mem_ctl.scala 621:16]
  assign io_iccm_wr_data = _T_3028 ? _T_3029 : _T_3036; // @[el2_ifu_mem_ctl.scala 626:19]
  assign io_iccm_wr_size = _T_2632 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 623:19]
  assign io_ic_hit_f = _T_255 | _T_256; // @[el2_ifu_mem_ctl.scala 280:15]
  assign io_ic_access_fault_f = _T_2402 & _T_309; // @[el2_ifu_mem_ctl.scala 375:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1267; // @[el2_ifu_mem_ctl.scala 376:29]
  assign io_iccm_rd_ecc_single_err = _T_3844 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 662:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 663:29]
  assign io_ic_error_start = _T_1191 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 338:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 184:28]
  assign io_iccm_dma_sb_error = _T_4 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 183:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 380:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 372:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 369:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 370:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9494; // @[el2_ifu_mem_ctl.scala 815:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2407; // @[el2_ifu_mem_ctl.scala 468:27]
  assign io_iccm_correction_state = _T_2435 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 503:28 el2_ifu_mem_ctl.scala 516:32 el2_ifu_mem_ctl.scala 523:32 el2_ifu_mem_ctl.scala 530:32]
  assign rvclkhdr_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_lib.scala 419:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_1_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_1_io_en = _T_1 | io_exu_flush_final; // @[el2_lib.scala 419:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_2_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_2_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_lib.scala 419:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_3_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_3_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_lib.scala 419:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_4_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_4_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_lib.scala 419:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_5_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_5_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_lib.scala 419:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_6_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_6_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_lib.scala 419:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_7_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_7_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_lib.scala 419:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_8_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_8_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_lib.scala 419:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_9_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_9_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_lib.scala 419:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_10_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_10_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_lib.scala 419:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_11_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_11_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_lib.scala 419:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_12_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_12_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_lib.scala 419:16]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_13_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_13_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_lib.scala 419:16]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_14_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_14_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_lib.scala 419:16]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_15_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_15_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_lib.scala 419:16]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_16_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_16_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_lib.scala 419:16]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_17_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_17_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_lib.scala 419:16]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_18_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_18_io_en = tag_valid_clken_0[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_19_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_19_io_en = tag_valid_clken_0[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_20_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_20_io_en = tag_valid_clken_1[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_21_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_21_io_en = tag_valid_clken_1[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_22_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_22_io_en = tag_valid_clken_2[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_23_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_23_io_en = tag_valid_clken_2[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_24_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_24_io_en = tag_valid_clken_3[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_25_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_25_io_en = tag_valid_clken_3[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  perr_state = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  err_stop_state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reset_all_tags = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  imb_ff = _RAND_16[30:0];
  _RAND_17 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_4981 = _RAND_19[6:0];
  _RAND_20 = {1{`RANDOM}};
  _T_4337 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4334 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4331 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4328 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4325 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4322 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4319 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4316 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4313 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4310 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4307 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4304 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4301 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4298 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4295 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4292 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4289 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4286 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4283 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4280 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4277 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4274 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4271 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4268 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4265 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4262 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4259 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4256 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4253 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4250 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4247 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4244 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4241 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4238 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4235 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4232 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4229 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4226 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4223 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4220 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4217 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4214 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4211 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4208 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4205 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4202 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4199 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4196 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4193 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4190 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_4187 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_4184 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_4181 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_4178 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_4175 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_4172 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_4169 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_4166 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_4163 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_4160 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4157 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4154 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4151 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4148 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_4145 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_4142 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_4139 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_4136 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4133 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4130 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4127 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4124 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4121 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4118 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4115 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4112 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_4109 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4106 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_4103 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_4100 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_4097 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_4094 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_4091 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_4088 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_4085 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_4082 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_4079 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_4076 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_4073 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_4070 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_4067 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_4064 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_4061 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_4058 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_4055 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_4052 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_4049 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_4046 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_4043 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_4040 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_4037 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_4034 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_4031 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_4028 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_4025 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_4022 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_4019 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_4016 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_4013 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4010 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4007 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4004 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4001 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_3998 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_3995 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3992 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3989 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3986 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3983 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3980 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3977 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3974 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3971 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3968 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3965 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3962 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3959 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3956 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_148[30:0];
  _RAND_149 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  reset_ic_ff = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  miss_addr = _RAND_155[25:0];
  _RAND_156 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_157[2:0];
  _RAND_158 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_158[0:0];
  _RAND_159 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  _T_1287 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  _T_1289 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  _T_1291 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  _T_1293 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  _T_1295 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  _T_1297 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  _T_1299 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  _T_1301 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  _T_1303 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  _T_1305 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  _T_1307 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  _T_1309 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  _T_1311 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  _T_1313 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  _T_1315 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  _T_1317 = _RAND_175[63:0];
  _RAND_176 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_436[0:0];
  _RAND_437 = {3{`RANDOM}};
  _T_1203 = _RAND_437[70:0];
  _RAND_438 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_438[5:0];
  _RAND_439 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_441[2:0];
  _RAND_442 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_444[0:0];
  _RAND_445 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_445[38:0];
  _RAND_446 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_447[2:0];
  _RAND_448 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_449[0:0];
  _RAND_450 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_450[63:0];
  _RAND_451 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_451[13:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_453[13:0];
  _RAND_454 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_454[6:0];
  _RAND_455 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  way_status_new_ff = _RAND_456[2:0];
  _RAND_457 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  ic_valid_ff = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  _T_9464 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  _T_9465 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  _T_9466 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  _T_9470 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_9471 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_9494 = _RAND_464[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_26) begin
        if (_T_28) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_33) begin
        if (_T_38) begin
          miss_state <= 3'h0;
        end else if (_T_42) begin
          miss_state <= 3'h3;
        end else if (_T_49) begin
          miss_state <= 3'h1;
        end else if (_T_53) begin
          miss_state <= 3'h0;
        end else if (_T_64) begin
          miss_state <= 3'h6;
        end else if (_T_72) begin
          miss_state <= 3'h0;
        end else if (_T_77) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_94) begin
        miss_state <= 3'h0;
      end else if (_T_98) begin
        if (_T_105) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_113) begin
        if (_T_118) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_124) begin
        if (_T_129) begin
          miss_state <= 3'h5;
        end else if (_T_135) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_143) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_34) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_152) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_34) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    reset_ic_ff <= _T_290 & _T_291;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_223) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2558) begin
      if (_T_223) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2554;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1287 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1287 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1289 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1289 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1291 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1291 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1293 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1293 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1295 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1295 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1297 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1297 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1299 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1299 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1301 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1301 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1303 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1303 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1305 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1305 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1307 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1307 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1309 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1309 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1311 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1311 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1313 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1313 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1315 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1315 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1317 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1317 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1203 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1203 <= {{5'd0}, _T_1202};
    end else begin
      _T_1203 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2507) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2582) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2626;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2410) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2412) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2422) begin
        perr_state <= 3'h0;
      end else if (_T_2425) begin
        if (_T_2427) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2431) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2435) begin
        err_stop_state <= 2'h1;
      end else if (_T_2440) begin
        if (_T_2442) begin
          err_stop_state <= 2'h0;
        end else if (_T_2463) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2467) begin
        if (_T_2442) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2484) begin
        if (_T_2488) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1348;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_4981 <= 7'h0;
    end else if (_T_3930) begin
      _T_4981 <= io_ic_debug_addr[9:3];
    end else begin
      _T_4981 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1388;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3865;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3040;
    end else begin
      iccm_dma_rdata <= _T_3041;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3861;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3930) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3933) begin
      way_status_new_ff <= _T_3937;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3933) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_9494 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9494 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_8;
    end
    if (reset) begin
      _T_9464 <= 1'h0;
    end else begin
      _T_9464 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_9465 <= 1'h0;
    end else begin
      _T_9465 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_9466 <= 1'h0;
    end else begin
      _T_9466 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_9470 <= 1'h0;
    end else begin
      _T_9470 <= _T_9469;
    end
    if (reset) begin
      _T_9471 <= 1'h0;
    end else begin
      _T_9471 <= bus_cmd_sent;
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk) begin
    if (reset) begin
      _T_4337 <= 3'h0;
    end else if (_T_3976) begin
      _T_4337 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4334 <= 3'h0;
    end else if (_T_3973) begin
      _T_4334 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4331 <= 3'h0;
    end else if (_T_3970) begin
      _T_4331 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4328 <= 3'h0;
    end else if (_T_3967) begin
      _T_4328 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4325 <= 3'h0;
    end else if (_T_3964) begin
      _T_4325 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4322 <= 3'h0;
    end else if (_T_3961) begin
      _T_4322 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4319 <= 3'h0;
    end else if (_T_3958) begin
      _T_4319 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4316 <= 3'h0;
    end else if (_T_3955) begin
      _T_4316 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk) begin
    if (reset) begin
      _T_4313 <= 3'h0;
    end else if (_T_3976) begin
      _T_4313 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4310 <= 3'h0;
    end else if (_T_3973) begin
      _T_4310 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4307 <= 3'h0;
    end else if (_T_3970) begin
      _T_4307 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4304 <= 3'h0;
    end else if (_T_3967) begin
      _T_4304 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4301 <= 3'h0;
    end else if (_T_3964) begin
      _T_4301 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4298 <= 3'h0;
    end else if (_T_3961) begin
      _T_4298 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4295 <= 3'h0;
    end else if (_T_3958) begin
      _T_4295 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4292 <= 3'h0;
    end else if (_T_3955) begin
      _T_4292 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk) begin
    if (reset) begin
      _T_4289 <= 3'h0;
    end else if (_T_3976) begin
      _T_4289 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4286 <= 3'h0;
    end else if (_T_3973) begin
      _T_4286 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4283 <= 3'h0;
    end else if (_T_3970) begin
      _T_4283 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4280 <= 3'h0;
    end else if (_T_3967) begin
      _T_4280 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4277 <= 3'h0;
    end else if (_T_3964) begin
      _T_4277 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4274 <= 3'h0;
    end else if (_T_3961) begin
      _T_4274 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4271 <= 3'h0;
    end else if (_T_3958) begin
      _T_4271 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4268 <= 3'h0;
    end else if (_T_3955) begin
      _T_4268 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk) begin
    if (reset) begin
      _T_4265 <= 3'h0;
    end else if (_T_3976) begin
      _T_4265 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4262 <= 3'h0;
    end else if (_T_3973) begin
      _T_4262 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4259 <= 3'h0;
    end else if (_T_3970) begin
      _T_4259 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4256 <= 3'h0;
    end else if (_T_3967) begin
      _T_4256 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4253 <= 3'h0;
    end else if (_T_3964) begin
      _T_4253 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4250 <= 3'h0;
    end else if (_T_3961) begin
      _T_4250 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4247 <= 3'h0;
    end else if (_T_3958) begin
      _T_4247 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4244 <= 3'h0;
    end else if (_T_3955) begin
      _T_4244 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk) begin
    if (reset) begin
      _T_4241 <= 3'h0;
    end else if (_T_3976) begin
      _T_4241 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4238 <= 3'h0;
    end else if (_T_3973) begin
      _T_4238 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4235 <= 3'h0;
    end else if (_T_3970) begin
      _T_4235 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4232 <= 3'h0;
    end else if (_T_3967) begin
      _T_4232 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4229 <= 3'h0;
    end else if (_T_3964) begin
      _T_4229 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4226 <= 3'h0;
    end else if (_T_3961) begin
      _T_4226 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4223 <= 3'h0;
    end else if (_T_3958) begin
      _T_4223 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4220 <= 3'h0;
    end else if (_T_3955) begin
      _T_4220 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk) begin
    if (reset) begin
      _T_4217 <= 3'h0;
    end else if (_T_3976) begin
      _T_4217 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4214 <= 3'h0;
    end else if (_T_3973) begin
      _T_4214 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4211 <= 3'h0;
    end else if (_T_3970) begin
      _T_4211 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4208 <= 3'h0;
    end else if (_T_3967) begin
      _T_4208 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4205 <= 3'h0;
    end else if (_T_3964) begin
      _T_4205 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4202 <= 3'h0;
    end else if (_T_3961) begin
      _T_4202 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4199 <= 3'h0;
    end else if (_T_3958) begin
      _T_4199 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4196 <= 3'h0;
    end else if (_T_3955) begin
      _T_4196 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk) begin
    if (reset) begin
      _T_4193 <= 3'h0;
    end else if (_T_3976) begin
      _T_4193 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4190 <= 3'h0;
    end else if (_T_3973) begin
      _T_4190 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4187 <= 3'h0;
    end else if (_T_3970) begin
      _T_4187 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4184 <= 3'h0;
    end else if (_T_3967) begin
      _T_4184 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4181 <= 3'h0;
    end else if (_T_3964) begin
      _T_4181 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4178 <= 3'h0;
    end else if (_T_3961) begin
      _T_4178 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4175 <= 3'h0;
    end else if (_T_3958) begin
      _T_4175 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4172 <= 3'h0;
    end else if (_T_3955) begin
      _T_4172 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk) begin
    if (reset) begin
      _T_4169 <= 3'h0;
    end else if (_T_3976) begin
      _T_4169 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4166 <= 3'h0;
    end else if (_T_3973) begin
      _T_4166 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4163 <= 3'h0;
    end else if (_T_3970) begin
      _T_4163 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4160 <= 3'h0;
    end else if (_T_3967) begin
      _T_4160 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4157 <= 3'h0;
    end else if (_T_3964) begin
      _T_4157 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4154 <= 3'h0;
    end else if (_T_3961) begin
      _T_4154 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4151 <= 3'h0;
    end else if (_T_3958) begin
      _T_4151 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4148 <= 3'h0;
    end else if (_T_3955) begin
      _T_4148 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk) begin
    if (reset) begin
      _T_4145 <= 3'h0;
    end else if (_T_3976) begin
      _T_4145 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4142 <= 3'h0;
    end else if (_T_3973) begin
      _T_4142 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4139 <= 3'h0;
    end else if (_T_3970) begin
      _T_4139 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4136 <= 3'h0;
    end else if (_T_3967) begin
      _T_4136 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4133 <= 3'h0;
    end else if (_T_3964) begin
      _T_4133 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4130 <= 3'h0;
    end else if (_T_3961) begin
      _T_4130 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4127 <= 3'h0;
    end else if (_T_3958) begin
      _T_4127 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4124 <= 3'h0;
    end else if (_T_3955) begin
      _T_4124 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk) begin
    if (reset) begin
      _T_4121 <= 3'h0;
    end else if (_T_3976) begin
      _T_4121 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4118 <= 3'h0;
    end else if (_T_3973) begin
      _T_4118 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4115 <= 3'h0;
    end else if (_T_3970) begin
      _T_4115 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4112 <= 3'h0;
    end else if (_T_3967) begin
      _T_4112 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4109 <= 3'h0;
    end else if (_T_3964) begin
      _T_4109 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4106 <= 3'h0;
    end else if (_T_3961) begin
      _T_4106 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4103 <= 3'h0;
    end else if (_T_3958) begin
      _T_4103 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4100 <= 3'h0;
    end else if (_T_3955) begin
      _T_4100 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk) begin
    if (reset) begin
      _T_4097 <= 3'h0;
    end else if (_T_3976) begin
      _T_4097 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4094 <= 3'h0;
    end else if (_T_3973) begin
      _T_4094 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4091 <= 3'h0;
    end else if (_T_3970) begin
      _T_4091 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4088 <= 3'h0;
    end else if (_T_3967) begin
      _T_4088 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4085 <= 3'h0;
    end else if (_T_3964) begin
      _T_4085 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4082 <= 3'h0;
    end else if (_T_3961) begin
      _T_4082 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4079 <= 3'h0;
    end else if (_T_3958) begin
      _T_4079 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4076 <= 3'h0;
    end else if (_T_3955) begin
      _T_4076 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk) begin
    if (reset) begin
      _T_4073 <= 3'h0;
    end else if (_T_3976) begin
      _T_4073 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4070 <= 3'h0;
    end else if (_T_3973) begin
      _T_4070 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4067 <= 3'h0;
    end else if (_T_3970) begin
      _T_4067 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4064 <= 3'h0;
    end else if (_T_3967) begin
      _T_4064 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4061 <= 3'h0;
    end else if (_T_3964) begin
      _T_4061 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4058 <= 3'h0;
    end else if (_T_3961) begin
      _T_4058 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4055 <= 3'h0;
    end else if (_T_3958) begin
      _T_4055 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4052 <= 3'h0;
    end else if (_T_3955) begin
      _T_4052 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk) begin
    if (reset) begin
      _T_4049 <= 3'h0;
    end else if (_T_3976) begin
      _T_4049 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4046 <= 3'h0;
    end else if (_T_3973) begin
      _T_4046 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4043 <= 3'h0;
    end else if (_T_3970) begin
      _T_4043 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4040 <= 3'h0;
    end else if (_T_3967) begin
      _T_4040 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4037 <= 3'h0;
    end else if (_T_3964) begin
      _T_4037 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4034 <= 3'h0;
    end else if (_T_3961) begin
      _T_4034 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4031 <= 3'h0;
    end else if (_T_3958) begin
      _T_4031 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4028 <= 3'h0;
    end else if (_T_3955) begin
      _T_4028 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk) begin
    if (reset) begin
      _T_4025 <= 3'h0;
    end else if (_T_3976) begin
      _T_4025 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4022 <= 3'h0;
    end else if (_T_3973) begin
      _T_4022 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4019 <= 3'h0;
    end else if (_T_3970) begin
      _T_4019 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4016 <= 3'h0;
    end else if (_T_3967) begin
      _T_4016 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4013 <= 3'h0;
    end else if (_T_3964) begin
      _T_4013 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4010 <= 3'h0;
    end else if (_T_3961) begin
      _T_4010 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4007 <= 3'h0;
    end else if (_T_3958) begin
      _T_4007 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4004 <= 3'h0;
    end else if (_T_3955) begin
      _T_4004 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk) begin
    if (reset) begin
      _T_4001 <= 3'h0;
    end else if (_T_3976) begin
      _T_4001 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3998 <= 3'h0;
    end else if (_T_3973) begin
      _T_3998 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3995 <= 3'h0;
    end else if (_T_3970) begin
      _T_3995 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3992 <= 3'h0;
    end else if (_T_3967) begin
      _T_3992 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3989 <= 3'h0;
    end else if (_T_3964) begin
      _T_3989 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3986 <= 3'h0;
    end else if (_T_3961) begin
      _T_3986 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3983 <= 3'h0;
    end else if (_T_3958) begin
      _T_3983 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3980 <= 3'h0;
    end else if (_T_3955) begin
      _T_3980 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk) begin
    if (reset) begin
      _T_3977 <= 3'h0;
    end else if (_T_3976) begin
      _T_3977 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3974 <= 3'h0;
    end else if (_T_3973) begin
      _T_3974 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3971 <= 3'h0;
    end else if (_T_3970) begin
      _T_3971 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3968 <= 3'h0;
    end else if (_T_3967) begin
      _T_3968 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3965 <= 3'h0;
    end else if (_T_3964) begin
      _T_3965 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3962 <= 3'h0;
    end else if (_T_3961) begin
      _T_3962 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3959 <= 3'h0;
    end else if (_T_3958) begin
      _T_3959 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3956 <= 3'h0;
    end else if (_T_3955) begin
      _T_3956 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5531) begin
      ic_tag_valid_out_1_0 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5545) begin
      ic_tag_valid_out_1_1 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5559) begin
      ic_tag_valid_out_1_2 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5573) begin
      ic_tag_valid_out_1_3 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5587) begin
      ic_tag_valid_out_1_4 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5601) begin
      ic_tag_valid_out_1_5 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5615) begin
      ic_tag_valid_out_1_6 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5629) begin
      ic_tag_valid_out_1_7 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5643) begin
      ic_tag_valid_out_1_8 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5657) begin
      ic_tag_valid_out_1_9 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5671) begin
      ic_tag_valid_out_1_10 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5685) begin
      ic_tag_valid_out_1_11 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5699) begin
      ic_tag_valid_out_1_12 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5713) begin
      ic_tag_valid_out_1_13 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5727) begin
      ic_tag_valid_out_1_14 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5741) begin
      ic_tag_valid_out_1_15 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5755) begin
      ic_tag_valid_out_1_16 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5769) begin
      ic_tag_valid_out_1_17 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5783) begin
      ic_tag_valid_out_1_18 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5797) begin
      ic_tag_valid_out_1_19 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5811) begin
      ic_tag_valid_out_1_20 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5825) begin
      ic_tag_valid_out_1_21 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5839) begin
      ic_tag_valid_out_1_22 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5853) begin
      ic_tag_valid_out_1_23 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5867) begin
      ic_tag_valid_out_1_24 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5881) begin
      ic_tag_valid_out_1_25 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5895) begin
      ic_tag_valid_out_1_26 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5909) begin
      ic_tag_valid_out_1_27 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_5923) begin
      ic_tag_valid_out_1_28 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_5937) begin
      ic_tag_valid_out_1_29 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_5951) begin
      ic_tag_valid_out_1_30 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_5965) begin
      ic_tag_valid_out_1_31 <= _T_5076;
    end
  end
  always @(posedge rvclkhdr_21_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6427) begin
      ic_tag_valid_out_1_32 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6441) begin
      ic_tag_valid_out_1_33 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6455) begin
      ic_tag_valid_out_1_34 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6469) begin
      ic_tag_valid_out_1_35 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6483) begin
      ic_tag_valid_out_1_36 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6497) begin
      ic_tag_valid_out_1_37 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6511) begin
      ic_tag_valid_out_1_38 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6525) begin
      ic_tag_valid_out_1_39 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6539) begin
      ic_tag_valid_out_1_40 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6553) begin
      ic_tag_valid_out_1_41 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6567) begin
      ic_tag_valid_out_1_42 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6581) begin
      ic_tag_valid_out_1_43 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6595) begin
      ic_tag_valid_out_1_44 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6609) begin
      ic_tag_valid_out_1_45 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6623) begin
      ic_tag_valid_out_1_46 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6637) begin
      ic_tag_valid_out_1_47 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6651) begin
      ic_tag_valid_out_1_48 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6665) begin
      ic_tag_valid_out_1_49 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6679) begin
      ic_tag_valid_out_1_50 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6693) begin
      ic_tag_valid_out_1_51 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6707) begin
      ic_tag_valid_out_1_52 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6721) begin
      ic_tag_valid_out_1_53 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6735) begin
      ic_tag_valid_out_1_54 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6749) begin
      ic_tag_valid_out_1_55 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6763) begin
      ic_tag_valid_out_1_56 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6777) begin
      ic_tag_valid_out_1_57 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6791) begin
      ic_tag_valid_out_1_58 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6805) begin
      ic_tag_valid_out_1_59 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6819) begin
      ic_tag_valid_out_1_60 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6833) begin
      ic_tag_valid_out_1_61 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_6847) begin
      ic_tag_valid_out_1_62 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_6861) begin
      ic_tag_valid_out_1_63 <= _T_5076;
    end
  end
  always @(posedge rvclkhdr_23_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7323) begin
      ic_tag_valid_out_1_64 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7337) begin
      ic_tag_valid_out_1_65 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7351) begin
      ic_tag_valid_out_1_66 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7365) begin
      ic_tag_valid_out_1_67 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7379) begin
      ic_tag_valid_out_1_68 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7393) begin
      ic_tag_valid_out_1_69 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7407) begin
      ic_tag_valid_out_1_70 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7421) begin
      ic_tag_valid_out_1_71 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7435) begin
      ic_tag_valid_out_1_72 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7449) begin
      ic_tag_valid_out_1_73 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7463) begin
      ic_tag_valid_out_1_74 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7477) begin
      ic_tag_valid_out_1_75 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7491) begin
      ic_tag_valid_out_1_76 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7505) begin
      ic_tag_valid_out_1_77 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7519) begin
      ic_tag_valid_out_1_78 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7533) begin
      ic_tag_valid_out_1_79 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7547) begin
      ic_tag_valid_out_1_80 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7561) begin
      ic_tag_valid_out_1_81 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7575) begin
      ic_tag_valid_out_1_82 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7589) begin
      ic_tag_valid_out_1_83 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7603) begin
      ic_tag_valid_out_1_84 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7617) begin
      ic_tag_valid_out_1_85 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7631) begin
      ic_tag_valid_out_1_86 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7645) begin
      ic_tag_valid_out_1_87 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7659) begin
      ic_tag_valid_out_1_88 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7673) begin
      ic_tag_valid_out_1_89 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7687) begin
      ic_tag_valid_out_1_90 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7701) begin
      ic_tag_valid_out_1_91 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7715) begin
      ic_tag_valid_out_1_92 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7729) begin
      ic_tag_valid_out_1_93 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7743) begin
      ic_tag_valid_out_1_94 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7757) begin
      ic_tag_valid_out_1_95 <= _T_5076;
    end
  end
  always @(posedge rvclkhdr_25_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8219) begin
      ic_tag_valid_out_1_96 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8233) begin
      ic_tag_valid_out_1_97 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8247) begin
      ic_tag_valid_out_1_98 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8261) begin
      ic_tag_valid_out_1_99 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8275) begin
      ic_tag_valid_out_1_100 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8289) begin
      ic_tag_valid_out_1_101 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8303) begin
      ic_tag_valid_out_1_102 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8317) begin
      ic_tag_valid_out_1_103 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8331) begin
      ic_tag_valid_out_1_104 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8345) begin
      ic_tag_valid_out_1_105 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8359) begin
      ic_tag_valid_out_1_106 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8373) begin
      ic_tag_valid_out_1_107 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8387) begin
      ic_tag_valid_out_1_108 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8401) begin
      ic_tag_valid_out_1_109 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8415) begin
      ic_tag_valid_out_1_110 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8429) begin
      ic_tag_valid_out_1_111 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8443) begin
      ic_tag_valid_out_1_112 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8457) begin
      ic_tag_valid_out_1_113 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8471) begin
      ic_tag_valid_out_1_114 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8485) begin
      ic_tag_valid_out_1_115 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8499) begin
      ic_tag_valid_out_1_116 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8513) begin
      ic_tag_valid_out_1_117 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8527) begin
      ic_tag_valid_out_1_118 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8541) begin
      ic_tag_valid_out_1_119 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8555) begin
      ic_tag_valid_out_1_120 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8569) begin
      ic_tag_valid_out_1_121 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8583) begin
      ic_tag_valid_out_1_122 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8597) begin
      ic_tag_valid_out_1_123 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8611) begin
      ic_tag_valid_out_1_124 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8625) begin
      ic_tag_valid_out_1_125 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8639) begin
      ic_tag_valid_out_1_126 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8653) begin
      ic_tag_valid_out_1_127 <= _T_5076;
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5083) begin
      ic_tag_valid_out_0_0 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5097) begin
      ic_tag_valid_out_0_1 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5111) begin
      ic_tag_valid_out_0_2 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5125) begin
      ic_tag_valid_out_0_3 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5139) begin
      ic_tag_valid_out_0_4 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5153) begin
      ic_tag_valid_out_0_5 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5167) begin
      ic_tag_valid_out_0_6 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5181) begin
      ic_tag_valid_out_0_7 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5195) begin
      ic_tag_valid_out_0_8 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5209) begin
      ic_tag_valid_out_0_9 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5223) begin
      ic_tag_valid_out_0_10 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5237) begin
      ic_tag_valid_out_0_11 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5251) begin
      ic_tag_valid_out_0_12 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5265) begin
      ic_tag_valid_out_0_13 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5279) begin
      ic_tag_valid_out_0_14 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5293) begin
      ic_tag_valid_out_0_15 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5307) begin
      ic_tag_valid_out_0_16 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5321) begin
      ic_tag_valid_out_0_17 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5335) begin
      ic_tag_valid_out_0_18 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5349) begin
      ic_tag_valid_out_0_19 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5363) begin
      ic_tag_valid_out_0_20 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5377) begin
      ic_tag_valid_out_0_21 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5391) begin
      ic_tag_valid_out_0_22 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5405) begin
      ic_tag_valid_out_0_23 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5419) begin
      ic_tag_valid_out_0_24 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5433) begin
      ic_tag_valid_out_0_25 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5447) begin
      ic_tag_valid_out_0_26 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5461) begin
      ic_tag_valid_out_0_27 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5475) begin
      ic_tag_valid_out_0_28 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5489) begin
      ic_tag_valid_out_0_29 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5503) begin
      ic_tag_valid_out_0_30 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5517) begin
      ic_tag_valid_out_0_31 <= _T_5076;
    end
  end
  always @(posedge rvclkhdr_20_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_5979) begin
      ic_tag_valid_out_0_32 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_5993) begin
      ic_tag_valid_out_0_33 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6007) begin
      ic_tag_valid_out_0_34 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6021) begin
      ic_tag_valid_out_0_35 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6035) begin
      ic_tag_valid_out_0_36 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6049) begin
      ic_tag_valid_out_0_37 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6063) begin
      ic_tag_valid_out_0_38 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6077) begin
      ic_tag_valid_out_0_39 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6091) begin
      ic_tag_valid_out_0_40 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6105) begin
      ic_tag_valid_out_0_41 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6119) begin
      ic_tag_valid_out_0_42 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6133) begin
      ic_tag_valid_out_0_43 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6147) begin
      ic_tag_valid_out_0_44 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6161) begin
      ic_tag_valid_out_0_45 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6175) begin
      ic_tag_valid_out_0_46 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6189) begin
      ic_tag_valid_out_0_47 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6203) begin
      ic_tag_valid_out_0_48 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6217) begin
      ic_tag_valid_out_0_49 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6231) begin
      ic_tag_valid_out_0_50 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6245) begin
      ic_tag_valid_out_0_51 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6259) begin
      ic_tag_valid_out_0_52 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6273) begin
      ic_tag_valid_out_0_53 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6287) begin
      ic_tag_valid_out_0_54 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6301) begin
      ic_tag_valid_out_0_55 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6315) begin
      ic_tag_valid_out_0_56 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6329) begin
      ic_tag_valid_out_0_57 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6343) begin
      ic_tag_valid_out_0_58 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6357) begin
      ic_tag_valid_out_0_59 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6371) begin
      ic_tag_valid_out_0_60 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6385) begin
      ic_tag_valid_out_0_61 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6399) begin
      ic_tag_valid_out_0_62 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6413) begin
      ic_tag_valid_out_0_63 <= _T_5076;
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_6875) begin
      ic_tag_valid_out_0_64 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_6889) begin
      ic_tag_valid_out_0_65 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_6903) begin
      ic_tag_valid_out_0_66 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_6917) begin
      ic_tag_valid_out_0_67 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_6931) begin
      ic_tag_valid_out_0_68 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_6945) begin
      ic_tag_valid_out_0_69 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_6959) begin
      ic_tag_valid_out_0_70 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_6973) begin
      ic_tag_valid_out_0_71 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_6987) begin
      ic_tag_valid_out_0_72 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7001) begin
      ic_tag_valid_out_0_73 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7015) begin
      ic_tag_valid_out_0_74 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7029) begin
      ic_tag_valid_out_0_75 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7043) begin
      ic_tag_valid_out_0_76 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7057) begin
      ic_tag_valid_out_0_77 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7071) begin
      ic_tag_valid_out_0_78 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7085) begin
      ic_tag_valid_out_0_79 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7099) begin
      ic_tag_valid_out_0_80 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7113) begin
      ic_tag_valid_out_0_81 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7127) begin
      ic_tag_valid_out_0_82 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7141) begin
      ic_tag_valid_out_0_83 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7155) begin
      ic_tag_valid_out_0_84 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7169) begin
      ic_tag_valid_out_0_85 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7183) begin
      ic_tag_valid_out_0_86 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7197) begin
      ic_tag_valid_out_0_87 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7211) begin
      ic_tag_valid_out_0_88 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7225) begin
      ic_tag_valid_out_0_89 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7239) begin
      ic_tag_valid_out_0_90 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7253) begin
      ic_tag_valid_out_0_91 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7267) begin
      ic_tag_valid_out_0_92 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7281) begin
      ic_tag_valid_out_0_93 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7295) begin
      ic_tag_valid_out_0_94 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7309) begin
      ic_tag_valid_out_0_95 <= _T_5076;
    end
  end
  always @(posedge rvclkhdr_24_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7771) begin
      ic_tag_valid_out_0_96 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_7785) begin
      ic_tag_valid_out_0_97 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_7799) begin
      ic_tag_valid_out_0_98 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_7813) begin
      ic_tag_valid_out_0_99 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_7827) begin
      ic_tag_valid_out_0_100 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_7841) begin
      ic_tag_valid_out_0_101 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_7855) begin
      ic_tag_valid_out_0_102 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_7869) begin
      ic_tag_valid_out_0_103 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_7883) begin
      ic_tag_valid_out_0_104 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_7897) begin
      ic_tag_valid_out_0_105 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_7911) begin
      ic_tag_valid_out_0_106 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_7925) begin
      ic_tag_valid_out_0_107 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_7939) begin
      ic_tag_valid_out_0_108 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_7953) begin
      ic_tag_valid_out_0_109 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_7967) begin
      ic_tag_valid_out_0_110 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_7981) begin
      ic_tag_valid_out_0_111 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_7995) begin
      ic_tag_valid_out_0_112 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8009) begin
      ic_tag_valid_out_0_113 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8023) begin
      ic_tag_valid_out_0_114 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8037) begin
      ic_tag_valid_out_0_115 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8051) begin
      ic_tag_valid_out_0_116 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8065) begin
      ic_tag_valid_out_0_117 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8079) begin
      ic_tag_valid_out_0_118 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8093) begin
      ic_tag_valid_out_0_119 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8107) begin
      ic_tag_valid_out_0_120 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8121) begin
      ic_tag_valid_out_0_121 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8135) begin
      ic_tag_valid_out_0_122 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8149) begin
      ic_tag_valid_out_0_123 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8163) begin
      ic_tag_valid_out_0_124 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8177) begin
      ic_tag_valid_out_0_125 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8191) begin
      ic_tag_valid_out_0_126 <= _T_5076;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8205) begin
      ic_tag_valid_out_0_127 <= _T_5076;
    end
  end
endmodule
