module el2_ifu_compress_ctl(
  input         clock,
  input         reset,
  input  [15:0] io_din,
  output [31:0] io_dout
);
  wire  _T_2 = ~io_din[14]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_4 = ~io_din[13]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_7 = ~io_din[6]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_9 = ~io_din[5]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_11 = io_din[15] & _T_2; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_12 = _T_11 & _T_4; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_13 = _T_12 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_14 = _T_13 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_15 = _T_14 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_16 = _T_15 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_23 = ~io_din[11]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_28 = _T_12 & _T_23; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_29 = _T_28 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_30 = _T_29 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  out_30 = _T_16 | _T_30; // @[el2_ifu_compress_ctl.scala 18:53]
  wire  _T_38 = ~io_din[10]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_40 = ~io_din[9]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_42 = ~io_din[8]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_44 = ~io_din[7]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_50 = ~io_din[4]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_52 = ~io_din[3]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_54 = ~io_din[2]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_56 = _T_2 & io_din[12]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_57 = _T_56 & _T_23; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_58 = _T_57 & _T_38; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_59 = _T_58 & _T_40; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_60 = _T_59 & _T_42; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_61 = _T_60 & _T_44; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_62 = _T_61 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_63 = _T_62 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_64 = _T_63 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_65 = _T_64 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_66 = _T_65 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  out_20 = _T_66 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_79 = _T_28 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_90 = _T_12 & _T_38; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_91 = _T_90 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_92 = _T_79 | _T_91; // @[el2_ifu_compress_ctl.scala 20:46]
  wire  _T_102 = _T_12 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_103 = _T_102 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_104 = _T_92 | _T_103; // @[el2_ifu_compress_ctl.scala 20:80]
  wire  _T_114 = _T_12 & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_115 = _T_114 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  out_14 = _T_104 | _T_115; // @[el2_ifu_compress_ctl.scala 20:113]
  wire  _T_128 = _T_12 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_129 = _T_128 & _T_38; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_130 = _T_129 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_142 = _T_128 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_143 = _T_142 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_144 = _T_130 | _T_143; // @[el2_ifu_compress_ctl.scala 22:50]
  wire  _T_147 = ~io_din[0]; // @[el2_ifu_compress_ctl.scala 22:101]
  wire  _T_148 = io_din[14] & _T_147; // @[el2_ifu_compress_ctl.scala 22:99]
  wire  out_13 = _T_144 | _T_148; // @[el2_ifu_compress_ctl.scala 22:86]
  wire  _T_161 = _T_102 & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_162 = _T_161 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_175 = _T_162 | _T_79; // @[el2_ifu_compress_ctl.scala 23:47]
  wire  _T_188 = _T_175 | _T_91; // @[el2_ifu_compress_ctl.scala 23:81]
  wire  _T_190 = ~io_din[15]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_194 = _T_190 & _T_2; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_195 = _T_194 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_196 = _T_188 | _T_195; // @[el2_ifu_compress_ctl.scala 23:115]
  wire  _T_200 = io_din[15] & io_din[14]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_201 = _T_200 & io_din[13]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  out_12 = _T_196 | _T_201; // @[el2_ifu_compress_ctl.scala 24:26]
  wire  _T_217 = _T_11 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_218 = _T_217 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_219 = _T_218 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_220 = _T_219 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_221 = _T_220 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_224 = _T_221 & _T_147; // @[el2_ifu_compress_ctl.scala 25:53]
  wire  _T_228 = _T_2 & io_din[13]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_229 = _T_224 | _T_228; // @[el2_ifu_compress_ctl.scala 25:67]
  wire  _T_234 = _T_200 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  out_6 = _T_229 | _T_234; // @[el2_ifu_compress_ctl.scala 25:88]
  wire  _T_239 = io_din[15] & _T_147; // @[el2_ifu_compress_ctl.scala 26:24]
  wire  _T_243 = io_din[15] & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_244 = _T_243 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_245 = _T_239 | _T_244; // @[el2_ifu_compress_ctl.scala 26:39]
  wire  _T_249 = io_din[13] & _T_42; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_250 = _T_245 | _T_249; // @[el2_ifu_compress_ctl.scala 26:63]
  wire  _T_253 = io_din[13] & io_din[7]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_254 = _T_250 | _T_253; // @[el2_ifu_compress_ctl.scala 26:83]
  wire  _T_257 = io_din[13] & io_din[9]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_258 = _T_254 | _T_257; // @[el2_ifu_compress_ctl.scala 26:102]
  wire  _T_261 = io_din[13] & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_262 = _T_258 | _T_261; // @[el2_ifu_compress_ctl.scala 27:22]
  wire  _T_265 = io_din[13] & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_266 = _T_262 | _T_265; // @[el2_ifu_compress_ctl.scala 27:42]
  wire  _T_271 = _T_266 | _T_228; // @[el2_ifu_compress_ctl.scala 27:62]
  wire  out_5 = _T_271 | _T_200; // @[el2_ifu_compress_ctl.scala 27:83]
  wire  _T_288 = _T_2 & _T_23; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_289 = _T_288 & _T_38; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_290 = _T_289 & _T_40; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_291 = _T_290 & _T_42; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_292 = _T_291 & _T_44; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_295 = _T_292 & _T_147; // @[el2_ifu_compress_ctl.scala 28:50]
  wire  _T_303 = _T_194 & _T_147; // @[el2_ifu_compress_ctl.scala 28:87]
  wire  _T_304 = _T_295 | _T_303; // @[el2_ifu_compress_ctl.scala 28:65]
  wire  _T_308 = _T_2 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_311 = _T_308 & _T_147; // @[el2_ifu_compress_ctl.scala 29:23]
  wire  _T_312 = _T_304 | _T_311; // @[el2_ifu_compress_ctl.scala 28:102]
  wire  _T_317 = _T_190 & io_din[14]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_318 = _T_317 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_319 = _T_312 | _T_318; // @[el2_ifu_compress_ctl.scala 29:38]
  wire  _T_323 = _T_2 & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_326 = _T_323 & _T_147; // @[el2_ifu_compress_ctl.scala 29:82]
  wire  _T_327 = _T_319 | _T_326; // @[el2_ifu_compress_ctl.scala 29:62]
  wire  _T_331 = _T_2 & io_din[4]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_334 = _T_331 & _T_147; // @[el2_ifu_compress_ctl.scala 30:23]
  wire  _T_335 = _T_327 | _T_334; // @[el2_ifu_compress_ctl.scala 29:97]
  wire  _T_339 = _T_2 & io_din[3]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_342 = _T_339 & _T_147; // @[el2_ifu_compress_ctl.scala 30:58]
  wire  _T_343 = _T_335 | _T_342; // @[el2_ifu_compress_ctl.scala 30:38]
  wire  _T_347 = _T_2 & io_din[2]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_350 = _T_347 & _T_147; // @[el2_ifu_compress_ctl.scala 30:93]
  wire  _T_351 = _T_343 | _T_350; // @[el2_ifu_compress_ctl.scala 30:73]
  wire  _T_357 = _T_2 & _T_4; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_358 = _T_357 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  out_4 = _T_351 | _T_358; // @[el2_ifu_compress_ctl.scala 30:108]
  wire  _T_380 = _T_56 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_381 = _T_380 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_382 = _T_381 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_383 = _T_382 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_384 = _T_383 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_385 = _T_384 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_386 = _T_385 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_403 = _T_56 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_404 = _T_403 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_405 = _T_404 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_406 = _T_405 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_407 = _T_406 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_408 = _T_407 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_409 = _T_408 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_410 = _T_386 | _T_409; // @[el2_ifu_compress_ctl.scala 33:59]
  wire  _T_427 = _T_56 & io_din[9]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_428 = _T_427 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_429 = _T_428 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_430 = _T_429 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_431 = _T_430 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_432 = _T_431 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_433 = _T_432 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_434 = _T_410 | _T_433; // @[el2_ifu_compress_ctl.scala 33:107]
  wire  _T_450 = _T_56 & io_din[8]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_451 = _T_450 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_452 = _T_451 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_453 = _T_452 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_454 = _T_453 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_455 = _T_454 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_456 = _T_455 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_457 = _T_434 | _T_456; // @[el2_ifu_compress_ctl.scala 34:48]
  wire  _T_474 = _T_56 & io_din[7]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_475 = _T_474 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_476 = _T_475 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_477 = _T_476 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_478 = _T_477 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_479 = _T_478 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_480 = _T_479 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_481 = _T_457 | _T_480; // @[el2_ifu_compress_ctl.scala 34:86]
  wire  _T_486 = ~io_din[12]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_498 = _T_11 & _T_486; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_499 = _T_498 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_500 = _T_499 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_501 = _T_500 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_502 = _T_501 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_503 = _T_502 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_506 = _T_503 & _T_147; // @[el2_ifu_compress_ctl.scala 35:42]
  wire  _T_507 = _T_481 | _T_506; // @[el2_ifu_compress_ctl.scala 34:125]
  wire  _T_513 = _T_190 & io_din[13]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_514 = _T_513 & _T_42; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_515 = _T_507 | _T_514; // @[el2_ifu_compress_ctl.scala 35:57]
  wire  _T_521 = _T_513 & io_din[7]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_522 = _T_515 | _T_521; // @[el2_ifu_compress_ctl.scala 35:80]
  wire  _T_528 = _T_513 & io_din[9]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_529 = _T_522 | _T_528; // @[el2_ifu_compress_ctl.scala 35:102]
  wire  _T_535 = _T_513 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_536 = _T_529 | _T_535; // @[el2_ifu_compress_ctl.scala 35:124]
  wire  _T_542 = _T_513 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_543 = _T_536 | _T_542; // @[el2_ifu_compress_ctl.scala 36:24]
  wire  out_2 = _T_543 | _T_228; // @[el2_ifu_compress_ctl.scala 36:47]
  wire [4:0] rs2d = io_din[6:2]; // @[el2_ifu_compress_ctl.scala 44:20]
  wire [4:0] rdd = io_din[11:7]; // @[el2_ifu_compress_ctl.scala 45:19]
  wire [4:0] rdpd = {2'h1,io_din[9:7]}; // @[Cat.scala 29:58]
  wire [4:0] rs2pd = {2'h1,io_din[4:2]}; // @[Cat.scala 29:58]
  wire  _T_556 = _T_308 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_563 = _T_317 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_564 = _T_563 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_565 = _T_556 | _T_564; // @[el2_ifu_compress_ctl.scala 49:33]
  wire  _T_571 = _T_323 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_572 = _T_565 | _T_571; // @[el2_ifu_compress_ctl.scala 49:58]
  wire  _T_579 = _T_317 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_580 = _T_579 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_581 = _T_572 | _T_580; // @[el2_ifu_compress_ctl.scala 49:79]
  wire  _T_587 = _T_331 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_588 = _T_581 | _T_587; // @[el2_ifu_compress_ctl.scala 49:104]
  wire  _T_595 = _T_317 & io_din[9]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_596 = _T_595 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_597 = _T_588 | _T_596; // @[el2_ifu_compress_ctl.scala 50:24]
  wire  _T_603 = _T_339 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_604 = _T_597 | _T_603; // @[el2_ifu_compress_ctl.scala 50:48]
  wire  _T_612 = _T_317 & _T_42; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_613 = _T_612 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_614 = _T_604 | _T_613; // @[el2_ifu_compress_ctl.scala 50:69]
  wire  _T_620 = _T_347 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_621 = _T_614 | _T_620; // @[el2_ifu_compress_ctl.scala 50:94]
  wire  _T_628 = _T_317 & io_din[7]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_629 = _T_628 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_630 = _T_621 | _T_629; // @[el2_ifu_compress_ctl.scala 51:22]
  wire  _T_634 = _T_190 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_635 = _T_630 | _T_634; // @[el2_ifu_compress_ctl.scala 51:46]
  wire  _T_641 = _T_190 & _T_4; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_642 = _T_641 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  rdrd = _T_635 | _T_642; // @[el2_ifu_compress_ctl.scala 51:65]
  wire  _T_650 = _T_380 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_658 = _T_403 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_659 = _T_650 | _T_658; // @[el2_ifu_compress_ctl.scala 53:38]
  wire  _T_667 = _T_427 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_668 = _T_659 | _T_667; // @[el2_ifu_compress_ctl.scala 53:63]
  wire  _T_676 = _T_450 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_677 = _T_668 | _T_676; // @[el2_ifu_compress_ctl.scala 53:87]
  wire  _T_685 = _T_474 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_686 = _T_677 | _T_685; // @[el2_ifu_compress_ctl.scala 53:111]
  wire  _T_702 = _T_2 & _T_486; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_703 = _T_702 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_704 = _T_703 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_705 = _T_704 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_706 = _T_705 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_707 = _T_706 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_708 = _T_707 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_709 = _T_686 | _T_708; // @[el2_ifu_compress_ctl.scala 54:27]
  wire  _T_716 = _T_56 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_717 = _T_716 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_718 = _T_709 | _T_717; // @[el2_ifu_compress_ctl.scala 54:65]
  wire  _T_725 = _T_56 & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_726 = _T_725 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_727 = _T_718 | _T_726; // @[el2_ifu_compress_ctl.scala 54:89]
  wire  _T_734 = _T_56 & io_din[4]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_735 = _T_734 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_736 = _T_727 | _T_735; // @[el2_ifu_compress_ctl.scala 54:113]
  wire  _T_743 = _T_56 & io_din[3]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_744 = _T_743 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_745 = _T_736 | _T_744; // @[el2_ifu_compress_ctl.scala 55:27]
  wire  _T_752 = _T_56 & io_din[2]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_753 = _T_752 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_754 = _T_745 | _T_753; // @[el2_ifu_compress_ctl.scala 55:51]
  wire  _T_763 = _T_194 & _T_4; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_764 = _T_763 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  rdrs1 = _T_754 | _T_764; // @[el2_ifu_compress_ctl.scala 55:75]
  wire  _T_768 = io_din[15] & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_769 = _T_768 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_773 = io_din[15] & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_774 = _T_773 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_775 = _T_769 | _T_774; // @[el2_ifu_compress_ctl.scala 57:34]
  wire  _T_779 = io_din[15] & io_din[4]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_780 = _T_779 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_781 = _T_775 | _T_780; // @[el2_ifu_compress_ctl.scala 57:54]
  wire  _T_785 = io_din[15] & io_din[3]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_786 = _T_785 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_787 = _T_781 | _T_786; // @[el2_ifu_compress_ctl.scala 57:74]
  wire  _T_791 = io_din[15] & io_din[2]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_792 = _T_791 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_793 = _T_787 | _T_792; // @[el2_ifu_compress_ctl.scala 57:94]
  wire  _T_798 = _T_200 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  rs2rs2 = _T_793 | _T_798; // @[el2_ifu_compress_ctl.scala 57:114]
  wire  rdprd = _T_12 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_811 = io_din[15] & _T_4; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_812 = _T_811 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_818 = _T_812 | _T_234; // @[el2_ifu_compress_ctl.scala 61:36]
  wire  _T_821 = ~io_din[1]; // @[el2_ifu_compress_ctl.scala 15:83]
  wire  _T_822 = io_din[14] & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_825 = _T_822 & _T_147; // @[el2_ifu_compress_ctl.scala 61:76]
  wire  rdprs1 = _T_818 | _T_825; // @[el2_ifu_compress_ctl.scala 61:57]
  wire  _T_837 = _T_128 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_838 = _T_837 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_842 = io_din[15] & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_845 = _T_842 & _T_147; // @[el2_ifu_compress_ctl.scala 63:66]
  wire  rs2prs2 = _T_838 | _T_845; // @[el2_ifu_compress_ctl.scala 63:47]
  wire  _T_850 = _T_190 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  rs2prd = _T_850 & _T_147; // @[el2_ifu_compress_ctl.scala 64:33]
  wire  _T_857 = _T_2 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  uimm9_2 = _T_857 & _T_147; // @[el2_ifu_compress_ctl.scala 65:34]
  wire  _T_866 = _T_317 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  ulwimm6_2 = _T_866 & _T_147; // @[el2_ifu_compress_ctl.scala 66:39]
  wire  ulwspimm7_2 = _T_317 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_888 = _T_317 & io_din[13]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_889 = _T_888 & _T_23; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_890 = _T_889 & _T_38; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_891 = _T_890 & _T_40; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_892 = _T_891 & io_din[8]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  rdeq2 = _T_892 & _T_44; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_981 = _T_450 & _T_7; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_982 = _T_981 & _T_9; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_983 = _T_982 & _T_50; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_984 = _T_983 & _T_52; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_985 = _T_984 & _T_54; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_986 = _T_985 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_987 = _T_434 | _T_986; // @[el2_ifu_compress_ctl.scala 70:42]
  wire  _T_1011 = _T_987 | _T_480; // @[el2_ifu_compress_ctl.scala 70:81]
  wire  _T_1018 = _T_194 & io_din[13]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  rdeq1 = _T_1011 | _T_1018; // @[el2_ifu_compress_ctl.scala 71:42]
  wire  _T_1041 = io_din[14] & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1042 = rdeq2 | _T_1041; // @[el2_ifu_compress_ctl.scala 72:53]
  wire  rs1eq2 = _T_1042 | uimm9_2; // @[el2_ifu_compress_ctl.scala 72:71]
  wire  _T_1083 = _T_357 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1084 = _T_1083 & _T_38; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1085 = _T_1084 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  simm5_0 = _T_1085 | _T_642; // @[el2_ifu_compress_ctl.scala 75:45]
  wire  _T_1103 = _T_888 & io_din[7]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1112 = _T_888 & _T_42; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1113 = _T_1103 | _T_1112; // @[el2_ifu_compress_ctl.scala 77:44]
  wire  _T_1121 = _T_888 & io_din[9]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1122 = _T_1113 | _T_1121; // @[el2_ifu_compress_ctl.scala 77:70]
  wire  _T_1130 = _T_888 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1131 = _T_1122 | _T_1130; // @[el2_ifu_compress_ctl.scala 77:95]
  wire  _T_1139 = _T_888 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  sluimm17_12 = _T_1131 | _T_1139; // @[el2_ifu_compress_ctl.scala 78:29]
  wire  uimm5_0 = _T_79 | _T_195; // @[el2_ifu_compress_ctl.scala 79:45]
  wire [4:0] _T_1185 = rdrd ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1186 = rdprd ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1187 = rs2prd ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1188 = rdeq1 ? 5'h1 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1189 = rdeq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1190 = _T_1185 | _T_1186; // @[Mux.scala 27:72]
  wire [4:0] _T_1191 = _T_1190 | _T_1187; // @[Mux.scala 27:72]
  wire [4:0] _T_1192 = _T_1191 | _T_1188; // @[Mux.scala 27:72]
  wire [4:0] l1_11 = _T_1192 | _T_1189; // @[Mux.scala 27:72]
  wire [4:0] _T_1204 = rdrs1 ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1205 = rdprs1 ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1206 = rs1eq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1207 = _T_1204 | _T_1205; // @[Mux.scala 27:72]
  wire [4:0] l1_19 = _T_1207 | _T_1206; // @[Mux.scala 27:72]
  wire [4:0] _T_1214 = {out_20,1'h0,1'h0,2'h0}; // @[el2_ifu_compress_ctl.scala 90:64]
  wire [4:0] _T_1217 = rs2rs2 ? rs2d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1218 = rs2prs2 ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1219 = _T_1217 | _T_1218; // @[Mux.scala 27:72]
  wire [4:0] l1_24 = _T_1214 | _T_1219; // @[el2_ifu_compress_ctl.scala 90:71]
  wire [14:0] _T_1228 = {out_14,out_13,out_12,l1_11,2'h3,out_2,_T_228,out_4,out_5,out_6}; // @[Cat.scala 29:58]
  wire [31:0] l1 = {4'h0,1'h0,out_30,1'h0,l1_24,l1_19,_T_1228}; // @[Cat.scala 29:58]
  wire [5:0] simm5d = {io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [5:0] simm9d = {io_din[12],io_din[4:3],io_din[5],io_din[2],io_din[6]}; // @[Cat.scala 29:58]
  wire [8:0] sjald_12 = io_din[12] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [19:0] sjald = {sjald_12,io_din[12],io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:4],io_din[3]}; // @[Cat.scala 29:58]
  wire [14:0] _T_1277 = io_din[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [19:0] sluimmd = {_T_1277,rs2d}; // @[Cat.scala 29:58]
  wire [6:0] _T_1283 = simm5d[5] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_1285 = {_T_1283,simm5d[4:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1288 = {2'h0,io_din[10:7],io_din[12:11],io_din[5],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [2:0] _T_1292 = simm9d[5] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_1295 = {_T_1292,simm9d[4:0],4'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1298 = {5'h0,io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1301 = {4'h0,io_din[3:2],io_din[12],io_din[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1303 = {6'h0,io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1308 = {sjald[19],sjald[9:0],sjald[10]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1310 = simm5_0 ? _T_1285 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1311 = uimm9_2 ? _T_1288 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1312 = rdeq2 ? _T_1295 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1313 = ulwimm6_2 ? _T_1298 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1314 = ulwspimm7_2 ? _T_1301 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1315 = uimm5_0 ? _T_1303 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1316 = _T_228 ? _T_1308 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1317 = sluimm17_12 ? sluimmd[19:8] : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1318 = _T_1310 | _T_1311; // @[Mux.scala 27:72]
  wire [11:0] _T_1319 = _T_1318 | _T_1312; // @[Mux.scala 27:72]
  wire [11:0] _T_1320 = _T_1319 | _T_1313; // @[Mux.scala 27:72]
  wire [11:0] _T_1321 = _T_1320 | _T_1314; // @[Mux.scala 27:72]
  wire [11:0] _T_1322 = _T_1321 | _T_1315; // @[Mux.scala 27:72]
  wire [11:0] _T_1323 = _T_1322 | _T_1316; // @[Mux.scala 27:72]
  wire [11:0] _T_1324 = _T_1323 | _T_1317; // @[Mux.scala 27:72]
  wire [11:0] l2_31 = l1[31:20] | _T_1324; // @[el2_ifu_compress_ctl.scala 106:25]
  wire [8:0] _T_1331 = _T_228 ? sjald[19:11] : 9'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1332 = sluimm17_12 ? sluimmd[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [8:0] _GEN_0 = {{1'd0}, _T_1332}; // @[Mux.scala 27:72]
  wire [8:0] _T_1333 = _T_1331 | _GEN_0; // @[Mux.scala 27:72]
  wire [8:0] _GEN_1 = {{1'd0}, l1[19:12]}; // @[el2_ifu_compress_ctl.scala 116:25]
  wire [8:0] l2_19 = _GEN_1 | _T_1333; // @[el2_ifu_compress_ctl.scala 116:25]
  wire [32:0] l2 = {l2_31,l2_19,l1[11:0]}; // @[Cat.scala 29:58]
  wire [8:0] sbr8d = {io_din[12],io_din[6],io_din[5],io_din[2],io_din[11],io_din[10],io_din[4],io_din[3],1'h0}; // @[Cat.scala 29:58]
  wire [6:0] uswimm6d = {io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [7:0] uswspimm7d = {io_din[8:7],io_din[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_1364 = sbr8d[8] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _T_1366 = {_T_1364,sbr8d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1369 = {5'h0,uswimm6d[6:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1372 = {4'h0,uswspimm7d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1373 = _T_234 ? _T_1366 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1374 = _T_845 ? _T_1369 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1375 = _T_798 ? _T_1372 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1376 = _T_1373 | _T_1374; // @[Mux.scala 27:72]
  wire [6:0] _T_1377 = _T_1376 | _T_1375; // @[Mux.scala 27:72]
  wire [6:0] l3_31 = l2[31:25] | _T_1377; // @[el2_ifu_compress_ctl.scala 122:25]
  wire [12:0] l3_24 = l2[24:12]; // @[el2_ifu_compress_ctl.scala 125:17]
  wire [4:0] _T_1383 = {sbr8d[4:1],sbr8d[8]}; // @[Cat.scala 29:58]
  wire [4:0] _T_1388 = _T_234 ? _T_1383 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1389 = _T_845 ? uswimm6d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1390 = _T_798 ? uswspimm7d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1391 = _T_1388 | _T_1389; // @[Mux.scala 27:72]
  wire [4:0] _T_1392 = _T_1391 | _T_1390; // @[Mux.scala 27:72]
  wire [4:0] l3_11 = l2[11:7] | _T_1392; // @[el2_ifu_compress_ctl.scala 126:24]
  wire [31:0] l3 = {l3_31,l3_24,l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire  _T_1403 = _T_4 & _T_486; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1404 = _T_1403 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1405 = _T_1404 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1408 = _T_1405 & _T_147; // @[el2_ifu_compress_ctl.scala 131:39]
  wire  _T_1416 = _T_1403 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1417 = _T_1416 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1420 = _T_1417 & _T_147; // @[el2_ifu_compress_ctl.scala 131:79]
  wire  _T_1421 = _T_1408 | _T_1420; // @[el2_ifu_compress_ctl.scala 131:54]
  wire  _T_1430 = _T_641 & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1431 = _T_1430 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1432 = _T_1421 | _T_1431; // @[el2_ifu_compress_ctl.scala 131:94]
  wire  _T_1440 = _T_1403 & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1441 = _T_1440 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1444 = _T_1441 & _T_147; // @[el2_ifu_compress_ctl.scala 132:55]
  wire  _T_1445 = _T_1432 | _T_1444; // @[el2_ifu_compress_ctl.scala 132:30]
  wire  _T_1453 = _T_1403 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1454 = _T_1453 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1457 = _T_1454 & _T_147; // @[el2_ifu_compress_ctl.scala 132:96]
  wire  _T_1458 = _T_1445 | _T_1457; // @[el2_ifu_compress_ctl.scala 132:70]
  wire  _T_1467 = _T_641 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1468 = _T_1467 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1469 = _T_1458 | _T_1468; // @[el2_ifu_compress_ctl.scala 132:111]
  wire  _T_1476 = io_din[15] & _T_486; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1477 = _T_1476 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1478 = _T_1477 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1479 = _T_1469 | _T_1478; // @[el2_ifu_compress_ctl.scala 133:29]
  wire  _T_1487 = _T_1403 & io_din[9]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1488 = _T_1487 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1491 = _T_1488 & _T_147; // @[el2_ifu_compress_ctl.scala 133:79]
  wire  _T_1492 = _T_1479 | _T_1491; // @[el2_ifu_compress_ctl.scala 133:54]
  wire  _T_1499 = _T_486 & io_din[6]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1500 = _T_1499 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1501 = _T_1500 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1502 = _T_1492 | _T_1501; // @[el2_ifu_compress_ctl.scala 133:94]
  wire  _T_1511 = _T_641 & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1512 = _T_1511 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1513 = _T_1502 | _T_1512; // @[el2_ifu_compress_ctl.scala 133:118]
  wire  _T_1521 = _T_1403 & io_din[8]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1522 = _T_1521 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1525 = _T_1522 & _T_147; // @[el2_ifu_compress_ctl.scala 134:28]
  wire  _T_1526 = _T_1513 | _T_1525; // @[el2_ifu_compress_ctl.scala 133:144]
  wire  _T_1533 = _T_486 & io_din[5]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1534 = _T_1533 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1535 = _T_1534 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1536 = _T_1526 | _T_1535; // @[el2_ifu_compress_ctl.scala 134:43]
  wire  _T_1545 = _T_641 & io_din[10]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1546 = _T_1545 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1547 = _T_1536 | _T_1546; // @[el2_ifu_compress_ctl.scala 134:67]
  wire  _T_1555 = _T_1403 & io_din[7]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1556 = _T_1555 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1559 = _T_1556 & _T_147; // @[el2_ifu_compress_ctl.scala 135:28]
  wire  _T_1560 = _T_1547 | _T_1559; // @[el2_ifu_compress_ctl.scala 134:94]
  wire  _T_1568 = io_din[12] & io_din[11]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1569 = _T_1568 & _T_38; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1570 = _T_1569 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1571 = _T_1570 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1572 = _T_1560 | _T_1571; // @[el2_ifu_compress_ctl.scala 135:43]
  wire  _T_1581 = _T_641 & io_din[9]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1582 = _T_1581 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1583 = _T_1572 | _T_1582; // @[el2_ifu_compress_ctl.scala 135:71]
  wire  _T_1591 = _T_1403 & io_din[4]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1592 = _T_1591 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1595 = _T_1592 & _T_147; // @[el2_ifu_compress_ctl.scala 136:28]
  wire  _T_1596 = _T_1583 | _T_1595; // @[el2_ifu_compress_ctl.scala 135:97]
  wire  _T_1602 = io_din[13] & io_din[12]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1603 = _T_1602 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1604 = _T_1603 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1605 = _T_1596 | _T_1604; // @[el2_ifu_compress_ctl.scala 136:43]
  wire  _T_1614 = _T_641 & io_din[8]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1615 = _T_1614 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1616 = _T_1605 | _T_1615; // @[el2_ifu_compress_ctl.scala 136:67]
  wire  _T_1624 = _T_1403 & io_din[3]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1625 = _T_1624 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1628 = _T_1625 & _T_147; // @[el2_ifu_compress_ctl.scala 137:28]
  wire  _T_1629 = _T_1616 | _T_1628; // @[el2_ifu_compress_ctl.scala 136:93]
  wire  _T_1635 = io_din[13] & io_din[4]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1636 = _T_1635 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1637 = _T_1636 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1638 = _T_1629 | _T_1637; // @[el2_ifu_compress_ctl.scala 137:43]
  wire  _T_1646 = _T_1403 & io_din[2]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1647 = _T_1646 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1650 = _T_1647 & _T_147; // @[el2_ifu_compress_ctl.scala 137:91]
  wire  _T_1651 = _T_1638 | _T_1650; // @[el2_ifu_compress_ctl.scala 137:66]
  wire  _T_1660 = _T_641 & io_din[7]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1661 = _T_1660 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1662 = _T_1651 | _T_1661; // @[el2_ifu_compress_ctl.scala 137:106]
  wire  _T_1668 = io_din[13] & io_din[3]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1669 = _T_1668 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1670 = _T_1669 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1671 = _T_1662 | _T_1670; // @[el2_ifu_compress_ctl.scala 138:29]
  wire  _T_1677 = io_din[13] & io_din[2]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1678 = _T_1677 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1679 = _T_1678 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1680 = _T_1671 | _T_1679; // @[el2_ifu_compress_ctl.scala 138:52]
  wire  _T_1686 = io_din[14] & _T_4; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1687 = _T_1686 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1688 = _T_1680 | _T_1687; // @[el2_ifu_compress_ctl.scala 138:75]
  wire  _T_1697 = _T_702 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1698 = _T_1697 & io_din[0]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1699 = _T_1688 | _T_1698; // @[el2_ifu_compress_ctl.scala 138:98]
  wire  _T_1706 = _T_811 & io_din[12]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1707 = _T_1706 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1710 = _T_1707 & _T_147; // @[el2_ifu_compress_ctl.scala 139:54]
  wire  _T_1711 = _T_1699 | _T_1710; // @[el2_ifu_compress_ctl.scala 139:29]
  wire  _T_1720 = _T_641 & _T_486; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1721 = _T_1720 & io_din[1]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1724 = _T_1721 & _T_147; // @[el2_ifu_compress_ctl.scala 139:96]
  wire  _T_1725 = _T_1711 | _T_1724; // @[el2_ifu_compress_ctl.scala 139:69]
  wire  _T_1734 = _T_641 & io_din[12]; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1735 = _T_1734 & _T_821; // @[el2_ifu_compress_ctl.scala 15:110]
  wire  _T_1736 = _T_1725 | _T_1735; // @[el2_ifu_compress_ctl.scala 139:111]
  wire  _T_1743 = _T_1686 & _T_147; // @[el2_ifu_compress_ctl.scala 140:50]
  wire  legal = _T_1736 | _T_1743; // @[el2_ifu_compress_ctl.scala 140:30]
  wire [31:0] _T_1745 = legal ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  assign io_dout = l3 & _T_1745; // @[el2_ifu_compress_ctl.scala 142:10]
endmodule
