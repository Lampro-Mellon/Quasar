module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 185:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 321:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 322:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 322:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 254:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 548:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 550:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 187:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 309:34]
  wire [4:0] _GEN_464 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 665:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_464 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 665:53]
  wire [1:0] _GEN_465 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 668:91]
  wire [1:0] _T_3121 = ic_fetch_val_shift_right[3:2] & _GEN_465; // @[el2_ifu_mem_ctl.scala 668:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 323:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 276:46]
  wire [1:0] _GEN_466 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 668:113]
  wire [1:0] _T_3122 = _T_3121 & _GEN_466; // @[el2_ifu_mem_ctl.scala 668:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 654:59]
  wire [1:0] _GEN_467 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 668:130]
  wire [1:0] _T_3123 = _T_3122 | _GEN_467; // @[el2_ifu_mem_ctl.scala 668:130]
  wire  _T_3124 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 668:154]
  wire [1:0] _GEN_468 = {{1'd0}, _T_3124}; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [1:0] _T_3125 = _T_3123 & _GEN_468; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [1:0] _T_3114 = ic_fetch_val_shift_right[1:0] & _GEN_465; // @[el2_ifu_mem_ctl.scala 668:91]
  wire [1:0] _T_3115 = _T_3114 & _GEN_466; // @[el2_ifu_mem_ctl.scala 668:113]
  wire [1:0] _T_3116 = _T_3115 | _GEN_467; // @[el2_ifu_mem_ctl.scala 668:130]
  wire [1:0] _T_3118 = _T_3116 & _GEN_468; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3125,_T_3118}; // @[Cat.scala 29:58]
  wire  _T_3225 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3226 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3227 = _T_3225 ^ _T_3226; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3235 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3236 = ^_T_3235; // @[el2_lib.scala 301:83]
  wire  _T_3237 = io_iccm_rd_data_ecc[37] ^ _T_3236; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3244 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3252 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3244}; // @[el2_lib.scala 301:103]
  wire  _T_3253 = ^_T_3252; // @[el2_lib.scala 301:110]
  wire  _T_3254 = io_iccm_rd_data_ecc[36] ^ _T_3253; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3261 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3269 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3261}; // @[el2_lib.scala 301:130]
  wire  _T_3270 = ^_T_3269; // @[el2_lib.scala 301:137]
  wire  _T_3271 = io_iccm_rd_data_ecc[35] ^ _T_3270; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3280 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3289 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3280}; // @[el2_lib.scala 301:157]
  wire  _T_3290 = ^_T_3289; // @[el2_lib.scala 301:164]
  wire  _T_3291 = io_iccm_rd_data_ecc[34] ^ _T_3290; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3300 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3309 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3300}; // @[el2_lib.scala 301:184]
  wire  _T_3310 = ^_T_3309; // @[el2_lib.scala 301:191]
  wire  _T_3311 = io_iccm_rd_data_ecc[33] ^ _T_3310; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3320 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3329 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3320}; // @[el2_lib.scala 301:211]
  wire  _T_3330 = ^_T_3329; // @[el2_lib.scala 301:218]
  wire  _T_3331 = io_iccm_rd_data_ecc[32] ^ _T_3330; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3337 = {_T_3227,_T_3237,_T_3254,_T_3271,_T_3291,_T_3311,_T_3331}; // @[Cat.scala 29:58]
  wire  _T_3338 = _T_3337 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3339 = iccm_ecc_word_enable[0] & _T_3338; // @[el2_lib.scala 302:32]
  wire  _T_3341 = _T_3339 & _T_3337[6]; // @[el2_lib.scala 302:53]
  wire  _T_3610 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3611 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3612 = _T_3610 ^ _T_3611; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3620 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3621 = ^_T_3620; // @[el2_lib.scala 301:83]
  wire  _T_3622 = io_iccm_rd_data_ecc[76] ^ _T_3621; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3629 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3637 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3629}; // @[el2_lib.scala 301:103]
  wire  _T_3638 = ^_T_3637; // @[el2_lib.scala 301:110]
  wire  _T_3639 = io_iccm_rd_data_ecc[75] ^ _T_3638; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3646 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3654 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3646}; // @[el2_lib.scala 301:130]
  wire  _T_3655 = ^_T_3654; // @[el2_lib.scala 301:137]
  wire  _T_3656 = io_iccm_rd_data_ecc[74] ^ _T_3655; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3665 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3674 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3665}; // @[el2_lib.scala 301:157]
  wire  _T_3675 = ^_T_3674; // @[el2_lib.scala 301:164]
  wire  _T_3676 = io_iccm_rd_data_ecc[73] ^ _T_3675; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3685 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3694 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3685}; // @[el2_lib.scala 301:184]
  wire  _T_3695 = ^_T_3694; // @[el2_lib.scala 301:191]
  wire  _T_3696 = io_iccm_rd_data_ecc[72] ^ _T_3695; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3705 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3714 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3705}; // @[el2_lib.scala 301:211]
  wire  _T_3715 = ^_T_3714; // @[el2_lib.scala 301:218]
  wire  _T_3716 = io_iccm_rd_data_ecc[71] ^ _T_3715; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3722 = {_T_3612,_T_3622,_T_3639,_T_3656,_T_3676,_T_3696,_T_3716}; // @[Cat.scala 29:58]
  wire  _T_3723 = _T_3722 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3724 = iccm_ecc_word_enable[1] & _T_3723; // @[el2_lib.scala 302:32]
  wire  _T_3726 = _T_3724 & _T_3722[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3341,_T_3726}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 190:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 632:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 192:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 477:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 192:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 192:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 192:72]
  wire  _T_2490 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2495 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2515 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 527:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 391:42]
  wire  _T_2517 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 527:79]
  wire  _T_2518 = _T_2515 | _T_2517; // @[el2_ifu_mem_ctl.scala 527:56]
  wire  _T_2519 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 527:122]
  wire  _T_2520 = ~_T_2519; // @[el2_ifu_mem_ctl.scala 527:101]
  wire  _T_2521 = _T_2518 & _T_2520; // @[el2_ifu_mem_ctl.scala 527:99]
  wire  _T_2522 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2536 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 534:45]
  wire  _T_2537 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 534:69]
  wire  _T_2538 = _T_2536 & _T_2537; // @[el2_ifu_mem_ctl.scala 534:67]
  wire  _T_2539 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_2522 ? _T_2538 : _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2495 ? _T_2521 : _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2490 ? 1'h0 : _GEN_59; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 192:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 194:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 194:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 284:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 284:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 700:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 275:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 325:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 275:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 275:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 284:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 284:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 284:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 284:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 547:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 589:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 616:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 311:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 597:56]
  wire  _T_2641 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 614:69]
  wire  _T_2642 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 614:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2641 : _T_2642; // @[el2_ifu_mem_ctl.scala 614:28]
  wire  _T_2588 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 593:68]
  wire  _T_2589 = ic_act_miss_f | _T_2588; // @[el2_ifu_mem_ctl.scala 593:48]
  wire  bus_reset_data_beat_cnt = _T_2589 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 593:91]
  wire  _T_2585 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 592:50]
  wire  _T_2586 = bus_ifu_wr_en_ff & _T_2585; // @[el2_ifu_mem_ctl.scala 592:48]
  wire  _T_2587 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 592:72]
  wire  bus_inc_data_beat_cnt = _T_2586 & _T_2587; // @[el2_ifu_mem_ctl.scala 592:70]
  wire [2:0] _T_2593 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 596:115]
  wire [2:0] _T_2595 = bus_inc_data_beat_cnt ? _T_2593 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2590 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 594:32]
  wire  _T_2591 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 594:57]
  wire  bus_hold_data_beat_cnt = _T_2590 & _T_2591; // @[el2_ifu_mem_ctl.scala 594:55]
  wire [2:0] _T_2596 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2595 | _T_2596; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 194:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 195:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 194:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 195:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 201:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 427:45]
  wire  _T_2120 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 448:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 404:60]
  wire  _T_2151 = _T_2120 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2124 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2152 = _T_2124 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2159 = _T_2151 | _T_2152; // @[Mux.scala 27:72]
  wire  _T_2128 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2153 = _T_2128 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2160 = _T_2159 | _T_2153; // @[Mux.scala 27:72]
  wire  _T_2132 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2154 = _T_2132 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2161 = _T_2160 | _T_2154; // @[Mux.scala 27:72]
  wire  _T_2136 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2155 = _T_2136 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2162 = _T_2161 | _T_2155; // @[Mux.scala 27:72]
  wire  _T_2140 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2156 = _T_2140 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2163 = _T_2162 | _T_2156; // @[Mux.scala 27:72]
  wire  _T_2144 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2157 = _T_2144 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2164 = _T_2163 | _T_2157; // @[Mux.scala 27:72]
  wire  _T_2148 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2158 = _T_2148 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2164 | _T_2158; // @[Mux.scala 27:72]
  wire  _T_2206 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 450:69]
  wire  _T_2207 = ic_miss_buff_data_valid_bypass_index & _T_2206; // @[el2_ifu_mem_ctl.scala 450:67]
  wire  _T_2209 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 450:91]
  wire  _T_2210 = _T_2207 & _T_2209; // @[el2_ifu_mem_ctl.scala 450:89]
  wire  _T_2215 = _T_2207 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 451:65]
  wire  _T_2216 = _T_2210 | _T_2215; // @[el2_ifu_mem_ctl.scala 450:112]
  wire  _T_2218 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 452:43]
  wire  _T_2221 = _T_2218 & _T_2209; // @[el2_ifu_mem_ctl.scala 452:65]
  wire  _T_2222 = _T_2216 | _T_2221; // @[el2_ifu_mem_ctl.scala 451:88]
  wire  _T_2226 = _T_2218 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 453:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 430:75]
  wire  _T_2166 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2190 = _T_2166 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2169 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2191 = _T_2169 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2190 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2172 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2192 = _T_2172 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2199 = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2193 = _T_2175 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2199 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2178 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2194 = _T_2178 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2181 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2195 = _T_2181 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2184 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2196 = _T_2184 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2187 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2197 = _T_2187 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2227 = _T_2226 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 453:87]
  wire  _T_2228 = _T_2222 | _T_2227; // @[el2_ifu_mem_ctl.scala 452:88]
  wire  _T_2232 = ic_miss_buff_data_valid_bypass_index & _T_2148; // @[el2_ifu_mem_ctl.scala 454:43]
  wire  miss_buff_hit_unq_f = _T_2228 | _T_2232; // @[el2_ifu_mem_ctl.scala 453:131]
  wire  _T_2248 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 459:55]
  wire  _T_2249 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 459:87]
  wire  _T_2250 = _T_2248 | _T_2249; // @[el2_ifu_mem_ctl.scala 459:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2250; // @[el2_ifu_mem_ctl.scala 459:41]
  wire  _T_2233 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 456:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 312:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 447:51]
  wire  _T_2234 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 456:68]
  wire  _T_2235 = miss_buff_hit_unq_f & _T_2234; // @[el2_ifu_mem_ctl.scala 456:66]
  wire  stream_hit_f = _T_2233 & _T_2235; // @[el2_ifu_mem_ctl.scala 456:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 279:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 279:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 599:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 626:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 205:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 205:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 205:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 205:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 207:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 208:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 209:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 209:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 209:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 197:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 209:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 209:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 210:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 210:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 210:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 210:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 211:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 212:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 209:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 208:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 207:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 206:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2245 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 458:60]
  wire  _T_2246 = _T_2245 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 458:94]
  wire  stream_eol_f = _T_2246 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 458:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 220:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 220:87]
  wire  _T_113 = _T_111 & _T_2587; // @[el2_ifu_mem_ctl.scala 220:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 220:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 224:48]
  wire  _T_126 = _T_124 & _T_2587; // @[el2_ifu_mem_ctl.scala 224:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 285:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 285:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 285:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 285:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 285:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 285:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 286:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 339:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 286:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 286:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 286:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:50]
  wire  _T_137 = _T_135 & _T_2587; // @[el2_ifu_mem_ctl.scala 228:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 287:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 288:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 288:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 287:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:35]
  wire  _T_143 = _T_141 & _T_2587; // @[el2_ifu_mem_ctl.scala 229:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 234:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 233:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 238:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 238:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 195:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 195:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 195:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 195:91]
  wire  _T_30 = ic_act_miss_f & _T_2587; // @[el2_ifu_mem_ctl.scala 202:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 213:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 213:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 213:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 213:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 217:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 217:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 221:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 225:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 230:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 235:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 235:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 255:95]
  wire  _T_175 = _T_2248 & _T_174; // @[el2_ifu_mem_ctl.scala 255:93]
  wire  crit_wd_byp_ok_ff = _T_2249 | _T_175; // @[el2_ifu_mem_ctl.scala 255:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 256:36]
  wire  _T_180 = _T_2248 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 256:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 256:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 256:70]
  wire  _T_184 = _T_2248 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 257:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 257:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 256:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 257:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 258:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 258:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 257:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 260:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:35]
  reg [6:0] _T_5166; // @[el2_ifu_mem_ctl.scala 728:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_5166[5:0]; // @[el2_ifu_mem_ctl.scala 727:27]
  wire [6:0] _GEN_473 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 724:121]
  wire  _T_5031 = _GEN_473 == 7'h7f; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5033 = _T_5031 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4522; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_4522[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_474 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5034 = _T_5033 & _GEN_474; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_5027 = _GEN_473 == 7'h7e; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5029 = _T_5027 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4518; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_4518[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_476 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5030 = _T_5029 & _GEN_476; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_5023 = _GEN_473 == 7'h7d; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5025 = _T_5023 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4514; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_4514[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_478 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5026 = _T_5025 & _GEN_478; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_5019 = _GEN_473 == 7'h7c; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5021 = _T_5019 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4510; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_4510[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_480 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5022 = _T_5021 & _GEN_480; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_5015 = _GEN_473 == 7'h7b; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5017 = _T_5015 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4506; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_4506[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_482 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5018 = _T_5017 & _GEN_482; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_5011 = _GEN_473 == 7'h7a; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5013 = _T_5011 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4502; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_4502[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_484 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5014 = _T_5013 & _GEN_484; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_5007 = _GEN_473 == 7'h79; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5009 = _T_5007 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4498; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_4498[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_486 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5010 = _T_5009 & _GEN_486; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_5003 = _GEN_473 == 7'h78; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5005 = _T_5003 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4494; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_4494[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_488 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5006 = _T_5005 & _GEN_488; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4999 = _GEN_473 == 7'h77; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_5001 = _T_4999 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4490; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_4490[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_490 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_5002 = _T_5001 & _GEN_490; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4995 = _GEN_473 == 7'h76; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4997 = _T_4995 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4486; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_4486[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_492 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4998 = _T_4997 & _GEN_492; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [59:0] _T_5043 = {_T_5034,_T_5030,_T_5026,_T_5022,_T_5018,_T_5014,_T_5010,_T_5006,_T_5002,_T_4998}; // @[Cat.scala 29:58]
  wire  _T_4991 = _GEN_473 == 7'h75; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4993 = _T_4991 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4482; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_4482[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_494 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4994 = _T_4993 & _GEN_494; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4987 = _GEN_473 == 7'h74; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4989 = _T_4987 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4478; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_4478[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_496 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4990 = _T_4989 & _GEN_496; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4983 = _GEN_473 == 7'h73; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4985 = _T_4983 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4474; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_4474[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_498 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4986 = _T_4985 & _GEN_498; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4979 = _GEN_473 == 7'h72; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4981 = _T_4979 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4470; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_4470[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_500 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4982 = _T_4981 & _GEN_500; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4975 = _GEN_473 == 7'h71; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4977 = _T_4975 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4466; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_4466[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_502 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4978 = _T_4977 & _GEN_502; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4971 = _GEN_473 == 7'h70; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4973 = _T_4971 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4462; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_4462[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_504 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4974 = _T_4973 & _GEN_504; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4967 = _GEN_473 == 7'h6f; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4969 = _T_4967 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4458; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_4458[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_506 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4970 = _T_4969 & _GEN_506; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4963 = _GEN_473 == 7'h6e; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4965 = _T_4963 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4454; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_4454[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_508 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4966 = _T_4965 & _GEN_508; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4959 = _GEN_473 == 7'h6d; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4961 = _T_4959 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4450; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_4450[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_510 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4962 = _T_4961 & _GEN_510; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [113:0] _T_5052 = {_T_5043,_T_4994,_T_4990,_T_4986,_T_4982,_T_4978,_T_4974,_T_4970,_T_4966,_T_4962}; // @[Cat.scala 29:58]
  wire  _T_4955 = _GEN_473 == 7'h6c; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4957 = _T_4955 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4446; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_4446[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_512 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4958 = _T_4957 & _GEN_512; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4951 = _GEN_473 == 7'h6b; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4953 = _T_4951 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4442; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_4442[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_514 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4954 = _T_4953 & _GEN_514; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4947 = _GEN_473 == 7'h6a; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4949 = _T_4947 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4438; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_4438[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_516 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4950 = _T_4949 & _GEN_516; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4943 = _GEN_473 == 7'h69; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4945 = _T_4943 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4434; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_4434[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_518 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4946 = _T_4945 & _GEN_518; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4939 = _GEN_473 == 7'h68; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4941 = _T_4939 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4430; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_4430[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_520 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4942 = _T_4941 & _GEN_520; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4935 = _GEN_473 == 7'h67; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4937 = _T_4935 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4426; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_4426[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_522 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4938 = _T_4937 & _GEN_522; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4931 = _GEN_473 == 7'h66; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4933 = _T_4931 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4422; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_4422[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_524 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4934 = _T_4933 & _GEN_524; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4927 = _GEN_473 == 7'h65; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4929 = _T_4927 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4418; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_4418[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_526 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4930 = _T_4929 & _GEN_526; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4923 = _GEN_473 == 7'h64; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4925 = _T_4923 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4414; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_4414[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_528 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4926 = _T_4925 & _GEN_528; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [167:0] _T_5061 = {_T_5052,_T_4958,_T_4954,_T_4950,_T_4946,_T_4942,_T_4938,_T_4934,_T_4930,_T_4926}; // @[Cat.scala 29:58]
  wire  _T_4919 = _GEN_473 == 7'h63; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4921 = _T_4919 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4410; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_4410[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_530 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4922 = _T_4921 & _GEN_530; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4915 = _GEN_473 == 7'h62; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4917 = _T_4915 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4406; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_4406[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_532 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4918 = _T_4917 & _GEN_532; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4911 = _GEN_473 == 7'h61; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4913 = _T_4911 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4402; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_4402[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_534 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4914 = _T_4913 & _GEN_534; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4907 = _GEN_473 == 7'h60; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4909 = _T_4907 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4398; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_4398[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_536 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4910 = _T_4909 & _GEN_536; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4903 = _GEN_473 == 7'h5f; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4905 = _T_4903 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4394; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_4394[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_538 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4906 = _T_4905 & _GEN_538; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4899 = _GEN_473 == 7'h5e; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4901 = _T_4899 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4390; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_4390[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_540 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4902 = _T_4901 & _GEN_540; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4895 = _GEN_473 == 7'h5d; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4897 = _T_4895 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4386; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_4386[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_542 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4898 = _T_4897 & _GEN_542; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4891 = _GEN_473 == 7'h5c; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4893 = _T_4891 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4382; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_4382[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_544 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4894 = _T_4893 & _GEN_544; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4887 = _GEN_473 == 7'h5b; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4889 = _T_4887 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4378; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_4378[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_546 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4890 = _T_4889 & _GEN_546; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [221:0] _T_5070 = {_T_5061,_T_4922,_T_4918,_T_4914,_T_4910,_T_4906,_T_4902,_T_4898,_T_4894,_T_4890}; // @[Cat.scala 29:58]
  wire  _T_4883 = _GEN_473 == 7'h5a; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4885 = _T_4883 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4374; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_4374[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_548 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4886 = _T_4885 & _GEN_548; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4879 = _GEN_473 == 7'h59; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4881 = _T_4879 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4370; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_4370[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_550 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4882 = _T_4881 & _GEN_550; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4875 = _GEN_473 == 7'h58; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4877 = _T_4875 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4366; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_4366[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_552 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4878 = _T_4877 & _GEN_552; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4871 = _GEN_473 == 7'h57; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4873 = _T_4871 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4362; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_4362[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_554 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4874 = _T_4873 & _GEN_554; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4867 = _GEN_473 == 7'h56; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4869 = _T_4867 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4358; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_4358[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_556 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4870 = _T_4869 & _GEN_556; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4863 = _GEN_473 == 7'h55; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4865 = _T_4863 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4354; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_4354[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_558 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4866 = _T_4865 & _GEN_558; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4859 = _GEN_473 == 7'h54; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4861 = _T_4859 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4350; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_4350[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_560 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4862 = _T_4861 & _GEN_560; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4855 = _GEN_473 == 7'h53; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4857 = _T_4855 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4346; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_4346[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_562 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4858 = _T_4857 & _GEN_562; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4851 = _GEN_473 == 7'h52; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4853 = _T_4851 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4342; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_4342[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_564 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4854 = _T_4853 & _GEN_564; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [275:0] _T_5079 = {_T_5070,_T_4886,_T_4882,_T_4878,_T_4874,_T_4870,_T_4866,_T_4862,_T_4858,_T_4854}; // @[Cat.scala 29:58]
  wire  _T_4847 = _GEN_473 == 7'h51; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4849 = _T_4847 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4338; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_4338[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_566 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4850 = _T_4849 & _GEN_566; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4843 = _GEN_473 == 7'h50; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4845 = _T_4843 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4334; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_4334[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_568 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4846 = _T_4845 & _GEN_568; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4839 = _GEN_473 == 7'h4f; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4841 = _T_4839 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4330; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_4330[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_570 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4842 = _T_4841 & _GEN_570; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4835 = _GEN_473 == 7'h4e; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4837 = _T_4835 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4326; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_4326[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_572 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4838 = _T_4837 & _GEN_572; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4831 = _GEN_473 == 7'h4d; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4833 = _T_4831 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4322; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_4322[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_574 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4834 = _T_4833 & _GEN_574; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4827 = _GEN_473 == 7'h4c; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4829 = _T_4827 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4318; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_4318[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_576 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4830 = _T_4829 & _GEN_576; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4823 = _GEN_473 == 7'h4b; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4825 = _T_4823 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4314; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_4314[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_578 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4826 = _T_4825 & _GEN_578; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4819 = _GEN_473 == 7'h4a; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4821 = _T_4819 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4310; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_4310[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_580 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4822 = _T_4821 & _GEN_580; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4815 = _GEN_473 == 7'h49; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4817 = _T_4815 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4306; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_4306[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_582 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4818 = _T_4817 & _GEN_582; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [329:0] _T_5088 = {_T_5079,_T_4850,_T_4846,_T_4842,_T_4838,_T_4834,_T_4830,_T_4826,_T_4822,_T_4818}; // @[Cat.scala 29:58]
  wire  _T_4811 = _GEN_473 == 7'h48; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4813 = _T_4811 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4302; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_4302[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_584 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4814 = _T_4813 & _GEN_584; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4807 = _GEN_473 == 7'h47; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4809 = _T_4807 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4298; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_4298[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_586 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4810 = _T_4809 & _GEN_586; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4803 = _GEN_473 == 7'h46; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4805 = _T_4803 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4294; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_4294[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_588 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4806 = _T_4805 & _GEN_588; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4799 = _GEN_473 == 7'h45; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4801 = _T_4799 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4290; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_4290[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_590 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4802 = _T_4801 & _GEN_590; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4795 = _GEN_473 == 7'h44; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4797 = _T_4795 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4286; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_4286[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_592 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4798 = _T_4797 & _GEN_592; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4791 = _GEN_473 == 7'h43; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4793 = _T_4791 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4282; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_4282[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_594 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4794 = _T_4793 & _GEN_594; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4787 = _GEN_473 == 7'h42; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4789 = _T_4787 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4278; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_4278[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_596 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4790 = _T_4789 & _GEN_596; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4783 = _GEN_473 == 7'h41; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4785 = _T_4783 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4274; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_4274[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_598 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4786 = _T_4785 & _GEN_598; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4779 = _GEN_473 == 7'h40; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4781 = _T_4779 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4270; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_4270[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4782 = _T_4781 & _GEN_600; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [383:0] _T_5097 = {_T_5088,_T_4814,_T_4810,_T_4806,_T_4802,_T_4798,_T_4794,_T_4790,_T_4786,_T_4782}; // @[Cat.scala 29:58]
  wire  _T_4775 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4777 = _T_4775 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4266; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_4266[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4778 = _T_4777 & _GEN_601; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4771 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4773 = _T_4771 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4262; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_4262[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4774 = _T_4773 & _GEN_602; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4767 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4769 = _T_4767 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4258; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_4258[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4770 = _T_4769 & _GEN_603; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4763 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4765 = _T_4763 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4254; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_4254[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4766 = _T_4765 & _GEN_604; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4759 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4761 = _T_4759 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4250; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_4250[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4762 = _T_4761 & _GEN_605; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4755 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4757 = _T_4755 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4246; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_4246[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4758 = _T_4757 & _GEN_606; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4751 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4753 = _T_4751 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4242; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_4242[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4754 = _T_4753 & _GEN_607; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4747 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4749 = _T_4747 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4238; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_4238[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4750 = _T_4749 & _GEN_608; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4743 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4745 = _T_4743 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4234; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_4234[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4746 = _T_4745 & _GEN_609; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [437:0] _T_5106 = {_T_5097,_T_4778,_T_4774,_T_4770,_T_4766,_T_4762,_T_4758,_T_4754,_T_4750,_T_4746}; // @[Cat.scala 29:58]
  wire  _T_4739 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4741 = _T_4739 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4230; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_4230[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4742 = _T_4741 & _GEN_610; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4735 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4737 = _T_4735 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4226; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_4226[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4738 = _T_4737 & _GEN_611; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4731 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4733 = _T_4731 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4222; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_4222[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4734 = _T_4733 & _GEN_612; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4727 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4729 = _T_4727 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4218; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_4218[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4730 = _T_4729 & _GEN_613; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4723 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4725 = _T_4723 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4214; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_4214[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4726 = _T_4725 & _GEN_614; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4719 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4721 = _T_4719 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4210; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_4210[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4722 = _T_4721 & _GEN_615; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4715 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4717 = _T_4715 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4206; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_4206[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4718 = _T_4717 & _GEN_616; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4711 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4713 = _T_4711 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4202; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_4202[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4714 = _T_4713 & _GEN_617; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4707 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4709 = _T_4707 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4198; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_4198[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4710 = _T_4709 & _GEN_618; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [491:0] _T_5115 = {_T_5106,_T_4742,_T_4738,_T_4734,_T_4730,_T_4726,_T_4722,_T_4718,_T_4714,_T_4710}; // @[Cat.scala 29:58]
  wire  _T_4703 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4705 = _T_4703 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4194; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_4194[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4706 = _T_4705 & _GEN_619; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4699 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4701 = _T_4699 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4190; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_4190[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4702 = _T_4701 & _GEN_620; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4695 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4697 = _T_4695 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4186; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_4186[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4698 = _T_4697 & _GEN_621; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4691 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4693 = _T_4691 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4182; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_4182[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4694 = _T_4693 & _GEN_622; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4687 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4689 = _T_4687 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4178; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_4178[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4690 = _T_4689 & _GEN_623; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4683 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4685 = _T_4683 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4174; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_4174[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4686 = _T_4685 & _GEN_624; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4679 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4681 = _T_4679 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4170; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_4170[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4682 = _T_4681 & _GEN_625; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4675 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4677 = _T_4675 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4166; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_4166[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4678 = _T_4677 & _GEN_626; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4671 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4673 = _T_4671 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4162; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_4162[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4674 = _T_4673 & _GEN_627; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [545:0] _T_5124 = {_T_5115,_T_4706,_T_4702,_T_4698,_T_4694,_T_4690,_T_4686,_T_4682,_T_4678,_T_4674}; // @[Cat.scala 29:58]
  wire  _T_4667 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4669 = _T_4667 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4158; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_4158[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4670 = _T_4669 & _GEN_628; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4663 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4665 = _T_4663 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4154; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_4154[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4666 = _T_4665 & _GEN_629; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4659 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4661 = _T_4659 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4150; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_4150[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4662 = _T_4661 & _GEN_630; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4655 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4657 = _T_4655 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4146; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_4146[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4658 = _T_4657 & _GEN_631; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4651 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4653 = _T_4651 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4142; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_4142[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4654 = _T_4653 & _GEN_632; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4647 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4649 = _T_4647 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4138; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_4138[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4650 = _T_4649 & _GEN_633; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4643 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4645 = _T_4643 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4134; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_4134[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4646 = _T_4645 & _GEN_634; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4639 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4641 = _T_4639 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4130; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_4130[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4642 = _T_4641 & _GEN_635; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4635 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4637 = _T_4635 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4126; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_4126[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4638 = _T_4637 & _GEN_636; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [599:0] _T_5133 = {_T_5124,_T_4670,_T_4666,_T_4662,_T_4658,_T_4654,_T_4650,_T_4646,_T_4642,_T_4638}; // @[Cat.scala 29:58]
  wire  _T_4631 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4633 = _T_4631 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4122; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_4122[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4634 = _T_4633 & _GEN_637; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4627 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4629 = _T_4627 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4118; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_4118[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4630 = _T_4629 & _GEN_638; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4623 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4625 = _T_4623 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4114; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_4114[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4626 = _T_4625 & _GEN_639; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4619 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4621 = _T_4619 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4110; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_4110[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4622 = _T_4621 & _GEN_640; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4615 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4617 = _T_4615 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4106; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_4106[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4618 = _T_4617 & _GEN_641; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4611 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4613 = _T_4611 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4102; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_4102[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4614 = _T_4613 & _GEN_642; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4607 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4609 = _T_4607 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4098; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_4098[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4610 = _T_4609 & _GEN_643; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4603 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4605 = _T_4603 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4094; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_4094[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4606 = _T_4605 & _GEN_644; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4599 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4601 = _T_4599 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4090; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_4090[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4602 = _T_4601 & _GEN_645; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [653:0] _T_5142 = {_T_5133,_T_4634,_T_4630,_T_4626,_T_4622,_T_4618,_T_4614,_T_4610,_T_4606,_T_4602}; // @[Cat.scala 29:58]
  wire  _T_4595 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4597 = _T_4595 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4086; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_4086[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4598 = _T_4597 & _GEN_646; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4591 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4593 = _T_4591 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4082; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_4082[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4594 = _T_4593 & _GEN_647; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4587 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4589 = _T_4587 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4078; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_4078[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4590 = _T_4589 & _GEN_648; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4583 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4585 = _T_4583 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4074; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_4074[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4586 = _T_4585 & _GEN_649; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4579 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4581 = _T_4579 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4070; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_4070[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4582 = _T_4581 & _GEN_650; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4575 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4577 = _T_4575 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4066; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_4066[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4578 = _T_4577 & _GEN_651; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4571 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4573 = _T_4571 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4062; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_4062[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4574 = _T_4573 & _GEN_652; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4567 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4569 = _T_4567 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4058; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_4058[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4570 = _T_4569 & _GEN_653; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4563 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4565 = _T_4563 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4054; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_4054[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4566 = _T_4565 & _GEN_654; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [707:0] _T_5151 = {_T_5142,_T_4598,_T_4594,_T_4590,_T_4586,_T_4582,_T_4578,_T_4574,_T_4570,_T_4566}; // @[Cat.scala 29:58]
  wire  _T_4559 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4561 = _T_4559 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4050; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_4050[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4562 = _T_4561 & _GEN_655; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4555 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4557 = _T_4555 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4046; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_4046[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4558 = _T_4557 & _GEN_656; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4551 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4553 = _T_4551 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4042; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_4042[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4554 = _T_4553 & _GEN_657; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4547 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4549 = _T_4547 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4038; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_4038[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4550 = _T_4549 & _GEN_658; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4543 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4545 = _T_4543 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4034; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_4034[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4546 = _T_4545 & _GEN_659; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4539 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4541 = _T_4539 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4030; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_4030[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4542 = _T_4541 & _GEN_660; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4535 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4537 = _T_4535 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4026; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_4026[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4538 = _T_4537 & _GEN_661; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4531 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4533 = _T_4531 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4022; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_4022[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4534 = _T_4533 & _GEN_662; // @[el2_ifu_mem_ctl.scala 724:130]
  wire  _T_4527 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4529 = _T_4527 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4018; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_4018[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4530 = _T_4529 & _GEN_663; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [761:0] _T_5160 = {_T_5151,_T_4562,_T_4558,_T_4554,_T_4550,_T_4546,_T_4542,_T_4538,_T_4534,_T_4530}; // @[Cat.scala 29:58]
  wire  _T_4523 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 724:121]
  wire [5:0] _T_4525 = _T_4523 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4014; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_4014[0]; // @[el2_ifu_mem_ctl.scala 721:30 el2_ifu_mem_ctl.scala 723:33]
  wire [5:0] _GEN_664 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [5:0] _T_4526 = _T_4525 & _GEN_664; // @[el2_ifu_mem_ctl.scala 724:130]
  wire [767:0] _T_5161 = {_T_5160,_T_4526}; // @[Cat.scala 29:58]
  wire  way_status = _T_5161[0]; // @[el2_ifu_mem_ctl.scala 724:16]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 263:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 265:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 272:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 277:59]
  wire  _T_214 = _T_212 | _T_2233; // @[el2_ifu_mem_ctl.scala 277:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 277:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 283:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 283:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 283:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 290:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 290:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 290:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 291:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 291:32]
  wire  _T_274 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 294:75]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 294:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2662 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 622:48]
  wire  _T_2663 = _T_2662 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 622:52]
  wire  bus_ifu_wr_data_error_ff = _T_2663 & miss_pending; // @[el2_ifu_mem_ctl.scala 622:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 367:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 366:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 294:145]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 294:143]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 297:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 298:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 317:30]
  wire  _T_10367 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 777:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 318:24]
  wire  _T_10369 = _T_10367 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 777:51]
  wire  _T_10371 = _T_10369 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 777:67]
  wire  _T_10373 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 777:86]
  wire  replace_way_mb_any_0 = _T_10371 | _T_10373; // @[el2_ifu_mem_ctl.scala 777:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10376 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 778:50]
  wire  _T_10378 = _T_10376 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 778:66]
  wire  _T_10380 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 778:85]
  wire  _T_10382 = _T_10380 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 778:100]
  wire  replace_way_mb_any_1 = _T_10378 | _T_10382; // @[el2_ifu_mem_ctl.scala 778:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 302:110]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 306:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 306:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 307:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 306:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 308:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 316:23]
  wire  _T_313 = _T_2248 & flush_final_f; // @[el2_ifu_mem_ctl.scala 320:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 320:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 320:53]
  wire  _T_2240 = ~_T_2235; // @[el2_ifu_mem_ctl.scala 457:46]
  wire  _T_2241 = _T_2233 & _T_2240; // @[el2_ifu_mem_ctl.scala 457:44]
  wire  stream_miss_f = _T_2241 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 457:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 320:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 320:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 326:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_2233; // @[el2_ifu_mem_ctl.scala 328:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 328:82]
  wire  _T_2254 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 462:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2254}; // @[Cat.scala 29:58]
  wire  _T_2255 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2279 = _T_2255 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2258 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2280 = _T_2258 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2287 = _T_2279 | _T_2280; // @[Mux.scala 27:72]
  wire  _T_2261 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2281 = _T_2261 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2287 | _T_2281; // @[Mux.scala 27:72]
  wire  _T_2264 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2282 = _T_2264 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2288 | _T_2282; // @[Mux.scala 27:72]
  wire  _T_2267 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2283 = _T_2267 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2289 | _T_2283; // @[Mux.scala 27:72]
  wire  _T_2270 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2284 = _T_2270 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2290 | _T_2284; // @[Mux.scala 27:72]
  wire  _T_2273 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2285 = _T_2273 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2291 | _T_2285; // @[Mux.scala 27:72]
  wire  _T_2276 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2286 = _T_2276 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2292 | _T_2286; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 464:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 332:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 332:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 619:61]
  wire  _T_2656 = ic_act_miss_f_delayed & _T_2249; // @[el2_ifu_mem_ctl.scala 620:53]
  wire  reset_tag_valid_for_miss = _T_2656 & _T_17; // @[el2_ifu_mem_ctl.scala 620:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 332:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 334:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 336:84]
  wire  _T_2650 = ~_T_2662; // @[el2_ifu_mem_ctl.scala 617:84]
  wire  _T_2651 = _T_100 & _T_2650; // @[el2_ifu_mem_ctl.scala 617:82]
  wire  bus_ifu_wr_en_ff_q = _T_2651 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 617:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 336:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 337:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_567 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 384:13]
  wire  _T_568 = ^_T_567; // @[el2_lib.scala 384:20]
  wire [6:0] _T_574 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_581 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 384:30]
  wire [14:0] _T_582 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_574}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_589 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 384:30]
  wire [30:0] _T_598 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_582}; // @[el2_lib.scala 384:30]
  wire  _T_599 = ^_T_598; // @[el2_lib.scala 384:37]
  wire [6:0] _T_605 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 384:47]
  wire [14:0] _T_613 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_605}; // @[el2_lib.scala 384:47]
  wire [30:0] _T_629 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_613}; // @[el2_lib.scala 384:47]
  wire  _T_630 = ^_T_629; // @[el2_lib.scala 384:54]
  wire [6:0] _T_636 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 384:64]
  wire [14:0] _T_644 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_636}; // @[el2_lib.scala 384:64]
  wire [30:0] _T_660 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_581,_T_644}; // @[el2_lib.scala 384:64]
  wire  _T_661 = ^_T_660; // @[el2_lib.scala 384:71]
  wire [7:0] _T_668 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 384:81]
  wire [16:0] _T_677 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_668}; // @[el2_lib.scala 384:81]
  wire [8:0] _T_685 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 384:81]
  wire [17:0] _T_694 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_685}; // @[el2_lib.scala 384:81]
  wire [34:0] _T_695 = {_T_694,_T_677}; // @[el2_lib.scala 384:81]
  wire  _T_696 = ^_T_695; // @[el2_lib.scala 384:88]
  wire [7:0] _T_703 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 384:98]
  wire [16:0] _T_712 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_703}; // @[el2_lib.scala 384:98]
  wire [8:0] _T_720 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 384:98]
  wire [17:0] _T_729 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_720}; // @[el2_lib.scala 384:98]
  wire [34:0] _T_730 = {_T_729,_T_712}; // @[el2_lib.scala 384:98]
  wire  _T_731 = ^_T_730; // @[el2_lib.scala 384:105]
  wire [7:0] _T_738 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 384:115]
  wire [16:0] _T_747 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_738}; // @[el2_lib.scala 384:115]
  wire [8:0] _T_755 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 384:115]
  wire [17:0] _T_764 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_755}; // @[el2_lib.scala 384:115]
  wire [34:0] _T_765 = {_T_764,_T_747}; // @[el2_lib.scala 384:115]
  wire  _T_766 = ^_T_765; // @[el2_lib.scala 384:122]
  wire [3:0] _T_2295 = {ifu_bus_rid_ff[2:1],_T_2254,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2296 = _T_2295 == 4'h0; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2343 = _T_2296 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2299 = _T_2295 == 4'h1; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2344 = _T_2299 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2343 | _T_2344; // @[Mux.scala 27:72]
  wire  _T_2302 = _T_2295 == 4'h2; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2345 = _T_2302 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2360 = _T_2359 | _T_2345; // @[Mux.scala 27:72]
  wire  _T_2305 = _T_2295 == 4'h3; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2346 = _T_2305 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2360 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2308 = _T_2295 == 4'h4; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2347 = _T_2308 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire  _T_2311 = _T_2295 == 4'h5; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2348 = _T_2311 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2363 = _T_2362 | _T_2348; // @[Mux.scala 27:72]
  wire  _T_2314 = _T_2295 == 4'h6; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2349 = _T_2314 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2364 = _T_2363 | _T_2349; // @[Mux.scala 27:72]
  wire  _T_2317 = _T_2295 == 4'h7; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2350 = _T_2317 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2365 = _T_2364 | _T_2350; // @[Mux.scala 27:72]
  wire  _T_2320 = _T_2295 == 4'h8; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2351 = _T_2320 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2366 = _T_2365 | _T_2351; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2295 == 4'h9; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2352 = _T_2323 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2367 = _T_2366 | _T_2352; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2295 == 4'ha; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2353 = _T_2326 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2368 = _T_2367 | _T_2353; // @[Mux.scala 27:72]
  wire  _T_2329 = _T_2295 == 4'hb; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2354 = _T_2329 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2369 = _T_2368 | _T_2354; // @[Mux.scala 27:72]
  wire  _T_2332 = _T_2295 == 4'hc; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2355 = _T_2332 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 27:72]
  wire  _T_2335 = _T_2295 == 4'hd; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2356 = _T_2335 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2371 = _T_2370 | _T_2356; // @[Mux.scala 27:72]
  wire  _T_2338 = _T_2295 == 4'he; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2357 = _T_2338 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2372 = _T_2371 | _T_2357; // @[Mux.scala 27:72]
  wire  _T_2341 = _T_2295 == 4'hf; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2358 = _T_2341 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2373 = _T_2372 | _T_2358; // @[Mux.scala 27:72]
  wire [3:0] _T_2375 = {ifu_bus_rid_ff[2:1],_T_2254,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2376 = _T_2375 == 4'h0; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2423 = _T_2376 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2375 == 4'h1; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2424 = _T_2379 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2439 = _T_2423 | _T_2424; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2375 == 4'h2; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2425 = _T_2382 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2440 = _T_2439 | _T_2425; // @[Mux.scala 27:72]
  wire  _T_2385 = _T_2375 == 4'h3; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2426 = _T_2385 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2441 = _T_2440 | _T_2426; // @[Mux.scala 27:72]
  wire  _T_2388 = _T_2375 == 4'h4; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2427 = _T_2388 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2442 = _T_2441 | _T_2427; // @[Mux.scala 27:72]
  wire  _T_2391 = _T_2375 == 4'h5; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2428 = _T_2391 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2443 = _T_2442 | _T_2428; // @[Mux.scala 27:72]
  wire  _T_2394 = _T_2375 == 4'h6; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2429 = _T_2394 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2444 = _T_2443 | _T_2429; // @[Mux.scala 27:72]
  wire  _T_2397 = _T_2375 == 4'h7; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2430 = _T_2397 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2445 = _T_2444 | _T_2430; // @[Mux.scala 27:72]
  wire  _T_2400 = _T_2375 == 4'h8; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2431 = _T_2400 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2446 = _T_2445 | _T_2431; // @[Mux.scala 27:72]
  wire  _T_2403 = _T_2375 == 4'h9; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2432 = _T_2403 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2447 = _T_2446 | _T_2432; // @[Mux.scala 27:72]
  wire  _T_2406 = _T_2375 == 4'ha; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2433 = _T_2406 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2448 = _T_2447 | _T_2433; // @[Mux.scala 27:72]
  wire  _T_2409 = _T_2375 == 4'hb; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2434 = _T_2409 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2449 = _T_2448 | _T_2434; // @[Mux.scala 27:72]
  wire  _T_2412 = _T_2375 == 4'hc; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2435 = _T_2412 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2450 = _T_2449 | _T_2435; // @[Mux.scala 27:72]
  wire  _T_2415 = _T_2375 == 4'hd; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2436 = _T_2415 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2451 = _T_2450 | _T_2436; // @[Mux.scala 27:72]
  wire  _T_2418 = _T_2375 == 4'he; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2437 = _T_2418 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2452 = _T_2451 | _T_2437; // @[Mux.scala 27:72]
  wire  _T_2421 = _T_2375 == 4'hf; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2438 = _T_2421 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2453 = _T_2452 | _T_2438; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [6:0] _T_989 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 384:13]
  wire  _T_990 = ^_T_989; // @[el2_lib.scala 384:20]
  wire [6:0] _T_996 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_1003 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 384:30]
  wire [14:0] _T_1004 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_996}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_1011 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 384:30]
  wire [30:0] _T_1020 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1004}; // @[el2_lib.scala 384:30]
  wire  _T_1021 = ^_T_1020; // @[el2_lib.scala 384:37]
  wire [6:0] _T_1027 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 384:47]
  wire [14:0] _T_1035 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1027}; // @[el2_lib.scala 384:47]
  wire [30:0] _T_1051 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1035}; // @[el2_lib.scala 384:47]
  wire  _T_1052 = ^_T_1051; // @[el2_lib.scala 384:54]
  wire [6:0] _T_1058 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 384:64]
  wire [14:0] _T_1066 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1058}; // @[el2_lib.scala 384:64]
  wire [30:0] _T_1082 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1003,_T_1066}; // @[el2_lib.scala 384:64]
  wire  _T_1083 = ^_T_1082; // @[el2_lib.scala 384:71]
  wire [7:0] _T_1090 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 384:81]
  wire [16:0] _T_1099 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1090}; // @[el2_lib.scala 384:81]
  wire [8:0] _T_1107 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 384:81]
  wire [17:0] _T_1116 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1107}; // @[el2_lib.scala 384:81]
  wire [34:0] _T_1117 = {_T_1116,_T_1099}; // @[el2_lib.scala 384:81]
  wire  _T_1118 = ^_T_1117; // @[el2_lib.scala 384:88]
  wire [7:0] _T_1125 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 384:98]
  wire [16:0] _T_1134 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1125}; // @[el2_lib.scala 384:98]
  wire [8:0] _T_1142 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 384:98]
  wire [17:0] _T_1151 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1142}; // @[el2_lib.scala 384:98]
  wire [34:0] _T_1152 = {_T_1151,_T_1134}; // @[el2_lib.scala 384:98]
  wire  _T_1153 = ^_T_1152; // @[el2_lib.scala 384:105]
  wire [7:0] _T_1160 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 384:115]
  wire [16:0] _T_1169 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1160}; // @[el2_lib.scala 384:115]
  wire [8:0] _T_1177 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 384:115]
  wire [17:0] _T_1186 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1177}; // @[el2_lib.scala 384:115]
  wire [34:0] _T_1187 = {_T_1186,_T_1169}; // @[el2_lib.scala 384:115]
  wire  _T_1188 = ^_T_1187; // @[el2_lib.scala 384:122]
  wire [70:0] _T_1233 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1232 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [141:0] _T_1234 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff,_T_1232}; // @[Cat.scala 29:58]
  wire [141:0] _T_1237 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453,_T_1233}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1234 : _T_1237; // @[el2_ifu_mem_ctl.scala 358:28]
  wire  _T_1196 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 348:56]
  wire  _T_1197 = _T_1196 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 348:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 412:28]
  wire  _T_1413 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 615:35]
  wire  _T_1282 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1339 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 403:118]
  wire  _T_1340 = ic_miss_buff_data_valid[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1340; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1436 = _T_1413 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1343 = ic_miss_buff_data_valid[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1343; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1437 = _T_1416 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1444 = _T_1436 | _T_1437; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1284 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1346 = ic_miss_buff_data_valid[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1346; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1438 = _T_1419 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1444 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1349 = ic_miss_buff_data_valid[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1349; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1439 = _T_1422 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1425 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1352 = ic_miss_buff_data_valid[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1352; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1440 = _T_1425 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1428 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1355 = ic_miss_buff_data_valid[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1355; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1441 = _T_1428 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1431 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1358 = ic_miss_buff_data_valid[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1358; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1442 = _T_1431 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1434 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1361 = ic_miss_buff_data_valid[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1361; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1443 = _T_1434 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1452 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 415:58]
  wire  _T_1453 = bypass_valid_value_check & _T_1452; // @[el2_ifu_mem_ctl.scala 415:56]
  wire  _T_1455 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 415:77]
  wire  _T_1456 = _T_1453 & _T_1455; // @[el2_ifu_mem_ctl.scala 415:75]
  wire  _T_1461 = _T_1453 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 416:75]
  wire  _T_1462 = _T_1456 | _T_1461; // @[el2_ifu_mem_ctl.scala 415:95]
  wire  _T_1464 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 417:56]
  wire  _T_1467 = _T_1464 & _T_1455; // @[el2_ifu_mem_ctl.scala 417:74]
  wire  _T_1468 = _T_1462 | _T_1467; // @[el2_ifu_mem_ctl.scala 416:94]
  wire  _T_1472 = _T_1464 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 418:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 413:70]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1489 = _T_1473 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1490 = _T_1475 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1497 = _T_1489 | _T_1490; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1491 = _T_1477 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1498 = _T_1497 | _T_1491; // @[Mux.scala 27:72]
  wire  _T_1479 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1492 = _T_1479 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1498 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1481 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1493 = _T_1481 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1499 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1483 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1494 = _T_1483 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1500 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1485 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1495 = _T_1485 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1501 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1487 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1496 = _T_1487 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1502 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1472 & _T_1503; // @[el2_ifu_mem_ctl.scala 418:69]
  wire  _T_1506 = _T_1468 | _T_1505; // @[el2_ifu_mem_ctl.scala 417:94]
  wire [4:0] _GEN_665 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 419:95]
  wire  _T_1509 = _GEN_665 == 5'h1f; // @[el2_ifu_mem_ctl.scala 419:95]
  wire  _T_1510 = bypass_valid_value_check & _T_1509; // @[el2_ifu_mem_ctl.scala 419:56]
  wire  bypass_data_ready_in = _T_1506 | _T_1510; // @[el2_ifu_mem_ctl.scala 418:181]
  wire  _T_1511 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 423:53]
  wire  _T_1512 = _T_1511 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 423:73]
  wire  _T_1514 = _T_1512 & _T_317; // @[el2_ifu_mem_ctl.scala 423:96]
  wire  _T_1516 = _T_1514 & _T_58; // @[el2_ifu_mem_ctl.scala 423:118]
  wire  _T_1518 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 424:73]
  wire  _T_1520 = _T_1518 & _T_317; // @[el2_ifu_mem_ctl.scala 424:96]
  wire  _T_1522 = _T_1520 & _T_58; // @[el2_ifu_mem_ctl.scala 424:118]
  wire  _T_1523 = _T_1516 | _T_1522; // @[el2_ifu_mem_ctl.scala 423:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 426:58]
  wire  _T_1524 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 425:54]
  wire  _T_1525 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 425:76]
  wire  _T_1526 = _T_1524 & _T_1525; // @[el2_ifu_mem_ctl.scala 425:74]
  wire  _T_1528 = _T_1526 & _T_317; // @[el2_ifu_mem_ctl.scala 425:96]
  wire  ic_crit_wd_rdy_new_in = _T_1523 | _T_1528; // @[el2_ifu_mem_ctl.scala 424:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 625:43]
  wire  _T_1249 = ic_crit_wd_rdy | _T_2233; // @[el2_ifu_mem_ctl.scala 371:38]
  wire  _T_1251 = _T_1249 | _T_2249; // @[el2_ifu_mem_ctl.scala 371:64]
  wire  _T_1252 = ~_T_1251; // @[el2_ifu_mem_ctl.scala 371:21]
  wire  _T_1253 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 371:98]
  wire  sel_ic_data = _T_1252 & _T_1253; // @[el2_ifu_mem_ctl.scala 371:96]
  wire  _T_2456 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 470:44]
  wire  _T_1622 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 437:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 409:60]
  wire  _T_1566 = _T_1413 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1416 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1566 | _T_1567; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1419 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1574 | _T_1568; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1422 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1575 | _T_1569; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1425 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1570; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1428 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1571; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1431 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1572; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1434 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1579 | _T_1573; // @[Mux.scala 27:72]
  wire  _T_1605 = _T_2166 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1606 = _T_2169 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1613 = _T_1605 | _T_1606; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_2172 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1614 = _T_1613 | _T_1607; // @[Mux.scala 27:72]
  wire  _T_1608 = _T_2175 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1615 = _T_1614 | _T_1608; // @[Mux.scala 27:72]
  wire  _T_1609 = _T_2178 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1616 = _T_1615 | _T_1609; // @[Mux.scala 27:72]
  wire  _T_1610 = _T_2181 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1617 = _T_1616 | _T_1610; // @[Mux.scala 27:72]
  wire  _T_1611 = _T_2184 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1618 = _T_1617 | _T_1611; // @[Mux.scala 27:72]
  wire  _T_1612 = _T_2187 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1618 | _T_1612; // @[Mux.scala 27:72]
  wire  _T_1623 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 439:70]
  wire  ifu_byp_data_err_new = _T_1622 ? ic_miss_buff_data_error_bypass : _T_1623; // @[el2_ifu_mem_ctl.scala 437:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 382:42]
  wire  _T_2457 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 470:91]
  wire  _T_2458 = ~_T_2457; // @[el2_ifu_mem_ctl.scala 470:60]
  wire  ic_rd_parity_final_err = _T_2456 & _T_2458; // @[el2_ifu_mem_ctl.scala 470:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9985 = _T_4523 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 752:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9987 = _T_4527 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10240 = _T_9985 | _T_9987; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9989 = _T_4531 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10241 = _T_10240 | _T_9989; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9991 = _T_4535 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10242 = _T_10241 | _T_9991; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9993 = _T_4539 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10243 = _T_10242 | _T_9993; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9995 = _T_4543 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10244 = _T_10243 | _T_9995; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9997 = _T_4547 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10245 = _T_10244 | _T_9997; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9999 = _T_4551 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10246 = _T_10245 | _T_9999; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_10001 = _T_4555 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10247 = _T_10246 | _T_10001; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_10003 = _T_4559 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10248 = _T_10247 | _T_10003; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_10005 = _T_4563 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10249 = _T_10248 | _T_10005; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_10007 = _T_4567 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10250 = _T_10249 | _T_10007; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_10009 = _T_4571 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10251 = _T_10250 | _T_10009; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_10011 = _T_4575 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10252 = _T_10251 | _T_10011; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_10013 = _T_4579 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10253 = _T_10252 | _T_10013; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_10015 = _T_4583 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10254 = _T_10253 | _T_10015; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_10017 = _T_4587 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10255 = _T_10254 | _T_10017; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_10019 = _T_4591 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10256 = _T_10255 | _T_10019; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_10021 = _T_4595 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10257 = _T_10256 | _T_10021; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_10023 = _T_4599 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10258 = _T_10257 | _T_10023; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_10025 = _T_4603 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10259 = _T_10258 | _T_10025; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_10027 = _T_4607 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10260 = _T_10259 | _T_10027; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_10029 = _T_4611 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10261 = _T_10260 | _T_10029; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_10031 = _T_4615 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10262 = _T_10261 | _T_10031; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_10033 = _T_4619 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10263 = _T_10262 | _T_10033; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_10035 = _T_4623 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10264 = _T_10263 | _T_10035; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_10037 = _T_4627 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10265 = _T_10264 | _T_10037; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_10039 = _T_4631 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10266 = _T_10265 | _T_10039; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_10041 = _T_4635 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10267 = _T_10266 | _T_10041; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_10043 = _T_4639 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10268 = _T_10267 | _T_10043; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_10045 = _T_4643 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10269 = _T_10268 | _T_10045; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_10047 = _T_4647 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10270 = _T_10269 | _T_10047; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_10049 = _T_4651 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10271 = _T_10270 | _T_10049; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_10051 = _T_4655 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10272 = _T_10271 | _T_10051; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_10053 = _T_4659 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10273 = _T_10272 | _T_10053; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_10055 = _T_4663 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10274 = _T_10273 | _T_10055; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_10057 = _T_4667 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10275 = _T_10274 | _T_10057; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_10059 = _T_4671 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10276 = _T_10275 | _T_10059; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_10061 = _T_4675 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10277 = _T_10276 | _T_10061; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_10063 = _T_4679 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10278 = _T_10277 | _T_10063; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_10065 = _T_4683 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10279 = _T_10278 | _T_10065; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_10067 = _T_4687 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10280 = _T_10279 | _T_10067; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_10069 = _T_4691 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10281 = _T_10280 | _T_10069; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_10071 = _T_4695 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10282 = _T_10281 | _T_10071; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_10073 = _T_4699 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10283 = _T_10282 | _T_10073; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_10075 = _T_4703 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10284 = _T_10283 | _T_10075; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_10077 = _T_4707 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10285 = _T_10284 | _T_10077; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_10079 = _T_4711 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10286 = _T_10285 | _T_10079; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_10081 = _T_4715 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10287 = _T_10286 | _T_10081; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_10083 = _T_4719 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10288 = _T_10287 | _T_10083; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_10085 = _T_4723 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10289 = _T_10288 | _T_10085; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_10087 = _T_4727 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10290 = _T_10289 | _T_10087; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_10089 = _T_4731 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10291 = _T_10290 | _T_10089; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_10091 = _T_4735 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10292 = _T_10291 | _T_10091; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_10093 = _T_4739 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10293 = _T_10292 | _T_10093; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_10095 = _T_4743 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10294 = _T_10293 | _T_10095; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_10097 = _T_4747 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10295 = _T_10294 | _T_10097; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_10099 = _T_4751 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10296 = _T_10295 | _T_10099; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_10101 = _T_4755 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10297 = _T_10296 | _T_10101; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_10103 = _T_4759 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10298 = _T_10297 | _T_10103; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_10105 = _T_4763 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10299 = _T_10298 | _T_10105; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_10107 = _T_4767 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10300 = _T_10299 | _T_10107; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_10109 = _T_4771 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10301 = _T_10300 | _T_10109; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_10111 = _T_4775 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10302 = _T_10301 | _T_10111; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_10113 = _T_4779 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10303 = _T_10302 | _T_10113; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_10115 = _T_4783 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10304 = _T_10303 | _T_10115; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_10117 = _T_4787 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10305 = _T_10304 | _T_10117; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_10119 = _T_4791 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10306 = _T_10305 | _T_10119; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_10121 = _T_4795 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10307 = _T_10306 | _T_10121; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_10123 = _T_4799 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10308 = _T_10307 | _T_10123; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_10125 = _T_4803 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10309 = _T_10308 | _T_10125; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_10127 = _T_4807 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10310 = _T_10309 | _T_10127; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_10129 = _T_4811 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10311 = _T_10310 | _T_10129; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_10131 = _T_4815 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10312 = _T_10311 | _T_10131; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_10133 = _T_4819 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10313 = _T_10312 | _T_10133; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_10135 = _T_4823 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10314 = _T_10313 | _T_10135; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_10137 = _T_4827 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10315 = _T_10314 | _T_10137; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_10139 = _T_4831 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10316 = _T_10315 | _T_10139; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_10141 = _T_4835 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10317 = _T_10316 | _T_10141; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_10143 = _T_4839 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10318 = _T_10317 | _T_10143; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_10145 = _T_4843 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10319 = _T_10318 | _T_10145; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_10147 = _T_4847 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10320 = _T_10319 | _T_10147; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_10149 = _T_4851 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10321 = _T_10320 | _T_10149; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_10151 = _T_4855 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10322 = _T_10321 | _T_10151; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_10153 = _T_4859 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10323 = _T_10322 | _T_10153; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_10155 = _T_4863 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10324 = _T_10323 | _T_10155; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_10157 = _T_4867 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10325 = _T_10324 | _T_10157; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_10159 = _T_4871 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10326 = _T_10325 | _T_10159; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_10161 = _T_4875 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10327 = _T_10326 | _T_10161; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_10163 = _T_4879 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10328 = _T_10327 | _T_10163; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_10165 = _T_4883 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10329 = _T_10328 | _T_10165; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_10167 = _T_4887 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10330 = _T_10329 | _T_10167; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_10169 = _T_4891 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10331 = _T_10330 | _T_10169; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_10171 = _T_4895 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10332 = _T_10331 | _T_10171; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_10173 = _T_4899 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10333 = _T_10332 | _T_10173; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_10175 = _T_4903 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10334 = _T_10333 | _T_10175; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_10177 = _T_4907 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10335 = _T_10334 | _T_10177; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_10179 = _T_4911 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10336 = _T_10335 | _T_10179; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_10181 = _T_4915 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10337 = _T_10336 | _T_10181; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_10183 = _T_4919 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10338 = _T_10337 | _T_10183; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_10185 = _T_4923 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10339 = _T_10338 | _T_10185; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_10187 = _T_4927 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10340 = _T_10339 | _T_10187; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_10189 = _T_4931 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10341 = _T_10340 | _T_10189; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_10191 = _T_4935 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10342 = _T_10341 | _T_10191; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_10193 = _T_4939 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10343 = _T_10342 | _T_10193; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_10195 = _T_4943 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10344 = _T_10343 | _T_10195; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_10197 = _T_4947 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10345 = _T_10344 | _T_10197; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_10199 = _T_4951 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10346 = _T_10345 | _T_10199; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_10201 = _T_4955 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10347 = _T_10346 | _T_10201; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_10203 = _T_4959 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10348 = _T_10347 | _T_10203; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_10205 = _T_4963 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10349 = _T_10348 | _T_10205; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_10207 = _T_4967 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10350 = _T_10349 | _T_10207; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_10209 = _T_4971 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10351 = _T_10350 | _T_10209; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_10211 = _T_4975 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10352 = _T_10351 | _T_10211; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_10213 = _T_4979 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10353 = _T_10352 | _T_10213; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_10215 = _T_4983 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10354 = _T_10353 | _T_10215; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_10217 = _T_4987 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10355 = _T_10354 | _T_10217; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_10219 = _T_4991 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10356 = _T_10355 | _T_10219; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_10221 = _T_4995 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10357 = _T_10356 | _T_10221; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_10223 = _T_4999 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10358 = _T_10357 | _T_10223; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_10225 = _T_5003 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10359 = _T_10358 | _T_10225; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_10227 = _T_5007 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10360 = _T_10359 | _T_10227; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_10229 = _T_5011 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10361 = _T_10360 | _T_10229; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_10231 = _T_5015 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10362 = _T_10361 | _T_10231; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_10233 = _T_5019 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10363 = _T_10362 | _T_10233; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_10235 = _T_5023 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10364 = _T_10363 | _T_10235; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_10237 = _T_5027 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10365 = _T_10364 | _T_10237; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_10239 = _T_5031 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_10366 = _T_10365 | _T_10239; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9602 = _T_4523 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 752:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9604 = _T_4527 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9857 = _T_9602 | _T_9604; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9606 = _T_4531 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9858 = _T_9857 | _T_9606; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9608 = _T_4535 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9859 = _T_9858 | _T_9608; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9610 = _T_4539 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9860 = _T_9859 | _T_9610; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9612 = _T_4543 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9861 = _T_9860 | _T_9612; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9614 = _T_4547 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9862 = _T_9861 | _T_9614; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9616 = _T_4551 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9863 = _T_9862 | _T_9616; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9618 = _T_4555 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9864 = _T_9863 | _T_9618; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9620 = _T_4559 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9865 = _T_9864 | _T_9620; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9622 = _T_4563 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9866 = _T_9865 | _T_9622; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9624 = _T_4567 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9867 = _T_9866 | _T_9624; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9626 = _T_4571 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9868 = _T_9867 | _T_9626; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9628 = _T_4575 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9869 = _T_9868 | _T_9628; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9630 = _T_4579 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9870 = _T_9869 | _T_9630; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9632 = _T_4583 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9871 = _T_9870 | _T_9632; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9634 = _T_4587 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9872 = _T_9871 | _T_9634; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9636 = _T_4591 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9873 = _T_9872 | _T_9636; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9638 = _T_4595 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9874 = _T_9873 | _T_9638; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9640 = _T_4599 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9875 = _T_9874 | _T_9640; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9642 = _T_4603 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9876 = _T_9875 | _T_9642; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9644 = _T_4607 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9877 = _T_9876 | _T_9644; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9646 = _T_4611 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9878 = _T_9877 | _T_9646; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9648 = _T_4615 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9879 = _T_9878 | _T_9648; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9650 = _T_4619 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9880 = _T_9879 | _T_9650; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9652 = _T_4623 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9881 = _T_9880 | _T_9652; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9654 = _T_4627 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9882 = _T_9881 | _T_9654; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9656 = _T_4631 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9883 = _T_9882 | _T_9656; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9658 = _T_4635 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9884 = _T_9883 | _T_9658; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9660 = _T_4639 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9885 = _T_9884 | _T_9660; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9662 = _T_4643 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9886 = _T_9885 | _T_9662; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9664 = _T_4647 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9887 = _T_9886 | _T_9664; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9666 = _T_4651 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9888 = _T_9887 | _T_9666; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9668 = _T_4655 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9889 = _T_9888 | _T_9668; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9670 = _T_4659 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9890 = _T_9889 | _T_9670; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9672 = _T_4663 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9891 = _T_9890 | _T_9672; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9674 = _T_4667 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9892 = _T_9891 | _T_9674; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9676 = _T_4671 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9893 = _T_9892 | _T_9676; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9678 = _T_4675 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9894 = _T_9893 | _T_9678; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9680 = _T_4679 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9895 = _T_9894 | _T_9680; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9682 = _T_4683 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9896 = _T_9895 | _T_9682; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9684 = _T_4687 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9897 = _T_9896 | _T_9684; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9686 = _T_4691 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9898 = _T_9897 | _T_9686; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9688 = _T_4695 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9899 = _T_9898 | _T_9688; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9690 = _T_4699 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9900 = _T_9899 | _T_9690; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9692 = _T_4703 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9901 = _T_9900 | _T_9692; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9694 = _T_4707 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9902 = _T_9901 | _T_9694; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9696 = _T_4711 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9903 = _T_9902 | _T_9696; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9698 = _T_4715 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9904 = _T_9903 | _T_9698; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9700 = _T_4719 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9905 = _T_9904 | _T_9700; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9702 = _T_4723 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9906 = _T_9905 | _T_9702; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9704 = _T_4727 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9907 = _T_9906 | _T_9704; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9706 = _T_4731 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9908 = _T_9907 | _T_9706; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9708 = _T_4735 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9909 = _T_9908 | _T_9708; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9710 = _T_4739 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9910 = _T_9909 | _T_9710; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9712 = _T_4743 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9911 = _T_9910 | _T_9712; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9714 = _T_4747 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9912 = _T_9911 | _T_9714; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9716 = _T_4751 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9913 = _T_9912 | _T_9716; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9718 = _T_4755 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9914 = _T_9913 | _T_9718; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9720 = _T_4759 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9915 = _T_9914 | _T_9720; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9722 = _T_4763 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9916 = _T_9915 | _T_9722; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9724 = _T_4767 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9917 = _T_9916 | _T_9724; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9726 = _T_4771 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9918 = _T_9917 | _T_9726; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9728 = _T_4775 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9919 = _T_9918 | _T_9728; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9730 = _T_4779 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9920 = _T_9919 | _T_9730; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9732 = _T_4783 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9921 = _T_9920 | _T_9732; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9734 = _T_4787 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9922 = _T_9921 | _T_9734; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9736 = _T_4791 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9923 = _T_9922 | _T_9736; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9738 = _T_4795 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9924 = _T_9923 | _T_9738; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9740 = _T_4799 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9925 = _T_9924 | _T_9740; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9742 = _T_4803 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9926 = _T_9925 | _T_9742; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9744 = _T_4807 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9927 = _T_9926 | _T_9744; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9746 = _T_4811 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9928 = _T_9927 | _T_9746; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9748 = _T_4815 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9929 = _T_9928 | _T_9748; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9750 = _T_4819 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9930 = _T_9929 | _T_9750; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9752 = _T_4823 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9931 = _T_9930 | _T_9752; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9754 = _T_4827 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9932 = _T_9931 | _T_9754; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9756 = _T_4831 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9933 = _T_9932 | _T_9756; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9758 = _T_4835 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9934 = _T_9933 | _T_9758; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9760 = _T_4839 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9935 = _T_9934 | _T_9760; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9762 = _T_4843 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9936 = _T_9935 | _T_9762; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9764 = _T_4847 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9937 = _T_9936 | _T_9764; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9766 = _T_4851 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9938 = _T_9937 | _T_9766; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9768 = _T_4855 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9939 = _T_9938 | _T_9768; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9770 = _T_4859 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9940 = _T_9939 | _T_9770; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9772 = _T_4863 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9941 = _T_9940 | _T_9772; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9774 = _T_4867 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9942 = _T_9941 | _T_9774; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9776 = _T_4871 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9943 = _T_9942 | _T_9776; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9778 = _T_4875 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9944 = _T_9943 | _T_9778; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9780 = _T_4879 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9945 = _T_9944 | _T_9780; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9782 = _T_4883 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9946 = _T_9945 | _T_9782; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9784 = _T_4887 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9947 = _T_9946 | _T_9784; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9786 = _T_4891 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9948 = _T_9947 | _T_9786; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9788 = _T_4895 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9949 = _T_9948 | _T_9788; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9790 = _T_4899 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9950 = _T_9949 | _T_9790; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9792 = _T_4903 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9951 = _T_9950 | _T_9792; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9794 = _T_4907 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9952 = _T_9951 | _T_9794; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9796 = _T_4911 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9953 = _T_9952 | _T_9796; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9798 = _T_4915 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9954 = _T_9953 | _T_9798; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9800 = _T_4919 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9955 = _T_9954 | _T_9800; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9802 = _T_4923 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9956 = _T_9955 | _T_9802; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9804 = _T_4927 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9957 = _T_9956 | _T_9804; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9806 = _T_4931 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9958 = _T_9957 | _T_9806; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9808 = _T_4935 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9959 = _T_9958 | _T_9808; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9810 = _T_4939 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9960 = _T_9959 | _T_9810; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9812 = _T_4943 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9961 = _T_9960 | _T_9812; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9814 = _T_4947 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9962 = _T_9961 | _T_9814; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9816 = _T_4951 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9963 = _T_9962 | _T_9816; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9818 = _T_4955 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9964 = _T_9963 | _T_9818; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9820 = _T_4959 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9965 = _T_9964 | _T_9820; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9822 = _T_4963 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9966 = _T_9965 | _T_9822; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9824 = _T_4967 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9967 = _T_9966 | _T_9824; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9826 = _T_4971 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9968 = _T_9967 | _T_9826; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9828 = _T_4975 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9969 = _T_9968 | _T_9828; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9830 = _T_4979 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9970 = _T_9969 | _T_9830; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9832 = _T_4983 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9971 = _T_9970 | _T_9832; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9834 = _T_4987 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9972 = _T_9971 | _T_9834; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9836 = _T_4991 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9973 = _T_9972 | _T_9836; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9838 = _T_4995 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9974 = _T_9973 | _T_9838; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9840 = _T_4999 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9975 = _T_9974 | _T_9840; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9842 = _T_5003 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9976 = _T_9975 | _T_9842; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9844 = _T_5007 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9977 = _T_9976 | _T_9844; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9846 = _T_5011 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9978 = _T_9977 | _T_9846; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9848 = _T_5015 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9979 = _T_9978 | _T_9848; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9850 = _T_5019 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9980 = _T_9979 | _T_9850; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9852 = _T_5023 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9981 = _T_9980 | _T_9852; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9854 = _T_5027 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9982 = _T_9981 | _T_9854; // @[el2_ifu_mem_ctl.scala 752:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9856 = _T_5031 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 752:10]
  wire  _T_9983 = _T_9982 | _T_9856; // @[el2_ifu_mem_ctl.scala 752:91]
  wire [1:0] ic_tag_valid_unq = {_T_10366,_T_9983}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 826:54]
  wire [1:0] _T_10406 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10407 = ic_debug_way_ff & _T_10406; // @[el2_ifu_mem_ctl.scala 807:67]
  wire [1:0] _T_10408 = ic_tag_valid_unq & _T_10407; // @[el2_ifu_mem_ctl.scala 807:48]
  wire  ic_debug_tag_val_rd_out = |_T_10408; // @[el2_ifu_mem_ctl.scala 807:115]
  wire [65:0] _T_1208 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1209; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2591; // @[el2_ifu_mem_ctl.scala 365:80]
  wire  _T_1247 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 370:98]
  wire  sel_byp_data = _T_1251 & _T_1247; // @[el2_ifu_mem_ctl.scala 370:96]
  wire [63:0] _T_1258 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1259 = _T_1258 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 377:64]
  wire [63:0] _T_1261 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2113 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 445:31]
  wire  _T_1626 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 441:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1627 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1675 = _T_1627 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1630 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1676 = _T_1630 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1675 | _T_1676; // @[Mux.scala 27:72]
  wire  _T_1633 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1677 = _T_1633 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1692 = _T_1691 | _T_1677; // @[Mux.scala 27:72]
  wire  _T_1636 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1678 = _T_1636 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1692 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1639 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1679 = _T_1639 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire  _T_1642 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1680 = _T_1642 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1695 = _T_1694 | _T_1680; // @[Mux.scala 27:72]
  wire  _T_1645 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1681 = _T_1645 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1696 = _T_1695 | _T_1681; // @[Mux.scala 27:72]
  wire  _T_1648 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1682 = _T_1648 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1697 = _T_1696 | _T_1682; // @[Mux.scala 27:72]
  wire  _T_1651 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1683 = _T_1651 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1698 = _T_1697 | _T_1683; // @[Mux.scala 27:72]
  wire  _T_1654 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1684 = _T_1654 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1699 = _T_1698 | _T_1684; // @[Mux.scala 27:72]
  wire  _T_1657 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1685 = _T_1657 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1700 = _T_1699 | _T_1685; // @[Mux.scala 27:72]
  wire  _T_1660 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1686 = _T_1660 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1701 = _T_1700 | _T_1686; // @[Mux.scala 27:72]
  wire  _T_1663 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1687 = _T_1663 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1702 = _T_1701 | _T_1687; // @[Mux.scala 27:72]
  wire  _T_1666 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1688 = _T_1666 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1703 = _T_1702 | _T_1688; // @[Mux.scala 27:72]
  wire  _T_1669 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1689 = _T_1669 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1704 = _T_1703 | _T_1689; // @[Mux.scala 27:72]
  wire  _T_1672 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1690 = _T_1672 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1705 = _T_1704 | _T_1690; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1707 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1755 = _T_1707 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1710 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1756 = _T_1710 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1755 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1713 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1757 = _T_1713 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1772 = _T_1771 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1716 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1758 = _T_1716 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1772 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1719 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1759 = _T_1719 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1722 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1760 = _T_1722 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1775 = _T_1774 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1725 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1761 = _T_1725 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1776 = _T_1775 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1728 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1762 = _T_1728 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1777 = _T_1776 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1731 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1763 = _T_1731 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1778 = _T_1777 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1734 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1764 = _T_1734 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1779 = _T_1778 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1737 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1765 = _T_1737 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1780 = _T_1779 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1740 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1766 = _T_1740 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1781 = _T_1780 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1743 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1767 = _T_1743 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1782 = _T_1781 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1746 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1768 = _T_1746 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1783 = _T_1782 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1749 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1769 = _T_1749 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1784 = _T_1783 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1752 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1770 = _T_1752 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1785 = _T_1784 | _T_1770; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1787 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1835 = _T_1787 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1790 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1836 = _T_1790 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1835 | _T_1836; // @[Mux.scala 27:72]
  wire  _T_1793 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1837 = _T_1793 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1852 = _T_1851 | _T_1837; // @[Mux.scala 27:72]
  wire  _T_1796 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1838 = _T_1796 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1852 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1799 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1839 = _T_1799 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire  _T_1802 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1840 = _T_1802 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1855 = _T_1854 | _T_1840; // @[Mux.scala 27:72]
  wire  _T_1805 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1841 = _T_1805 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1856 = _T_1855 | _T_1841; // @[Mux.scala 27:72]
  wire  _T_1808 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1842 = _T_1808 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1857 = _T_1856 | _T_1842; // @[Mux.scala 27:72]
  wire  _T_1811 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1843 = _T_1811 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1858 = _T_1857 | _T_1843; // @[Mux.scala 27:72]
  wire  _T_1814 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1844 = _T_1814 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1859 = _T_1858 | _T_1844; // @[Mux.scala 27:72]
  wire  _T_1817 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1845 = _T_1817 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1860 = _T_1859 | _T_1845; // @[Mux.scala 27:72]
  wire  _T_1820 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1846 = _T_1820 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1861 = _T_1860 | _T_1846; // @[Mux.scala 27:72]
  wire  _T_1823 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1847 = _T_1823 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1862 = _T_1861 | _T_1847; // @[Mux.scala 27:72]
  wire  _T_1826 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1848 = _T_1826 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1863 = _T_1862 | _T_1848; // @[Mux.scala 27:72]
  wire  _T_1829 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1849 = _T_1829 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1864 = _T_1863 | _T_1849; // @[Mux.scala 27:72]
  wire  _T_1832 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1850 = _T_1832 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1865 = _T_1864 | _T_1850; // @[Mux.scala 27:72]
  wire [79:0] _T_1868 = {_T_1705,_T_1785,_T_1865}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1869 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1917 = _T_1869 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1918 = _T_1872 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1917 | _T_1918; // @[Mux.scala 27:72]
  wire  _T_1875 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1919 = _T_1875 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1934 = _T_1933 | _T_1919; // @[Mux.scala 27:72]
  wire  _T_1878 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1920 = _T_1878 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1934 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1881 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1921 = _T_1881 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire  _T_1884 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1922 = _T_1884 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1937 = _T_1936 | _T_1922; // @[Mux.scala 27:72]
  wire  _T_1887 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1923 = _T_1887 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1938 = _T_1937 | _T_1923; // @[Mux.scala 27:72]
  wire  _T_1890 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1924 = _T_1890 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1939 = _T_1938 | _T_1924; // @[Mux.scala 27:72]
  wire  _T_1893 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1925 = _T_1893 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1940 = _T_1939 | _T_1925; // @[Mux.scala 27:72]
  wire  _T_1896 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1926 = _T_1896 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1941 = _T_1940 | _T_1926; // @[Mux.scala 27:72]
  wire  _T_1899 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1927 = _T_1899 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1942 = _T_1941 | _T_1927; // @[Mux.scala 27:72]
  wire  _T_1902 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1928 = _T_1902 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1943 = _T_1942 | _T_1928; // @[Mux.scala 27:72]
  wire  _T_1905 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1929 = _T_1905 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1944 = _T_1943 | _T_1929; // @[Mux.scala 27:72]
  wire  _T_1908 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1930 = _T_1908 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1945 = _T_1944 | _T_1930; // @[Mux.scala 27:72]
  wire  _T_1911 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1931 = _T_1911 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1946 = _T_1945 | _T_1931; // @[Mux.scala 27:72]
  wire  _T_1914 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1932 = _T_1914 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1947 = _T_1946 | _T_1932; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1627 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1630 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_1997 | _T_1998; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1633 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_2013 | _T_1999; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1636 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_2014 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1639 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1642 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2017 = _T_2016 | _T_2002; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_1645 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2018 = _T_2017 | _T_2003; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_1648 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2019 = _T_2018 | _T_2004; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_1651 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2020 = _T_2019 | _T_2005; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_1654 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2021 = _T_2020 | _T_2006; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_1657 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2022 = _T_2021 | _T_2007; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_1660 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2023 = _T_2022 | _T_2008; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_1663 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2024 = _T_2023 | _T_2009; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_1666 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2025 = _T_2024 | _T_2010; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_1669 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2026 = _T_2025 | _T_2011; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_1672 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2027 = _T_2026 | _T_2012; // @[Mux.scala 27:72]
  wire [79:0] _T_2110 = {_T_1947,_T_2027,_T_1785}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1626 ? _T_1868 : _T_2110; // @[el2_ifu_mem_ctl.scala 441:37]
  wire [79:0] _T_2115 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2113 ? ic_byp_data_only_pre_new : _T_2115; // @[el2_ifu_mem_ctl.scala 445:30]
  wire [79:0] _GEN_794 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 377:109]
  wire [79:0] _T_1262 = _GEN_794 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 377:109]
  wire [79:0] _GEN_795 = {{16'd0}, _T_1259}; // @[el2_ifu_mem_ctl.scala 377:83]
  wire [79:0] ic_premux_data = _GEN_795 | _T_1262; // @[el2_ifu_mem_ctl.scala 377:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 384:38]
  wire [1:0] _T_1271 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 388:8]
  wire  _T_1273 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 390:45]
  wire  _T_1275 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 390:80]
  wire  _T_1276 = ~_T_1275; // @[el2_ifu_mem_ctl.scala 390:71]
  wire  _T_1277 = _T_1273 & _T_1276; // @[el2_ifu_mem_ctl.scala 390:69]
  wire  _T_1278 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 390:131]
  wire  _T_1279 = _T_1277 & _T_1278; // @[el2_ifu_mem_ctl.scala 390:114]
  wire [7:0] _T_1368 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1373 = ic_miss_buff_data_error[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  _T_2659 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 621:47]
  wire  _T_2660 = _T_2659 & _T_13; // @[el2_ifu_mem_ctl.scala 621:50]
  wire  bus_ifu_wr_data_error = _T_2660 & miss_pending; // @[el2_ifu_mem_ctl.scala 621:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1373; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1377 = ic_miss_buff_data_error[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1377; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1381 = ic_miss_buff_data_error[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1381; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1385 = ic_miss_buff_data_error[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1385; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1389 = ic_miss_buff_data_error[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1389; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1393 = ic_miss_buff_data_error[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1393; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1397 = ic_miss_buff_data_error[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1397; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1401 = ic_miss_buff_data_error[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1401; // @[el2_ifu_mem_ctl.scala 407:72]
  wire [7:0] _T_1408 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2465 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2473 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 490:65]
  wire  _T_2474 = _T_2473 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 490:88]
  wire  _T_2476 = _T_2474 & _T_2587; // @[el2_ifu_mem_ctl.scala 490:112]
  wire  _T_2477 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2478 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 495:50]
  wire  _T_2480 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2486 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2488 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_2486 | _T_2488; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2480 ? _T_2478 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_2477 ? _T_2478 : _GEN_41; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2465 ? _T_2476 : _GEN_43; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2465 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2479 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 496:56]
  wire  _GEN_44 = _T_2477 & _T_2479; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2465 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 481:58]
  wire  _T_2462 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 480:49]
  wire  _T_2467 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 489:87]
  wire  _T_2481 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 499:54]
  wire  _T_2482 = _T_2481 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 499:84]
  wire  _T_2491 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 520:66]
  wire  _T_2492 = io_dec_tlu_flush_err_wb & _T_2491; // @[el2_ifu_mem_ctl.scala 520:52]
  wire  _T_2494 = _T_2492 & _T_2587; // @[el2_ifu_mem_ctl.scala 520:81]
  wire  _T_2496 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 523:59]
  wire  _T_2497 = _T_2496 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 523:86]
  wire  _T_2511 = _T_2496 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 526:81]
  wire  _T_2512 = _T_2511 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 526:103]
  wire  _T_2513 = _T_2512 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 526:126]
  wire  _T_2533 = _T_2511 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 533:103]
  wire  _T_2540 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 538:62]
  wire  _T_2541 = io_dec_tlu_flush_lower_wb & _T_2540; // @[el2_ifu_mem_ctl.scala 538:60]
  wire  _T_2542 = _T_2541 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 538:88]
  wire  _T_2543 = _T_2542 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 538:115]
  wire  _GEN_51 = _T_2539 & _T_2497; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_2522 ? _T_2533 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_2522 | _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2495 ? _T_2513 : _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_2495 | _GEN_56; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2490 ? _T_2494 : _GEN_58; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2555 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 555:64]
  wire  _T_2557 = _T_2555 & _T_2587; // @[el2_ifu_mem_ctl.scala 555:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2559 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 555:133]
  wire  _T_2560 = _T_2559 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 555:164]
  wire  _T_2561 = _T_2560 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 555:184]
  wire  _T_2562 = _T_2561 & miss_pending; // @[el2_ifu_mem_ctl.scala 555:204]
  wire  _T_2563 = ~_T_2562; // @[el2_ifu_mem_ctl.scala 555:112]
  wire  ifc_bus_ic_req_ff_in = _T_2557 & _T_2563; // @[el2_ifu_mem_ctl.scala 555:110]
  wire  _T_2564 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 556:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 587:45]
  wire  _T_2581 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 590:35]
  wire  _T_2582 = _T_2581 & miss_pending; // @[el2_ifu_mem_ctl.scala 590:53]
  wire  bus_cmd_sent = _T_2582 & _T_2587; // @[el2_ifu_mem_ctl.scala 590:68]
  wire [2:0] _T_2572 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2574 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2576 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 588:51]
  wire  _T_2602 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 598:73]
  wire  _T_2603 = _T_2588 & _T_2602; // @[el2_ifu_mem_ctl.scala 598:71]
  wire  _T_2605 = last_data_recieved_ff & _T_1339; // @[el2_ifu_mem_ctl.scala 598:114]
  wire  last_data_recieved_in = _T_2603 | _T_2605; // @[el2_ifu_mem_ctl.scala 598:89]
  wire [2:0] _T_2611 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 603:45]
  wire  _T_2614 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 604:81]
  wire  _T_2615 = _T_2614 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 604:97]
  wire  _T_2617 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 606:48]
  wire  _T_2618 = _T_2617 & miss_pending; // @[el2_ifu_mem_ctl.scala 606:68]
  wire  bus_inc_cmd_beat_cnt = _T_2618 & _T_2587; // @[el2_ifu_mem_ctl.scala 606:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 608:57]
  wire  _T_2622 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 609:31]
  wire  _T_2623 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 609:71]
  wire  _T_2624 = _T_2623 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 609:87]
  wire  _T_2625 = ~_T_2624; // @[el2_ifu_mem_ctl.scala 609:55]
  wire  bus_hold_cmd_beat_cnt = _T_2622 & _T_2625; // @[el2_ifu_mem_ctl.scala 609:53]
  wire  _T_2626 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 610:46]
  wire  bus_cmd_beat_en = _T_2626 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 610:62]
  wire [2:0] _T_2629 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 612:46]
  wire [2:0] _T_2631 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2632 = bus_inc_cmd_beat_cnt ? _T_2629 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2633 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2635 = _T_2631 | _T_2632; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2635 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2639 = _T_2615 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 613:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 624:62]
  wire  _T_2667 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 629:50]
  wire  _T_2668 = io_ifc_dma_access_ok & _T_2667; // @[el2_ifu_mem_ctl.scala 629:47]
  wire  _T_2669 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 629:70]
  wire  ifc_dma_access_ok_d = _T_2668 & _T_2669; // @[el2_ifu_mem_ctl.scala 629:68]
  wire  _T_2673 = _T_2668 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 630:72]
  wire  _T_2674 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 630:111]
  wire  _T_2675 = _T_2673 & _T_2674; // @[el2_ifu_mem_ctl.scala 630:97]
  wire  ifc_dma_access_q_ok = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 630:127]
  wire  _T_2678 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 633:40]
  wire  _T_2679 = _T_2678 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 633:58]
  wire  _T_2682 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 634:60]
  wire  _T_2683 = _T_2678 & _T_2682; // @[el2_ifu_mem_ctl.scala 634:58]
  wire  _T_2684 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 634:104]
  wire [2:0] _T_2689 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2795 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2804 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2795}; // @[el2_lib.scala 268:22]
  wire  _T_2805 = ^_T_2804; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2813 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2822 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2813}; // @[el2_lib.scala 268:39]
  wire  _T_2823 = ^_T_2822; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2831 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2840 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2831}; // @[el2_lib.scala 268:56]
  wire  _T_2841 = ^_T_2840; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2847 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2855 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2847}; // @[el2_lib.scala 268:73]
  wire  _T_2856 = ^_T_2855; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2870 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2847}; // @[el2_lib.scala 268:90]
  wire  _T_2871 = ^_T_2870; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2876 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2877 = ^_T_2876; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2882 = {_T_2805,_T_2823,_T_2841,_T_2856,_T_2871,_T_2877}; // @[Cat.scala 29:58]
  wire  _T_2883 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2884 = ^_T_2882; // @[el2_lib.scala 269:23]
  wire  _T_2885 = _T_2883 ^ _T_2884; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2991 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_3000 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2991}; // @[el2_lib.scala 268:22]
  wire  _T_3001 = ^_T_3000; // @[el2_lib.scala 268:29]
  wire [8:0] _T_3009 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_3018 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_3009}; // @[el2_lib.scala 268:39]
  wire  _T_3019 = ^_T_3018; // @[el2_lib.scala 268:46]
  wire [8:0] _T_3027 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_3036 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_3027}; // @[el2_lib.scala 268:56]
  wire  _T_3037 = ^_T_3036; // @[el2_lib.scala 268:63]
  wire [6:0] _T_3043 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_3051 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_3043}; // @[el2_lib.scala 268:73]
  wire  _T_3052 = ^_T_3051; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3066 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_3043}; // @[el2_lib.scala 268:90]
  wire  _T_3067 = ^_T_3066; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3072 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3073 = ^_T_3072; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3078 = {_T_3001,_T_3019,_T_3037,_T_3052,_T_3067,_T_3073}; // @[Cat.scala 29:58]
  wire  _T_3079 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3080 = ^_T_3078; // @[el2_lib.scala 269:23]
  wire  _T_3081 = _T_3079 ^ _T_3080; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3082 = {_T_3081,_T_3001,_T_3019,_T_3037,_T_3052,_T_3067,_T_3073}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2885,_T_2805,_T_2823,_T_2841,_T_2856,_T_2871,_T_2877,_T_3082}; // @[Cat.scala 29:58]
  wire  _T_3084 = ~_T_2678; // @[el2_ifu_mem_ctl.scala 639:45]
  wire  _T_3085 = iccm_correct_ecc & _T_3084; // @[el2_ifu_mem_ctl.scala 639:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3086 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3093 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 653:53]
  wire  _T_3425 = _T_3337[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3423 = _T_3337[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3421 = _T_3337[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3419 = _T_3337[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3417 = _T_3337[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3415 = _T_3337[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3413 = _T_3337[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3411 = _T_3337[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3409 = _T_3337[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3407 = _T_3337[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3483 = {_T_3425,_T_3423,_T_3421,_T_3419,_T_3417,_T_3415,_T_3413,_T_3411,_T_3409,_T_3407}; // @[el2_lib.scala 310:69]
  wire  _T_3405 = _T_3337[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3403 = _T_3337[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3401 = _T_3337[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3399 = _T_3337[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3397 = _T_3337[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3395 = _T_3337[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3393 = _T_3337[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3391 = _T_3337[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3389 = _T_3337[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3387 = _T_3337[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3474 = {_T_3405,_T_3403,_T_3401,_T_3399,_T_3397,_T_3395,_T_3393,_T_3391,_T_3389,_T_3387}; // @[el2_lib.scala 310:69]
  wire  _T_3385 = _T_3337[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3383 = _T_3337[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3381 = _T_3337[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3379 = _T_3337[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3377 = _T_3337[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3375 = _T_3337[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3373 = _T_3337[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3371 = _T_3337[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3369 = _T_3337[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3367 = _T_3337[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3464 = {_T_3385,_T_3383,_T_3381,_T_3379,_T_3377,_T_3375,_T_3373,_T_3371,_T_3369,_T_3367}; // @[el2_lib.scala 310:69]
  wire  _T_3365 = _T_3337[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3363 = _T_3337[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3361 = _T_3337[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3359 = _T_3337[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3357 = _T_3337[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3355 = _T_3337[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3353 = _T_3337[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3351 = _T_3337[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3349 = _T_3337[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3465 = {_T_3464,_T_3365,_T_3363,_T_3361,_T_3359,_T_3357,_T_3355,_T_3353,_T_3351,_T_3349}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3485 = {_T_3483,_T_3474,_T_3465}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3440 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3446 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3440}; // @[Cat.scala 29:58]
  wire [38:0] _T_3486 = _T_3485 ^ _T_3446; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3487 = _T_3341 ? _T_3486 : _T_3446; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3487[37:32],_T_3487[30:16],_T_3487[14:8],_T_3487[6:4],_T_3487[2]}; // @[Cat.scala 29:58]
  wire  _T_3810 = _T_3722[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3808 = _T_3722[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3806 = _T_3722[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3804 = _T_3722[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3802 = _T_3722[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3800 = _T_3722[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3798 = _T_3722[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3796 = _T_3722[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3794 = _T_3722[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3792 = _T_3722[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3868 = {_T_3810,_T_3808,_T_3806,_T_3804,_T_3802,_T_3800,_T_3798,_T_3796,_T_3794,_T_3792}; // @[el2_lib.scala 310:69]
  wire  _T_3790 = _T_3722[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3788 = _T_3722[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3786 = _T_3722[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3784 = _T_3722[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3782 = _T_3722[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3780 = _T_3722[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3778 = _T_3722[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3776 = _T_3722[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3774 = _T_3722[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3772 = _T_3722[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3859 = {_T_3790,_T_3788,_T_3786,_T_3784,_T_3782,_T_3780,_T_3778,_T_3776,_T_3774,_T_3772}; // @[el2_lib.scala 310:69]
  wire  _T_3770 = _T_3722[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3768 = _T_3722[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3766 = _T_3722[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3764 = _T_3722[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3762 = _T_3722[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3760 = _T_3722[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3758 = _T_3722[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3756 = _T_3722[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3754 = _T_3722[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3752 = _T_3722[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3849 = {_T_3770,_T_3768,_T_3766,_T_3764,_T_3762,_T_3760,_T_3758,_T_3756,_T_3754,_T_3752}; // @[el2_lib.scala 310:69]
  wire  _T_3750 = _T_3722[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3748 = _T_3722[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3746 = _T_3722[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3744 = _T_3722[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3742 = _T_3722[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3740 = _T_3722[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3738 = _T_3722[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3736 = _T_3722[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3734 = _T_3722[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3850 = {_T_3849,_T_3750,_T_3748,_T_3746,_T_3744,_T_3742,_T_3740,_T_3738,_T_3736,_T_3734}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3870 = {_T_3868,_T_3859,_T_3850}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3825 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3831 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3825}; // @[Cat.scala 29:58]
  wire [38:0] _T_3871 = _T_3870 ^ _T_3831; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3872 = _T_3726 ? _T_3871 : _T_3831; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3872[37:32],_T_3872[30:16],_T_3872[14:8],_T_3872[6:4],_T_3872[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 645:35]
  wire  _T_3345 = ~_T_3337[6]; // @[el2_lib.scala 303:55]
  wire  _T_3346 = _T_3339 & _T_3345; // @[el2_lib.scala 303:53]
  wire  _T_3730 = ~_T_3722[6]; // @[el2_lib.scala 303:55]
  wire  _T_3731 = _T_3724 & _T_3730; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3346,_T_3731}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 647:53]
  wire [63:0] _T_3097 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3098 = {iccm_dma_rdata_1_muxed,_T_3487[37:32],_T_3487[30:16],_T_3487[14:8],_T_3487[6:4],_T_3487[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 649:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 650:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 655:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 659:70]
  wire  _T_3103 = _T_2678 & _T_2667; // @[el2_ifu_mem_ctl.scala 662:65]
  wire  _T_3106 = _T_3084 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 663:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3107 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3109 = _T_3106 ? {{1'd0}, _T_3107} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 663:8]
  wire [31:0] _T_3110 = _T_3103 ? io_dma_mem_addr : {{16'd0}, _T_3109}; // @[el2_ifu_mem_ctl.scala 662:25]
  wire  _T_3499 = _T_3337 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3500 = _T_3487[38] ^ _T_3499; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3500,_T_3487[31],_T_3487[15],_T_3487[7],_T_3487[3],_T_3487[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3884 = _T_3722 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3885 = _T_3872[38] ^ _T_3884; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3885,_T_3872[31],_T_3872[15],_T_3872[7],_T_3872[3],_T_3872[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3901 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 675:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 677:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 678:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 686:62]
  wire  _T_3909 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 680:76]
  wire  _T_3910 = io_iccm_rd_ecc_single_err & _T_3909; // @[el2_ifu_mem_ctl.scala 680:74]
  wire  _T_3912 = _T_3910 & _T_317; // @[el2_ifu_mem_ctl.scala 680:104]
  wire  iccm_ecc_write_status = _T_3912 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 680:127]
  wire  _T_3913 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 681:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3913 & _T_317; // @[el2_ifu_mem_ctl.scala 681:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 685:51]
  wire [13:0] _T_3918 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 684:102]
  wire [38:0] _T_3922 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3927 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 689:41]
  wire  _T_3928 = io_ifc_fetch_req_bf & _T_3927; // @[el2_ifu_mem_ctl.scala 689:39]
  wire  _T_3929 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 689:72]
  wire  _T_3930 = _T_3928 & _T_3929; // @[el2_ifu_mem_ctl.scala 689:70]
  wire  _T_3932 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 690:34]
  wire  _T_3933 = _T_2233 & _T_3932; // @[el2_ifu_mem_ctl.scala 690:32]
  wire  _T_3936 = _T_2249 & _T_3932; // @[el2_ifu_mem_ctl.scala 691:37]
  wire  _T_3937 = _T_3933 | _T_3936; // @[el2_ifu_mem_ctl.scala 690:88]
  wire  _T_3938 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 692:19]
  wire  _T_3940 = _T_3938 & _T_3932; // @[el2_ifu_mem_ctl.scala 692:41]
  wire  _T_3941 = _T_3937 | _T_3940; // @[el2_ifu_mem_ctl.scala 691:88]
  wire  _T_3942 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 693:19]
  wire  _T_3944 = _T_3942 & _T_3932; // @[el2_ifu_mem_ctl.scala 693:35]
  wire  _T_3945 = _T_3941 | _T_3944; // @[el2_ifu_mem_ctl.scala 692:88]
  wire  _T_3948 = _T_2248 & _T_3932; // @[el2_ifu_mem_ctl.scala 694:38]
  wire  _T_3949 = _T_3945 | _T_3948; // @[el2_ifu_mem_ctl.scala 693:88]
  wire  _T_3951 = _T_2249 & miss_state_en; // @[el2_ifu_mem_ctl.scala 695:37]
  wire  _T_3952 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 695:71]
  wire  _T_3953 = _T_3951 & _T_3952; // @[el2_ifu_mem_ctl.scala 695:54]
  wire  _T_3954 = _T_3949 | _T_3953; // @[el2_ifu_mem_ctl.scala 694:57]
  wire  _T_3955 = ~_T_3954; // @[el2_ifu_mem_ctl.scala 690:5]
  wire  _T_3956 = _T_3930 & _T_3955; // @[el2_ifu_mem_ctl.scala 689:96]
  wire  _T_3957 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 696:28]
  wire  _T_3959 = _T_3957 & _T_3927; // @[el2_ifu_mem_ctl.scala 696:50]
  wire  _T_3961 = _T_3959 & _T_3929; // @[el2_ifu_mem_ctl.scala 696:81]
  wire [1:0] _T_3964 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10391 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 784:74]
  wire  bus_wren_1 = _T_10391 & miss_pending; // @[el2_ifu_mem_ctl.scala 784:98]
  wire  _T_10390 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 784:74]
  wire  bus_wren_0 = _T_10390 & miss_pending; // @[el2_ifu_mem_ctl.scala 784:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3970 = ~_T_108; // @[el2_ifu_mem_ctl.scala 699:106]
  wire  _T_3971 = _T_2233 & _T_3970; // @[el2_ifu_mem_ctl.scala 699:104]
  wire  _T_3972 = _T_2249 | _T_3971; // @[el2_ifu_mem_ctl.scala 699:77]
  wire  _T_3976 = ~_T_51; // @[el2_ifu_mem_ctl.scala 699:172]
  wire  _T_3977 = _T_3972 & _T_3976; // @[el2_ifu_mem_ctl.scala 699:170]
  wire  _T_3978 = ~_T_3977; // @[el2_ifu_mem_ctl.scala 699:44]
  wire  _T_3982 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 702:64]
  wire  _T_3983 = ~_T_3982; // @[el2_ifu_mem_ctl.scala 702:50]
  wire  _T_3984 = _T_276 & _T_3983; // @[el2_ifu_mem_ctl.scala 702:48]
  wire  _T_3985 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 702:81]
  wire  ic_valid = _T_3984 & _T_3985; // @[el2_ifu_mem_ctl.scala 702:79]
  wire  _T_3987 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 703:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 706:14]
  wire  _T_3990 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 709:74]
  wire  _T_10388 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 783:45]
  wire  way_status_wr_en = _T_10388 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 783:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3990; // @[el2_ifu_mem_ctl.scala 709:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:14]
  wire [2:0] _T_3994 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 715:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 779:41]
  wire  way_status_new = _T_10388 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 782:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 717:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 719:132]
  wire  _T_4011 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4012 = _T_4011 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4013 = _T_4012 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4015 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4016 = _T_4015 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4017 = _T_4016 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4019 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4020 = _T_4019 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4021 = _T_4020 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4023 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4024 = _T_4023 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4025 = _T_4024 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4027 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4028 = _T_4027 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4029 = _T_4028 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4031 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4032 = _T_4031 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4033 = _T_4032 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4035 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4036 = _T_4035 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4037 = _T_4036 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4039 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 723:93]
  wire  _T_4040 = _T_4039 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 723:102]
  wire  _T_4041 = _T_4040 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4045 = _T_4012 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4049 = _T_4016 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4053 = _T_4020 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4057 = _T_4024 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4061 = _T_4028 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4065 = _T_4032 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4069 = _T_4036 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4073 = _T_4040 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4077 = _T_4012 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4081 = _T_4016 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4085 = _T_4020 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4089 = _T_4024 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4093 = _T_4028 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4097 = _T_4032 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4101 = _T_4036 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4105 = _T_4040 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4109 = _T_4012 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4113 = _T_4016 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4117 = _T_4020 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4121 = _T_4024 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4125 = _T_4028 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4129 = _T_4032 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4133 = _T_4036 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4137 = _T_4040 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4141 = _T_4012 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4145 = _T_4016 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4149 = _T_4020 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4153 = _T_4024 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4157 = _T_4028 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4161 = _T_4032 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4165 = _T_4036 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4169 = _T_4040 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4173 = _T_4012 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4177 = _T_4016 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4181 = _T_4020 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4185 = _T_4024 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4189 = _T_4028 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4193 = _T_4032 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4197 = _T_4036 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4201 = _T_4040 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4205 = _T_4012 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4209 = _T_4016 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4213 = _T_4020 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4217 = _T_4024 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4221 = _T_4028 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4225 = _T_4032 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4229 = _T_4036 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4233 = _T_4040 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4237 = _T_4012 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4241 = _T_4016 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4245 = _T_4020 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4249 = _T_4024 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4253 = _T_4028 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4257 = _T_4032 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4261 = _T_4036 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4265 = _T_4040 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4269 = _T_4012 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4273 = _T_4016 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4277 = _T_4020 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4281 = _T_4024 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4285 = _T_4028 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4289 = _T_4032 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4293 = _T_4036 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4297 = _T_4040 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4301 = _T_4012 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4305 = _T_4016 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4309 = _T_4020 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4313 = _T_4024 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4317 = _T_4028 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4321 = _T_4032 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4325 = _T_4036 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4329 = _T_4040 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4333 = _T_4012 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4337 = _T_4016 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4341 = _T_4020 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4345 = _T_4024 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4349 = _T_4028 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4353 = _T_4032 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4357 = _T_4036 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4361 = _T_4040 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4365 = _T_4012 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4369 = _T_4016 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4373 = _T_4020 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4377 = _T_4024 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4381 = _T_4028 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4385 = _T_4032 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4389 = _T_4036 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4393 = _T_4040 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4397 = _T_4012 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4401 = _T_4016 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4405 = _T_4020 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4409 = _T_4024 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4413 = _T_4028 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4417 = _T_4032 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4421 = _T_4036 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4425 = _T_4040 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4429 = _T_4012 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4433 = _T_4016 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4437 = _T_4020 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4441 = _T_4024 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4445 = _T_4028 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4449 = _T_4032 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4453 = _T_4036 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4457 = _T_4040 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4461 = _T_4012 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4465 = _T_4016 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4469 = _T_4020 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4473 = _T_4024 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4477 = _T_4028 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4481 = _T_4032 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4485 = _T_4036 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4489 = _T_4040 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4493 = _T_4012 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4497 = _T_4016 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4501 = _T_4020 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4505 = _T_4024 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4509 = _T_4028 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4513 = _T_4032 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4517 = _T_4036 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_4521 = _T_4040 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 723:124]
  wire  _T_10394 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 786:84]
  wire  _T_10395 = _T_10394 & miss_pending; // @[el2_ifu_mem_ctl.scala 786:108]
  wire  bus_wren_last_1 = _T_10395 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 786:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 787:84]
  wire  _T_10397 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 788:73]
  wire  _T_10392 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 786:84]
  wire  _T_10393 = _T_10392 & miss_pending; // @[el2_ifu_mem_ctl.scala 786:108]
  wire  bus_wren_last_0 = _T_10393 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 786:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 787:84]
  wire  _T_10396 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 788:73]
  wire [1:0] ifu_tag_wren = {_T_10397,_T_10396}; // @[Cat.scala 29:58]
  wire [1:0] _T_10432 = _T_3990 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10432 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 822:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 732:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 734:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 738:14]
  wire  _T_5170 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 742:82]
  wire  _T_5172 = _T_5170 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5174 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 743:74]
  wire  _T_5176 = _T_5174 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5177 = _T_5172 | _T_5176; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5178 = _T_5177 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire  _T_5182 = _T_5170 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5186 = _T_5174 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5187 = _T_5182 | _T_5186; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5188 = _T_5187 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire [1:0] tag_valid_clken_0 = {_T_5188,_T_5178}; // @[Cat.scala 29:58]
  wire  _T_5190 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 742:82]
  wire  _T_5192 = _T_5190 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5194 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 743:74]
  wire  _T_5196 = _T_5194 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5197 = _T_5192 | _T_5196; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5198 = _T_5197 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire  _T_5202 = _T_5190 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5206 = _T_5194 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5207 = _T_5202 | _T_5206; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5208 = _T_5207 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire [1:0] tag_valid_clken_1 = {_T_5208,_T_5198}; // @[Cat.scala 29:58]
  wire  _T_5210 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 742:82]
  wire  _T_5212 = _T_5210 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5214 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 743:74]
  wire  _T_5216 = _T_5214 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5217 = _T_5212 | _T_5216; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5218 = _T_5217 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire  _T_5222 = _T_5210 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5226 = _T_5214 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5227 = _T_5222 | _T_5226; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5228 = _T_5227 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire [1:0] tag_valid_clken_2 = {_T_5228,_T_5218}; // @[Cat.scala 29:58]
  wire  _T_5230 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 742:82]
  wire  _T_5232 = _T_5230 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5234 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 743:74]
  wire  _T_5236 = _T_5234 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5237 = _T_5232 | _T_5236; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5238 = _T_5237 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire  _T_5242 = _T_5230 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:91]
  wire  _T_5246 = _T_5234 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 743:83]
  wire  _T_5247 = _T_5242 | _T_5246; // @[el2_ifu_mem_ctl.scala 742:113]
  wire  _T_5248 = _T_5247 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 743:106]
  wire [1:0] tag_valid_clken_3 = {_T_5248,_T_5238}; // @[Cat.scala 29:58]
  wire  _T_5251 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 748:64]
  wire  _T_5252 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 748:91]
  wire  _T_5253 = _T_5251 & _T_5252; // @[el2_ifu_mem_ctl.scala 748:89]
  wire  _T_5256 = _T_4523 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5257 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5259 = _T_5257 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5260 = _T_5259 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5262 = _T_5260 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5263 = _T_5256 | _T_5262; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5273 = _T_4527 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5274 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5276 = _T_5274 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5277 = _T_5276 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5279 = _T_5277 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5280 = _T_5273 | _T_5279; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5290 = _T_4531 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5291 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5293 = _T_5291 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5294 = _T_5293 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5296 = _T_5294 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5297 = _T_5290 | _T_5296; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5307 = _T_4535 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5308 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5310 = _T_5308 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5311 = _T_5310 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5313 = _T_5311 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5314 = _T_5307 | _T_5313; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5324 = _T_4539 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5325 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5327 = _T_5325 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5328 = _T_5327 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5330 = _T_5328 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5331 = _T_5324 | _T_5330; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5341 = _T_4543 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5342 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5344 = _T_5342 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5345 = _T_5344 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5347 = _T_5345 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5348 = _T_5341 | _T_5347; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5358 = _T_4547 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5359 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5361 = _T_5359 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5362 = _T_5361 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5364 = _T_5362 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5365 = _T_5358 | _T_5364; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5375 = _T_4551 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5376 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5378 = _T_5376 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5379 = _T_5378 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5381 = _T_5379 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5382 = _T_5375 | _T_5381; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5392 = _T_4555 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5393 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5395 = _T_5393 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5396 = _T_5395 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5398 = _T_5396 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5399 = _T_5392 | _T_5398; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5409 = _T_4559 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5410 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5412 = _T_5410 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5413 = _T_5412 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5415 = _T_5413 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5416 = _T_5409 | _T_5415; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5426 = _T_4563 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5427 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5429 = _T_5427 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5430 = _T_5429 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5432 = _T_5430 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5433 = _T_5426 | _T_5432; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5443 = _T_4567 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5444 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5446 = _T_5444 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5447 = _T_5446 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5449 = _T_5447 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5450 = _T_5443 | _T_5449; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5460 = _T_4571 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5461 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5463 = _T_5461 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5464 = _T_5463 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5466 = _T_5464 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5467 = _T_5460 | _T_5466; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5477 = _T_4575 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5478 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5480 = _T_5478 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5481 = _T_5480 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5483 = _T_5481 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5484 = _T_5477 | _T_5483; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5494 = _T_4579 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5495 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5497 = _T_5495 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5498 = _T_5497 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5500 = _T_5498 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5501 = _T_5494 | _T_5500; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5511 = _T_4583 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5512 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5514 = _T_5512 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5515 = _T_5514 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5517 = _T_5515 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5518 = _T_5511 | _T_5517; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5528 = _T_4587 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5529 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5531 = _T_5529 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5532 = _T_5531 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5534 = _T_5532 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5535 = _T_5528 | _T_5534; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5545 = _T_4591 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5546 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5548 = _T_5546 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5549 = _T_5548 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5551 = _T_5549 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5552 = _T_5545 | _T_5551; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5562 = _T_4595 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5563 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5565 = _T_5563 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5566 = _T_5565 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5568 = _T_5566 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5569 = _T_5562 | _T_5568; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5579 = _T_4599 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5580 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5582 = _T_5580 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5583 = _T_5582 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5585 = _T_5583 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5586 = _T_5579 | _T_5585; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5596 = _T_4603 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5597 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5599 = _T_5597 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5600 = _T_5599 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5602 = _T_5600 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5603 = _T_5596 | _T_5602; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5613 = _T_4607 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5614 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5616 = _T_5614 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5617 = _T_5616 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5619 = _T_5617 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5620 = _T_5613 | _T_5619; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5630 = _T_4611 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5631 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5633 = _T_5631 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5634 = _T_5633 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5636 = _T_5634 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5637 = _T_5630 | _T_5636; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5647 = _T_4615 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5648 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5650 = _T_5648 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5651 = _T_5650 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5653 = _T_5651 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5654 = _T_5647 | _T_5653; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5664 = _T_4619 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5665 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5667 = _T_5665 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5668 = _T_5667 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5670 = _T_5668 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5671 = _T_5664 | _T_5670; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5681 = _T_4623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5682 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5684 = _T_5682 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5685 = _T_5684 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5687 = _T_5685 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5688 = _T_5681 | _T_5687; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5698 = _T_4627 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5699 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5701 = _T_5699 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5702 = _T_5701 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5704 = _T_5702 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5705 = _T_5698 | _T_5704; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5715 = _T_4631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5716 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5718 = _T_5716 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5719 = _T_5718 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5721 = _T_5719 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5722 = _T_5715 | _T_5721; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5732 = _T_4635 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5733 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5735 = _T_5733 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5736 = _T_5735 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5738 = _T_5736 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5739 = _T_5732 | _T_5738; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5749 = _T_4639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5750 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5752 = _T_5750 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5753 = _T_5752 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5755 = _T_5753 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5756 = _T_5749 | _T_5755; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5766 = _T_4643 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5767 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5769 = _T_5767 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5770 = _T_5769 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5772 = _T_5770 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5773 = _T_5766 | _T_5772; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5783 = _T_4647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5784 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_5786 = _T_5784 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5787 = _T_5786 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5789 = _T_5787 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5790 = _T_5783 | _T_5789; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5800 = _T_4523 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5803 = _T_5257 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5804 = _T_5803 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5806 = _T_5804 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5807 = _T_5800 | _T_5806; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5817 = _T_4527 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5820 = _T_5274 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5821 = _T_5820 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5823 = _T_5821 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5824 = _T_5817 | _T_5823; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5834 = _T_4531 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5837 = _T_5291 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5838 = _T_5837 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5840 = _T_5838 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5841 = _T_5834 | _T_5840; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5851 = _T_4535 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5854 = _T_5308 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5855 = _T_5854 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5857 = _T_5855 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5858 = _T_5851 | _T_5857; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5868 = _T_4539 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5871 = _T_5325 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5872 = _T_5871 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5874 = _T_5872 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5875 = _T_5868 | _T_5874; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5885 = _T_4543 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5888 = _T_5342 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5889 = _T_5888 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5891 = _T_5889 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5892 = _T_5885 | _T_5891; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5902 = _T_4547 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5905 = _T_5359 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5906 = _T_5905 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5908 = _T_5906 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5909 = _T_5902 | _T_5908; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5919 = _T_4551 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5922 = _T_5376 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5923 = _T_5922 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5925 = _T_5923 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5926 = _T_5919 | _T_5925; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5936 = _T_4555 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5939 = _T_5393 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5940 = _T_5939 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5942 = _T_5940 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5943 = _T_5936 | _T_5942; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5953 = _T_4559 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5956 = _T_5410 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5957 = _T_5956 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5959 = _T_5957 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5960 = _T_5953 | _T_5959; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5970 = _T_4563 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5973 = _T_5427 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5974 = _T_5973 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5976 = _T_5974 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5977 = _T_5970 | _T_5976; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_5987 = _T_4567 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_5990 = _T_5444 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_5991 = _T_5990 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_5993 = _T_5991 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_5994 = _T_5987 | _T_5993; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6004 = _T_4571 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6007 = _T_5461 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6008 = _T_6007 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6010 = _T_6008 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6011 = _T_6004 | _T_6010; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6021 = _T_4575 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6024 = _T_5478 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6025 = _T_6024 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6027 = _T_6025 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6028 = _T_6021 | _T_6027; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6038 = _T_4579 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6041 = _T_5495 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6042 = _T_6041 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6044 = _T_6042 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6045 = _T_6038 | _T_6044; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6055 = _T_4583 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6058 = _T_5512 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6059 = _T_6058 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6061 = _T_6059 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6062 = _T_6055 | _T_6061; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6072 = _T_4587 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6075 = _T_5529 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6076 = _T_6075 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6078 = _T_6076 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6079 = _T_6072 | _T_6078; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6089 = _T_4591 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6092 = _T_5546 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6093 = _T_6092 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6095 = _T_6093 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6096 = _T_6089 | _T_6095; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6106 = _T_4595 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6109 = _T_5563 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6110 = _T_6109 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6112 = _T_6110 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6113 = _T_6106 | _T_6112; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6123 = _T_4599 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6126 = _T_5580 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6127 = _T_6126 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6129 = _T_6127 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6130 = _T_6123 | _T_6129; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6140 = _T_4603 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6143 = _T_5597 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6144 = _T_6143 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6146 = _T_6144 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6147 = _T_6140 | _T_6146; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6157 = _T_4607 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6160 = _T_5614 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6161 = _T_6160 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6163 = _T_6161 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6164 = _T_6157 | _T_6163; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6174 = _T_4611 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6177 = _T_5631 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6178 = _T_6177 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6180 = _T_6178 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6181 = _T_6174 | _T_6180; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6191 = _T_4615 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6194 = _T_5648 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6195 = _T_6194 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6197 = _T_6195 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6198 = _T_6191 | _T_6197; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6208 = _T_4619 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6211 = _T_5665 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6212 = _T_6211 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6214 = _T_6212 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6215 = _T_6208 | _T_6214; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6225 = _T_4623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6228 = _T_5682 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6229 = _T_6228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6231 = _T_6229 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6232 = _T_6225 | _T_6231; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6242 = _T_4627 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6245 = _T_5699 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6246 = _T_6245 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6248 = _T_6246 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6249 = _T_6242 | _T_6248; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6259 = _T_4631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6262 = _T_5716 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6263 = _T_6262 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6265 = _T_6263 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6266 = _T_6259 | _T_6265; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6276 = _T_4635 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6279 = _T_5733 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6280 = _T_6279 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6282 = _T_6280 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6283 = _T_6276 | _T_6282; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6293 = _T_4639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6296 = _T_5750 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6297 = _T_6296 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6299 = _T_6297 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6300 = _T_6293 | _T_6299; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6310 = _T_4643 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6313 = _T_5767 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6314 = _T_6313 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6316 = _T_6314 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6317 = _T_6310 | _T_6316; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6327 = _T_4647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6330 = _T_5784 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6331 = _T_6330 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6333 = _T_6331 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6334 = _T_6327 | _T_6333; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6344 = _T_4651 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6345 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6347 = _T_6345 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6348 = _T_6347 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6350 = _T_6348 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6351 = _T_6344 | _T_6350; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6361 = _T_4655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6362 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6364 = _T_6362 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6365 = _T_6364 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6367 = _T_6365 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6368 = _T_6361 | _T_6367; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6378 = _T_4659 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6379 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6381 = _T_6379 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6382 = _T_6381 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6384 = _T_6382 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6385 = _T_6378 | _T_6384; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6395 = _T_4663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6396 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6398 = _T_6396 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6399 = _T_6398 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6401 = _T_6399 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6402 = _T_6395 | _T_6401; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6412 = _T_4667 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6413 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6415 = _T_6413 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6416 = _T_6415 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6418 = _T_6416 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6419 = _T_6412 | _T_6418; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6429 = _T_4671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6430 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6432 = _T_6430 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6433 = _T_6432 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6435 = _T_6433 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6436 = _T_6429 | _T_6435; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6446 = _T_4675 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6447 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6449 = _T_6447 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6450 = _T_6449 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6452 = _T_6450 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6453 = _T_6446 | _T_6452; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6463 = _T_4679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6464 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6466 = _T_6464 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6467 = _T_6466 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6469 = _T_6467 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6470 = _T_6463 | _T_6469; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6480 = _T_4683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6481 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6483 = _T_6481 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6484 = _T_6483 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6486 = _T_6484 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6487 = _T_6480 | _T_6486; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6497 = _T_4687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6498 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6500 = _T_6498 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6501 = _T_6500 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6503 = _T_6501 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6504 = _T_6497 | _T_6503; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6514 = _T_4691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6515 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6517 = _T_6515 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6518 = _T_6517 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6520 = _T_6518 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6521 = _T_6514 | _T_6520; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6531 = _T_4695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6532 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6534 = _T_6532 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6535 = _T_6534 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6537 = _T_6535 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6538 = _T_6531 | _T_6537; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6548 = _T_4699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6549 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6551 = _T_6549 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6552 = _T_6551 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6554 = _T_6552 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6555 = _T_6548 | _T_6554; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6565 = _T_4703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6566 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6568 = _T_6566 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6569 = _T_6568 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6571 = _T_6569 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6572 = _T_6565 | _T_6571; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6582 = _T_4707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6583 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6585 = _T_6583 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6586 = _T_6585 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6588 = _T_6586 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6589 = _T_6582 | _T_6588; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6599 = _T_4711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6600 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6602 = _T_6600 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6603 = _T_6602 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6605 = _T_6603 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6606 = _T_6599 | _T_6605; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6616 = _T_4715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6617 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6619 = _T_6617 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6620 = _T_6619 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6622 = _T_6620 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6623 = _T_6616 | _T_6622; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6633 = _T_4719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6634 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6636 = _T_6634 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6637 = _T_6636 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6639 = _T_6637 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6640 = _T_6633 | _T_6639; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6650 = _T_4723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6651 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6653 = _T_6651 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6654 = _T_6653 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6656 = _T_6654 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6657 = _T_6650 | _T_6656; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6667 = _T_4727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6668 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6670 = _T_6668 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6671 = _T_6670 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6673 = _T_6671 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6674 = _T_6667 | _T_6673; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6684 = _T_4731 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6685 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6687 = _T_6685 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6688 = _T_6687 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6690 = _T_6688 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6691 = _T_6684 | _T_6690; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6701 = _T_4735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6702 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6704 = _T_6702 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6705 = _T_6704 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6707 = _T_6705 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6708 = _T_6701 | _T_6707; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6718 = _T_4739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6719 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6721 = _T_6719 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6722 = _T_6721 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6724 = _T_6722 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6725 = _T_6718 | _T_6724; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6735 = _T_4743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6736 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6738 = _T_6736 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6739 = _T_6738 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6741 = _T_6739 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6742 = _T_6735 | _T_6741; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6752 = _T_4747 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6753 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6755 = _T_6753 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6756 = _T_6755 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6758 = _T_6756 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6759 = _T_6752 | _T_6758; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6769 = _T_4751 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6770 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6772 = _T_6770 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6773 = _T_6772 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6775 = _T_6773 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6776 = _T_6769 | _T_6775; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6786 = _T_4755 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6787 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6789 = _T_6787 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6790 = _T_6789 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6792 = _T_6790 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6793 = _T_6786 | _T_6792; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6803 = _T_4759 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6804 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6806 = _T_6804 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6807 = _T_6806 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6809 = _T_6807 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6810 = _T_6803 | _T_6809; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6820 = _T_4763 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6821 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6823 = _T_6821 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6824 = _T_6823 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6826 = _T_6824 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6827 = _T_6820 | _T_6826; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6837 = _T_4767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6838 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6840 = _T_6838 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6841 = _T_6840 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6843 = _T_6841 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6844 = _T_6837 | _T_6843; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6854 = _T_4771 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6855 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6857 = _T_6855 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6858 = _T_6857 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6860 = _T_6858 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6861 = _T_6854 | _T_6860; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6871 = _T_4775 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6872 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_6874 = _T_6872 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6875 = _T_6874 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6877 = _T_6875 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6878 = _T_6871 | _T_6877; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6888 = _T_4651 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6891 = _T_6345 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6892 = _T_6891 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6894 = _T_6892 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6895 = _T_6888 | _T_6894; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6905 = _T_4655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6908 = _T_6362 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6909 = _T_6908 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6911 = _T_6909 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6912 = _T_6905 | _T_6911; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6922 = _T_4659 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6925 = _T_6379 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6926 = _T_6925 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6928 = _T_6926 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6929 = _T_6922 | _T_6928; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6939 = _T_4663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6942 = _T_6396 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6943 = _T_6942 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6945 = _T_6943 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6946 = _T_6939 | _T_6945; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6956 = _T_4667 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6959 = _T_6413 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6960 = _T_6959 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6962 = _T_6960 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6963 = _T_6956 | _T_6962; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6973 = _T_4671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6976 = _T_6430 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6977 = _T_6976 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6979 = _T_6977 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6980 = _T_6973 | _T_6979; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_6990 = _T_4675 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_6993 = _T_6447 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_6994 = _T_6993 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_6996 = _T_6994 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_6997 = _T_6990 | _T_6996; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7007 = _T_4679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7010 = _T_6464 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7011 = _T_7010 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7013 = _T_7011 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7014 = _T_7007 | _T_7013; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7024 = _T_4683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7027 = _T_6481 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7028 = _T_7027 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7030 = _T_7028 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7031 = _T_7024 | _T_7030; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7041 = _T_4687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7044 = _T_6498 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7045 = _T_7044 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7047 = _T_7045 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7048 = _T_7041 | _T_7047; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7058 = _T_4691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7061 = _T_6515 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7062 = _T_7061 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7064 = _T_7062 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7065 = _T_7058 | _T_7064; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7075 = _T_4695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7078 = _T_6532 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7079 = _T_7078 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7081 = _T_7079 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7082 = _T_7075 | _T_7081; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7092 = _T_4699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7095 = _T_6549 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7096 = _T_7095 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7098 = _T_7096 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7099 = _T_7092 | _T_7098; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7109 = _T_4703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7112 = _T_6566 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7113 = _T_7112 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7115 = _T_7113 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7116 = _T_7109 | _T_7115; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7126 = _T_4707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7129 = _T_6583 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7130 = _T_7129 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7132 = _T_7130 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7133 = _T_7126 | _T_7132; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7143 = _T_4711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7146 = _T_6600 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7147 = _T_7146 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7149 = _T_7147 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7150 = _T_7143 | _T_7149; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7160 = _T_4715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7163 = _T_6617 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7164 = _T_7163 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7166 = _T_7164 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7167 = _T_7160 | _T_7166; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7177 = _T_4719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7180 = _T_6634 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7181 = _T_7180 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7183 = _T_7181 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7184 = _T_7177 | _T_7183; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7194 = _T_4723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7197 = _T_6651 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7198 = _T_7197 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7200 = _T_7198 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7201 = _T_7194 | _T_7200; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7211 = _T_4727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7214 = _T_6668 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7215 = _T_7214 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7217 = _T_7215 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7218 = _T_7211 | _T_7217; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7228 = _T_4731 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7231 = _T_6685 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7232 = _T_7231 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7234 = _T_7232 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7235 = _T_7228 | _T_7234; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7245 = _T_4735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7248 = _T_6702 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7249 = _T_7248 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7251 = _T_7249 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7252 = _T_7245 | _T_7251; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7262 = _T_4739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7265 = _T_6719 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7266 = _T_7265 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7268 = _T_7266 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7269 = _T_7262 | _T_7268; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7279 = _T_4743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7282 = _T_6736 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7283 = _T_7282 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7285 = _T_7283 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7286 = _T_7279 | _T_7285; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7296 = _T_4747 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7299 = _T_6753 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7300 = _T_7299 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7302 = _T_7300 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7303 = _T_7296 | _T_7302; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7313 = _T_4751 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7316 = _T_6770 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7317 = _T_7316 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7319 = _T_7317 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7320 = _T_7313 | _T_7319; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7330 = _T_4755 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7333 = _T_6787 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7334 = _T_7333 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7336 = _T_7334 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7337 = _T_7330 | _T_7336; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7347 = _T_4759 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7350 = _T_6804 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7351 = _T_7350 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7353 = _T_7351 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7354 = _T_7347 | _T_7353; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7364 = _T_4763 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7367 = _T_6821 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7368 = _T_7367 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7370 = _T_7368 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7371 = _T_7364 | _T_7370; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7381 = _T_4767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7384 = _T_6838 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7385 = _T_7384 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7387 = _T_7385 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7388 = _T_7381 | _T_7387; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7398 = _T_4771 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7401 = _T_6855 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7402 = _T_7401 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7404 = _T_7402 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7405 = _T_7398 | _T_7404; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7415 = _T_4775 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7418 = _T_6872 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7419 = _T_7418 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7421 = _T_7419 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7422 = _T_7415 | _T_7421; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7432 = _T_4779 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire [6:0] _GEN_797 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7433 = _GEN_797 == 7'h40; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7435 = _T_7433 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7436 = _T_7435 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7438 = _T_7436 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7439 = _T_7432 | _T_7438; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7449 = _T_4783 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7450 = _GEN_797 == 7'h41; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7452 = _T_7450 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7453 = _T_7452 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7455 = _T_7453 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7456 = _T_7449 | _T_7455; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7466 = _T_4787 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7467 = _GEN_797 == 7'h42; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7469 = _T_7467 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7470 = _T_7469 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7472 = _T_7470 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7473 = _T_7466 | _T_7472; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7483 = _T_4791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7484 = _GEN_797 == 7'h43; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7486 = _T_7484 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7487 = _T_7486 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7489 = _T_7487 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7490 = _T_7483 | _T_7489; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7500 = _T_4795 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7501 = _GEN_797 == 7'h44; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7503 = _T_7501 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7504 = _T_7503 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7506 = _T_7504 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7507 = _T_7500 | _T_7506; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7517 = _T_4799 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7518 = _GEN_797 == 7'h45; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7520 = _T_7518 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7521 = _T_7520 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7523 = _T_7521 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7524 = _T_7517 | _T_7523; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7534 = _T_4803 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7535 = _GEN_797 == 7'h46; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7537 = _T_7535 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7538 = _T_7537 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7540 = _T_7538 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7541 = _T_7534 | _T_7540; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7551 = _T_4807 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7552 = _GEN_797 == 7'h47; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7554 = _T_7552 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7555 = _T_7554 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7557 = _T_7555 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7558 = _T_7551 | _T_7557; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7568 = _T_4811 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7569 = _GEN_797 == 7'h48; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7571 = _T_7569 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7572 = _T_7571 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7574 = _T_7572 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7575 = _T_7568 | _T_7574; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7585 = _T_4815 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7586 = _GEN_797 == 7'h49; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7588 = _T_7586 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7589 = _T_7588 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7591 = _T_7589 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7592 = _T_7585 | _T_7591; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7602 = _T_4819 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7603 = _GEN_797 == 7'h4a; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7605 = _T_7603 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7606 = _T_7605 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7608 = _T_7606 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7609 = _T_7602 | _T_7608; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7619 = _T_4823 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7620 = _GEN_797 == 7'h4b; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7622 = _T_7620 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7623 = _T_7622 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7625 = _T_7623 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7626 = _T_7619 | _T_7625; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7636 = _T_4827 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7637 = _GEN_797 == 7'h4c; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7639 = _T_7637 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7640 = _T_7639 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7642 = _T_7640 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7643 = _T_7636 | _T_7642; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7653 = _T_4831 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7654 = _GEN_797 == 7'h4d; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7656 = _T_7654 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7657 = _T_7656 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7659 = _T_7657 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7660 = _T_7653 | _T_7659; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7670 = _T_4835 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7671 = _GEN_797 == 7'h4e; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7673 = _T_7671 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7674 = _T_7673 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7676 = _T_7674 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7677 = _T_7670 | _T_7676; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7687 = _T_4839 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7688 = _GEN_797 == 7'h4f; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7690 = _T_7688 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7691 = _T_7690 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7693 = _T_7691 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7694 = _T_7687 | _T_7693; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7704 = _T_4843 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7705 = _GEN_797 == 7'h50; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7707 = _T_7705 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7708 = _T_7707 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7710 = _T_7708 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7711 = _T_7704 | _T_7710; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7721 = _T_4847 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7722 = _GEN_797 == 7'h51; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7724 = _T_7722 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7725 = _T_7724 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7727 = _T_7725 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7728 = _T_7721 | _T_7727; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7738 = _T_4851 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7739 = _GEN_797 == 7'h52; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7741 = _T_7739 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7742 = _T_7741 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7744 = _T_7742 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7745 = _T_7738 | _T_7744; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7755 = _T_4855 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7756 = _GEN_797 == 7'h53; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7758 = _T_7756 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7759 = _T_7758 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7761 = _T_7759 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7762 = _T_7755 | _T_7761; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7772 = _T_4859 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7773 = _GEN_797 == 7'h54; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7775 = _T_7773 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7776 = _T_7775 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7778 = _T_7776 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7779 = _T_7772 | _T_7778; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7789 = _T_4863 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7790 = _GEN_797 == 7'h55; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7792 = _T_7790 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7793 = _T_7792 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7795 = _T_7793 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7796 = _T_7789 | _T_7795; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7806 = _T_4867 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7807 = _GEN_797 == 7'h56; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7809 = _T_7807 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7810 = _T_7809 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7812 = _T_7810 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7813 = _T_7806 | _T_7812; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7823 = _T_4871 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7824 = _GEN_797 == 7'h57; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7826 = _T_7824 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7827 = _T_7826 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7829 = _T_7827 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7830 = _T_7823 | _T_7829; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7840 = _T_4875 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7841 = _GEN_797 == 7'h58; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7843 = _T_7841 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7844 = _T_7843 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7846 = _T_7844 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7847 = _T_7840 | _T_7846; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7857 = _T_4879 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7858 = _GEN_797 == 7'h59; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7860 = _T_7858 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7861 = _T_7860 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7863 = _T_7861 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7864 = _T_7857 | _T_7863; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7874 = _T_4883 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7875 = _GEN_797 == 7'h5a; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7877 = _T_7875 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7878 = _T_7877 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7880 = _T_7878 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7881 = _T_7874 | _T_7880; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7891 = _T_4887 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7892 = _GEN_797 == 7'h5b; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7894 = _T_7892 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7895 = _T_7894 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7897 = _T_7895 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7898 = _T_7891 | _T_7897; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7908 = _T_4891 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7909 = _GEN_797 == 7'h5c; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7911 = _T_7909 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7912 = _T_7911 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7914 = _T_7912 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7915 = _T_7908 | _T_7914; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7925 = _T_4895 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7926 = _GEN_797 == 7'h5d; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7928 = _T_7926 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7929 = _T_7928 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7931 = _T_7929 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7932 = _T_7925 | _T_7931; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7942 = _T_4899 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7943 = _GEN_797 == 7'h5e; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7945 = _T_7943 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7946 = _T_7945 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7948 = _T_7946 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7949 = _T_7942 | _T_7948; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7959 = _T_4903 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7960 = _GEN_797 == 7'h5f; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_7962 = _T_7960 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7963 = _T_7962 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7965 = _T_7963 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7966 = _T_7959 | _T_7965; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7976 = _T_4779 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7979 = _T_7433 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7980 = _T_7979 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7982 = _T_7980 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_7983 = _T_7976 | _T_7982; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_7993 = _T_4783 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_7996 = _T_7450 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_7997 = _T_7996 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_7999 = _T_7997 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8000 = _T_7993 | _T_7999; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8010 = _T_4787 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8013 = _T_7467 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8014 = _T_8013 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8016 = _T_8014 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8017 = _T_8010 | _T_8016; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8027 = _T_4791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8030 = _T_7484 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8031 = _T_8030 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8033 = _T_8031 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8034 = _T_8027 | _T_8033; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8044 = _T_4795 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8047 = _T_7501 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8048 = _T_8047 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8050 = _T_8048 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8051 = _T_8044 | _T_8050; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8061 = _T_4799 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8064 = _T_7518 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8065 = _T_8064 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8067 = _T_8065 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8068 = _T_8061 | _T_8067; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8078 = _T_4803 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8081 = _T_7535 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8082 = _T_8081 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8084 = _T_8082 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8085 = _T_8078 | _T_8084; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8095 = _T_4807 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8098 = _T_7552 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8099 = _T_8098 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8101 = _T_8099 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8102 = _T_8095 | _T_8101; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8112 = _T_4811 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8115 = _T_7569 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8116 = _T_8115 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8118 = _T_8116 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8119 = _T_8112 | _T_8118; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8129 = _T_4815 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8132 = _T_7586 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8133 = _T_8132 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8135 = _T_8133 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8136 = _T_8129 | _T_8135; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8146 = _T_4819 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8149 = _T_7603 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8150 = _T_8149 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8152 = _T_8150 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8153 = _T_8146 | _T_8152; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8163 = _T_4823 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8166 = _T_7620 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8167 = _T_8166 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8169 = _T_8167 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8170 = _T_8163 | _T_8169; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8180 = _T_4827 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8183 = _T_7637 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8184 = _T_8183 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8186 = _T_8184 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8187 = _T_8180 | _T_8186; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8197 = _T_4831 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8200 = _T_7654 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8201 = _T_8200 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8203 = _T_8201 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8204 = _T_8197 | _T_8203; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8214 = _T_4835 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8217 = _T_7671 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8218 = _T_8217 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8220 = _T_8218 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8221 = _T_8214 | _T_8220; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8231 = _T_4839 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8234 = _T_7688 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8235 = _T_8234 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8237 = _T_8235 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8238 = _T_8231 | _T_8237; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8248 = _T_4843 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8251 = _T_7705 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8252 = _T_8251 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8254 = _T_8252 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8255 = _T_8248 | _T_8254; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8265 = _T_4847 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8268 = _T_7722 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8269 = _T_8268 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8271 = _T_8269 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8272 = _T_8265 | _T_8271; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8282 = _T_4851 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8285 = _T_7739 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8286 = _T_8285 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8288 = _T_8286 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8289 = _T_8282 | _T_8288; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8299 = _T_4855 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8302 = _T_7756 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8303 = _T_8302 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8305 = _T_8303 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8306 = _T_8299 | _T_8305; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8316 = _T_4859 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8319 = _T_7773 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8320 = _T_8319 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8322 = _T_8320 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8323 = _T_8316 | _T_8322; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8333 = _T_4863 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8336 = _T_7790 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8337 = _T_8336 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8339 = _T_8337 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8340 = _T_8333 | _T_8339; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8350 = _T_4867 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8353 = _T_7807 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8354 = _T_8353 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8356 = _T_8354 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8357 = _T_8350 | _T_8356; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8367 = _T_4871 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8370 = _T_7824 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8371 = _T_8370 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8373 = _T_8371 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8374 = _T_8367 | _T_8373; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8384 = _T_4875 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8387 = _T_7841 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8388 = _T_8387 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8390 = _T_8388 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8391 = _T_8384 | _T_8390; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8401 = _T_4879 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8404 = _T_7858 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8405 = _T_8404 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8407 = _T_8405 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8408 = _T_8401 | _T_8407; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8418 = _T_4883 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8421 = _T_7875 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8422 = _T_8421 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8424 = _T_8422 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8425 = _T_8418 | _T_8424; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8435 = _T_4887 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8438 = _T_7892 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8439 = _T_8438 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8441 = _T_8439 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8442 = _T_8435 | _T_8441; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8452 = _T_4891 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8455 = _T_7909 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8456 = _T_8455 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8458 = _T_8456 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8459 = _T_8452 | _T_8458; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8469 = _T_4895 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8472 = _T_7926 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8473 = _T_8472 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8475 = _T_8473 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8476 = _T_8469 | _T_8475; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8486 = _T_4899 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8489 = _T_7943 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8490 = _T_8489 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8492 = _T_8490 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8493 = _T_8486 | _T_8492; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8503 = _T_4903 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8506 = _T_7960 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8507 = _T_8506 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8509 = _T_8507 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8510 = _T_8503 | _T_8509; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8520 = _T_4907 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8521 = _GEN_797 == 7'h60; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8523 = _T_8521 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8524 = _T_8523 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8526 = _T_8524 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8527 = _T_8520 | _T_8526; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8537 = _T_4911 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8538 = _GEN_797 == 7'h61; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8540 = _T_8538 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8541 = _T_8540 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8543 = _T_8541 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8544 = _T_8537 | _T_8543; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8554 = _T_4915 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8555 = _GEN_797 == 7'h62; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8557 = _T_8555 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8558 = _T_8557 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8560 = _T_8558 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8561 = _T_8554 | _T_8560; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8571 = _T_4919 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8572 = _GEN_797 == 7'h63; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8574 = _T_8572 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8575 = _T_8574 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8577 = _T_8575 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8578 = _T_8571 | _T_8577; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8588 = _T_4923 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8589 = _GEN_797 == 7'h64; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8591 = _T_8589 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8592 = _T_8591 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8594 = _T_8592 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8595 = _T_8588 | _T_8594; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8605 = _T_4927 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8606 = _GEN_797 == 7'h65; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8608 = _T_8606 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8609 = _T_8608 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8611 = _T_8609 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8612 = _T_8605 | _T_8611; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8622 = _T_4931 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8623 = _GEN_797 == 7'h66; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8625 = _T_8623 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8626 = _T_8625 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8628 = _T_8626 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8629 = _T_8622 | _T_8628; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8639 = _T_4935 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8640 = _GEN_797 == 7'h67; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8642 = _T_8640 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8643 = _T_8642 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8645 = _T_8643 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8646 = _T_8639 | _T_8645; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8656 = _T_4939 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8657 = _GEN_797 == 7'h68; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8659 = _T_8657 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8660 = _T_8659 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8662 = _T_8660 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8663 = _T_8656 | _T_8662; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8673 = _T_4943 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8674 = _GEN_797 == 7'h69; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8676 = _T_8674 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8677 = _T_8676 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8679 = _T_8677 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8680 = _T_8673 | _T_8679; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8690 = _T_4947 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8691 = _GEN_797 == 7'h6a; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8693 = _T_8691 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8694 = _T_8693 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8696 = _T_8694 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8697 = _T_8690 | _T_8696; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8707 = _T_4951 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8708 = _GEN_797 == 7'h6b; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8710 = _T_8708 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8711 = _T_8710 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8713 = _T_8711 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8714 = _T_8707 | _T_8713; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8724 = _T_4955 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8725 = _GEN_797 == 7'h6c; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8727 = _T_8725 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8728 = _T_8727 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8730 = _T_8728 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8731 = _T_8724 | _T_8730; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8741 = _T_4959 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8742 = _GEN_797 == 7'h6d; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8744 = _T_8742 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8745 = _T_8744 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8747 = _T_8745 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8748 = _T_8741 | _T_8747; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8758 = _T_4963 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8759 = _GEN_797 == 7'h6e; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8761 = _T_8759 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8762 = _T_8761 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8764 = _T_8762 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8765 = _T_8758 | _T_8764; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8775 = _T_4967 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8776 = _GEN_797 == 7'h6f; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8778 = _T_8776 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8779 = _T_8778 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8781 = _T_8779 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8782 = _T_8775 | _T_8781; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8792 = _T_4971 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8793 = _GEN_797 == 7'h70; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8795 = _T_8793 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8796 = _T_8795 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8798 = _T_8796 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8799 = _T_8792 | _T_8798; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8809 = _T_4975 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8810 = _GEN_797 == 7'h71; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8812 = _T_8810 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8813 = _T_8812 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8815 = _T_8813 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8816 = _T_8809 | _T_8815; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8826 = _T_4979 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8827 = _GEN_797 == 7'h72; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8829 = _T_8827 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8830 = _T_8829 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8832 = _T_8830 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8833 = _T_8826 | _T_8832; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8843 = _T_4983 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8844 = _GEN_797 == 7'h73; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8846 = _T_8844 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8847 = _T_8846 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8849 = _T_8847 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8850 = _T_8843 | _T_8849; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8860 = _T_4987 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8861 = _GEN_797 == 7'h74; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8863 = _T_8861 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8864 = _T_8863 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8866 = _T_8864 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8867 = _T_8860 | _T_8866; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8877 = _T_4991 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8878 = _GEN_797 == 7'h75; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8880 = _T_8878 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8881 = _T_8880 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8883 = _T_8881 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8884 = _T_8877 | _T_8883; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8894 = _T_4995 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8895 = _GEN_797 == 7'h76; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8897 = _T_8895 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8898 = _T_8897 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8900 = _T_8898 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8901 = _T_8894 | _T_8900; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8911 = _T_4999 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8912 = _GEN_797 == 7'h77; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8914 = _T_8912 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8915 = _T_8914 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8917 = _T_8915 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8918 = _T_8911 | _T_8917; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8928 = _T_5003 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8929 = _GEN_797 == 7'h78; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8931 = _T_8929 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8932 = _T_8931 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8934 = _T_8932 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8935 = _T_8928 | _T_8934; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8945 = _T_5007 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8946 = _GEN_797 == 7'h79; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8948 = _T_8946 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8949 = _T_8948 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8951 = _T_8949 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8952 = _T_8945 | _T_8951; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8962 = _T_5011 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8963 = _GEN_797 == 7'h7a; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8965 = _T_8963 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8966 = _T_8965 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8968 = _T_8966 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8969 = _T_8962 | _T_8968; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8979 = _T_5015 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8980 = _GEN_797 == 7'h7b; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8982 = _T_8980 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_8983 = _T_8982 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_8985 = _T_8983 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_8986 = _T_8979 | _T_8985; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_8996 = _T_5019 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_8997 = _GEN_797 == 7'h7c; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_8999 = _T_8997 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9000 = _T_8999 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9002 = _T_9000 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9003 = _T_8996 | _T_9002; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9013 = _T_5023 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9014 = _GEN_797 == 7'h7d; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_9016 = _T_9014 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9017 = _T_9016 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9019 = _T_9017 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9020 = _T_9013 | _T_9019; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9030 = _T_5027 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9031 = _GEN_797 == 7'h7e; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_9033 = _T_9031 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9034 = _T_9033 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9036 = _T_9034 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9037 = _T_9030 | _T_9036; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9047 = _T_5031 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9048 = _GEN_797 == 7'h7f; // @[el2_ifu_mem_ctl.scala 749:101]
  wire  _T_9050 = _T_9048 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9051 = _T_9050 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9053 = _T_9051 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9054 = _T_9047 | _T_9053; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9064 = _T_4907 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9067 = _T_8521 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9068 = _T_9067 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9070 = _T_9068 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9071 = _T_9064 | _T_9070; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9081 = _T_4911 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9084 = _T_8538 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9085 = _T_9084 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9087 = _T_9085 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9088 = _T_9081 | _T_9087; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9098 = _T_4915 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9101 = _T_8555 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9102 = _T_9101 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9104 = _T_9102 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9105 = _T_9098 | _T_9104; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9115 = _T_4919 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9118 = _T_8572 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9119 = _T_9118 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9121 = _T_9119 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9122 = _T_9115 | _T_9121; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9132 = _T_4923 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9135 = _T_8589 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9136 = _T_9135 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9138 = _T_9136 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9139 = _T_9132 | _T_9138; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9149 = _T_4927 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9152 = _T_8606 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9153 = _T_9152 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9155 = _T_9153 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9156 = _T_9149 | _T_9155; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9166 = _T_4931 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9169 = _T_8623 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9170 = _T_9169 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9172 = _T_9170 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9173 = _T_9166 | _T_9172; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9183 = _T_4935 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9186 = _T_8640 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9187 = _T_9186 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9189 = _T_9187 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9190 = _T_9183 | _T_9189; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9200 = _T_4939 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9203 = _T_8657 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9204 = _T_9203 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9206 = _T_9204 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9207 = _T_9200 | _T_9206; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9217 = _T_4943 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9220 = _T_8674 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9221 = _T_9220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9223 = _T_9221 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9224 = _T_9217 | _T_9223; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9234 = _T_4947 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9237 = _T_8691 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9238 = _T_9237 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9240 = _T_9238 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9241 = _T_9234 | _T_9240; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9251 = _T_4951 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9254 = _T_8708 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9255 = _T_9254 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9257 = _T_9255 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9258 = _T_9251 | _T_9257; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9268 = _T_4955 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9271 = _T_8725 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9272 = _T_9271 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9274 = _T_9272 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9275 = _T_9268 | _T_9274; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9285 = _T_4959 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9288 = _T_8742 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9289 = _T_9288 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9291 = _T_9289 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9292 = _T_9285 | _T_9291; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9302 = _T_4963 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9305 = _T_8759 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9306 = _T_9305 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9308 = _T_9306 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9309 = _T_9302 | _T_9308; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9319 = _T_4967 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9322 = _T_8776 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9323 = _T_9322 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9325 = _T_9323 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9326 = _T_9319 | _T_9325; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9336 = _T_4971 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9339 = _T_8793 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9340 = _T_9339 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9342 = _T_9340 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9343 = _T_9336 | _T_9342; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9353 = _T_4975 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9356 = _T_8810 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9357 = _T_9356 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9359 = _T_9357 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9360 = _T_9353 | _T_9359; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9370 = _T_4979 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9373 = _T_8827 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9374 = _T_9373 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9376 = _T_9374 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9377 = _T_9370 | _T_9376; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9387 = _T_4983 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9390 = _T_8844 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9391 = _T_9390 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9393 = _T_9391 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9394 = _T_9387 | _T_9393; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9404 = _T_4987 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9407 = _T_8861 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9408 = _T_9407 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9410 = _T_9408 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9411 = _T_9404 | _T_9410; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9421 = _T_4991 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9424 = _T_8878 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9425 = _T_9424 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9427 = _T_9425 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9428 = _T_9421 | _T_9427; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9438 = _T_4995 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9441 = _T_8895 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9442 = _T_9441 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9444 = _T_9442 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9445 = _T_9438 | _T_9444; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9455 = _T_4999 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9458 = _T_8912 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9459 = _T_9458 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9461 = _T_9459 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9462 = _T_9455 | _T_9461; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9472 = _T_5003 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9475 = _T_8929 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9476 = _T_9475 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9478 = _T_9476 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9479 = _T_9472 | _T_9478; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9489 = _T_5007 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9492 = _T_8946 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9493 = _T_9492 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9495 = _T_9493 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9496 = _T_9489 | _T_9495; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9506 = _T_5011 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9509 = _T_8963 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9510 = _T_9509 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9512 = _T_9510 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9513 = _T_9506 | _T_9512; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9523 = _T_5015 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9526 = _T_8980 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9527 = _T_9526 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9529 = _T_9527 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9530 = _T_9523 | _T_9529; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9540 = _T_5019 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9543 = _T_8997 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9544 = _T_9543 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9546 = _T_9544 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9547 = _T_9540 | _T_9546; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9557 = _T_5023 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9560 = _T_9014 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9561 = _T_9560 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9563 = _T_9561 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9564 = _T_9557 | _T_9563; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9574 = _T_5027 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9577 = _T_9031 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9578 = _T_9577 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9580 = _T_9578 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9581 = _T_9574 | _T_9580; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_9591 = _T_5031 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 749:58]
  wire  _T_9594 = _T_9048 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:123]
  wire  _T_9595 = _T_9594 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:145]
  wire  _T_9597 = _T_9595 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 749:163]
  wire  _T_9598 = _T_9591 | _T_9597; // @[el2_ifu_mem_ctl.scala 749:80]
  wire  _T_10400 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 804:63]
  wire  _T_10401 = _T_10400 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 804:85]
  wire [1:0] _T_10403 = _T_10401 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10410; // @[el2_ifu_mem_ctl.scala 809:57]
  reg  _T_10411; // @[el2_ifu_mem_ctl.scala 810:56]
  reg  _T_10412; // @[el2_ifu_mem_ctl.scala 811:59]
  wire  _T_10413 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 812:80]
  wire  _T_10414 = ifu_bus_arvalid_ff & _T_10413; // @[el2_ifu_mem_ctl.scala 812:78]
  wire  _T_10415 = _T_10414 & miss_pending; // @[el2_ifu_mem_ctl.scala 812:100]
  reg  _T_10416; // @[el2_ifu_mem_ctl.scala 812:58]
  reg  _T_10417; // @[el2_ifu_mem_ctl.scala 813:58]
  wire  _T_10420 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 820:71]
  wire  _T_10422 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 820:124]
  wire  _T_10424 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 821:50]
  wire  _T_10426 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 821:103]
  wire [3:0] _T_10429 = {_T_10420,_T_10422,_T_10424,_T_10426}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 823:53]
  reg  _T_10440; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 329:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 328:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 192:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3978; // @[el2_ifu_mem_ctl.scala 699:21]
  assign io_ifu_pmu_ic_miss = _T_10410; // @[el2_ifu_mem_ctl.scala 809:22]
  assign io_ifu_pmu_ic_hit = _T_10411; // @[el2_ifu_mem_ctl.scala 810:21]
  assign io_ifu_pmu_bus_error = _T_10412; // @[el2_ifu_mem_ctl.scala 811:24]
  assign io_ifu_pmu_bus_busy = _T_10416; // @[el2_ifu_mem_ctl.scala 812:23]
  assign io_ifu_pmu_bus_trxn = _T_10417; // @[el2_ifu_mem_ctl.scala 813:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 142:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 141:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 136:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 140:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 138:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 151:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 144:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 135:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 143:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 152:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 561:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2572; // @[el2_ifu_mem_ctl.scala 562:19]
  assign io_ifu_axi_araddr = _T_2574 & _T_2576; // @[el2_ifu_mem_ctl.scala 563:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 566:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 564:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 567:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 565:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 145:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 568:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 658:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 656:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 660:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 651:20]
  assign io_iccm_ready = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 631:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 338:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3964; // @[el2_ifu_mem_ctl.scala 698:15]
  assign io_ic_rd_en = _T_3956 | _T_3961; // @[el2_ifu_mem_ctl.scala 689:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 345:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 345:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 346:23]
  assign io_ifu_ic_debug_rd_data = _T_1209; // @[el2_ifu_mem_ctl.scala 354:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 816:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 818:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 819:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 817:25]
  assign io_ic_debug_way = _T_10429[1:0]; // @[el2_ifu_mem_ctl.scala 820:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10403; // @[el2_ifu_mem_ctl.scala 804:19]
  assign io_iccm_rw_addr = _T_3110[14:0]; // @[el2_ifu_mem_ctl.scala 662:19]
  assign io_iccm_wren = _T_2679 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 633:16]
  assign io_iccm_rden = _T_2683 | _T_2684; // @[el2_ifu_mem_ctl.scala 634:16]
  assign io_iccm_wr_data = _T_3085 ? _T_3086 : _T_3093; // @[el2_ifu_mem_ctl.scala 639:19]
  assign io_iccm_wr_size = _T_2689 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 636:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 290:15]
  assign io_ic_access_fault_f = _T_2457 & _T_317; // @[el2_ifu_mem_ctl.scala 386:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1271; // @[el2_ifu_mem_ctl.scala 387:29]
  assign io_iccm_rd_ecc_single_err = _T_3901 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 675:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 676:29]
  assign io_ic_error_start = _T_1197 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 348:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 190:24]
  assign io_ic_fetch_val_f = {_T_1279,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 390:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 383:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 380:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 381:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10440; // @[el2_ifu_mem_ctl.scala 827:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2462; // @[el2_ifu_mem_ctl.scala 480:27]
  assign io_iccm_correction_state = _T_2490 ? 1'h0 : _GEN_60; // @[el2_ifu_mem_ctl.scala 515:28 el2_ifu_mem_ctl.scala 528:32 el2_ifu_mem_ctl.scala 535:32 el2_ifu_mem_ctl.scala 542:32]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_5166 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4522 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4518 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4514 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4510 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4506 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4502 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4498 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4494 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4490 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4486 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4482 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4478 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4474 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4470 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4466 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4462 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4458 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4454 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4450 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4446 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4442 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4438 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4434 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4430 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4426 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4422 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4418 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4414 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4410 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4406 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4402 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4398 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4394 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4390 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4386 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4382 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4378 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4374 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4370 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4366 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4362 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4358 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4354 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4350 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4346 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4342 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4338 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4334 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_4330 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_4326 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_4322 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_4318 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_4314 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_4310 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_4306 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_4302 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_4298 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_4294 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4290 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4286 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4282 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4278 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_4274 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_4270 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_4266 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_4262 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4258 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4254 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4250 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4246 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4242 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4238 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4234 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4230 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_4226 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4222 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_4218 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_4214 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_4210 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_4206 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_4202 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_4198 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_4194 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_4190 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_4186 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_4182 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_4178 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_4174 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_4170 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_4166 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_4162 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_4158 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_4154 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_4150 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_4146 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_4142 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_4138 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_4134 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_4130 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_4126 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_4122 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_4118 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_4114 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_4110 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_4106 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_4102 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_4098 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4094 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4090 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4086 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4082 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_4078 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_4074 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_4070 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_4066 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_4062 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_4058 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_4054 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_4050 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_4046 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_4042 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_4038 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_4034 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_4030 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_4026 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_4022 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_4018 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_4014 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_1209 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_10410 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10411 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10412 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10416 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10417 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10440 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_4522 <= 3'h0;
    end else if (_T_4521) begin
      _T_4522 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4518 <= 3'h0;
    end else if (_T_4517) begin
      _T_4518 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4514 <= 3'h0;
    end else if (_T_4513) begin
      _T_4514 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4510 <= 3'h0;
    end else if (_T_4509) begin
      _T_4510 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4506 <= 3'h0;
    end else if (_T_4505) begin
      _T_4506 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4502 <= 3'h0;
    end else if (_T_4501) begin
      _T_4502 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4498 <= 3'h0;
    end else if (_T_4497) begin
      _T_4498 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4494 <= 3'h0;
    end else if (_T_4493) begin
      _T_4494 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4490 <= 3'h0;
    end else if (_T_4489) begin
      _T_4490 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4486 <= 3'h0;
    end else if (_T_4485) begin
      _T_4486 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4482 <= 3'h0;
    end else if (_T_4481) begin
      _T_4482 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4478 <= 3'h0;
    end else if (_T_4477) begin
      _T_4478 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4474 <= 3'h0;
    end else if (_T_4473) begin
      _T_4474 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4470 <= 3'h0;
    end else if (_T_4469) begin
      _T_4470 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4466 <= 3'h0;
    end else if (_T_4465) begin
      _T_4466 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4462 <= 3'h0;
    end else if (_T_4461) begin
      _T_4462 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4458 <= 3'h0;
    end else if (_T_4457) begin
      _T_4458 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4454 <= 3'h0;
    end else if (_T_4453) begin
      _T_4454 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4450 <= 3'h0;
    end else if (_T_4449) begin
      _T_4450 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4446 <= 3'h0;
    end else if (_T_4445) begin
      _T_4446 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4442 <= 3'h0;
    end else if (_T_4441) begin
      _T_4442 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4438 <= 3'h0;
    end else if (_T_4437) begin
      _T_4438 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4434 <= 3'h0;
    end else if (_T_4433) begin
      _T_4434 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4430 <= 3'h0;
    end else if (_T_4429) begin
      _T_4430 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4426 <= 3'h0;
    end else if (_T_4425) begin
      _T_4426 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4422 <= 3'h0;
    end else if (_T_4421) begin
      _T_4422 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4418 <= 3'h0;
    end else if (_T_4417) begin
      _T_4418 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4414 <= 3'h0;
    end else if (_T_4413) begin
      _T_4414 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4410 <= 3'h0;
    end else if (_T_4409) begin
      _T_4410 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4406 <= 3'h0;
    end else if (_T_4405) begin
      _T_4406 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4402 <= 3'h0;
    end else if (_T_4401) begin
      _T_4402 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4398 <= 3'h0;
    end else if (_T_4397) begin
      _T_4398 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4394 <= 3'h0;
    end else if (_T_4393) begin
      _T_4394 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4390 <= 3'h0;
    end else if (_T_4389) begin
      _T_4390 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4386 <= 3'h0;
    end else if (_T_4385) begin
      _T_4386 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4382 <= 3'h0;
    end else if (_T_4381) begin
      _T_4382 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4378 <= 3'h0;
    end else if (_T_4377) begin
      _T_4378 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4374 <= 3'h0;
    end else if (_T_4373) begin
      _T_4374 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4370 <= 3'h0;
    end else if (_T_4369) begin
      _T_4370 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4366 <= 3'h0;
    end else if (_T_4365) begin
      _T_4366 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4362 <= 3'h0;
    end else if (_T_4361) begin
      _T_4362 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4358 <= 3'h0;
    end else if (_T_4357) begin
      _T_4358 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4354 <= 3'h0;
    end else if (_T_4353) begin
      _T_4354 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4350 <= 3'h0;
    end else if (_T_4349) begin
      _T_4350 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4346 <= 3'h0;
    end else if (_T_4345) begin
      _T_4346 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4342 <= 3'h0;
    end else if (_T_4341) begin
      _T_4342 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4338 <= 3'h0;
    end else if (_T_4337) begin
      _T_4338 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4334 <= 3'h0;
    end else if (_T_4333) begin
      _T_4334 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4330 <= 3'h0;
    end else if (_T_4329) begin
      _T_4330 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4326 <= 3'h0;
    end else if (_T_4325) begin
      _T_4326 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4322 <= 3'h0;
    end else if (_T_4321) begin
      _T_4322 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4318 <= 3'h0;
    end else if (_T_4317) begin
      _T_4318 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4314 <= 3'h0;
    end else if (_T_4313) begin
      _T_4314 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4310 <= 3'h0;
    end else if (_T_4309) begin
      _T_4310 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4306 <= 3'h0;
    end else if (_T_4305) begin
      _T_4306 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4302 <= 3'h0;
    end else if (_T_4301) begin
      _T_4302 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4298 <= 3'h0;
    end else if (_T_4297) begin
      _T_4298 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4294 <= 3'h0;
    end else if (_T_4293) begin
      _T_4294 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4290 <= 3'h0;
    end else if (_T_4289) begin
      _T_4290 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4286 <= 3'h0;
    end else if (_T_4285) begin
      _T_4286 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4282 <= 3'h0;
    end else if (_T_4281) begin
      _T_4282 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4278 <= 3'h0;
    end else if (_T_4277) begin
      _T_4278 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4274 <= 3'h0;
    end else if (_T_4273) begin
      _T_4274 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4270 <= 3'h0;
    end else if (_T_4269) begin
      _T_4270 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4266 <= 3'h0;
    end else if (_T_4265) begin
      _T_4266 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4262 <= 3'h0;
    end else if (_T_4261) begin
      _T_4262 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4258 <= 3'h0;
    end else if (_T_4257) begin
      _T_4258 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4254 <= 3'h0;
    end else if (_T_4253) begin
      _T_4254 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4250 <= 3'h0;
    end else if (_T_4249) begin
      _T_4250 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4246 <= 3'h0;
    end else if (_T_4245) begin
      _T_4246 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4242 <= 3'h0;
    end else if (_T_4241) begin
      _T_4242 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4238 <= 3'h0;
    end else if (_T_4237) begin
      _T_4238 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4234 <= 3'h0;
    end else if (_T_4233) begin
      _T_4234 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4230 <= 3'h0;
    end else if (_T_4229) begin
      _T_4230 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4226 <= 3'h0;
    end else if (_T_4225) begin
      _T_4226 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4222 <= 3'h0;
    end else if (_T_4221) begin
      _T_4222 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4218 <= 3'h0;
    end else if (_T_4217) begin
      _T_4218 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4214 <= 3'h0;
    end else if (_T_4213) begin
      _T_4214 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4210 <= 3'h0;
    end else if (_T_4209) begin
      _T_4210 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4206 <= 3'h0;
    end else if (_T_4205) begin
      _T_4206 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4202 <= 3'h0;
    end else if (_T_4201) begin
      _T_4202 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4198 <= 3'h0;
    end else if (_T_4197) begin
      _T_4198 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4194 <= 3'h0;
    end else if (_T_4193) begin
      _T_4194 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4190 <= 3'h0;
    end else if (_T_4189) begin
      _T_4190 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4186 <= 3'h0;
    end else if (_T_4185) begin
      _T_4186 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4182 <= 3'h0;
    end else if (_T_4181) begin
      _T_4182 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4178 <= 3'h0;
    end else if (_T_4177) begin
      _T_4178 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4174 <= 3'h0;
    end else if (_T_4173) begin
      _T_4174 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4170 <= 3'h0;
    end else if (_T_4169) begin
      _T_4170 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4166 <= 3'h0;
    end else if (_T_4165) begin
      _T_4166 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4162 <= 3'h0;
    end else if (_T_4161) begin
      _T_4162 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4158 <= 3'h0;
    end else if (_T_4157) begin
      _T_4158 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4154 <= 3'h0;
    end else if (_T_4153) begin
      _T_4154 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4150 <= 3'h0;
    end else if (_T_4149) begin
      _T_4150 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4146 <= 3'h0;
    end else if (_T_4145) begin
      _T_4146 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4142 <= 3'h0;
    end else if (_T_4141) begin
      _T_4142 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4138 <= 3'h0;
    end else if (_T_4137) begin
      _T_4138 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4134 <= 3'h0;
    end else if (_T_4133) begin
      _T_4134 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4130 <= 3'h0;
    end else if (_T_4129) begin
      _T_4130 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4126 <= 3'h0;
    end else if (_T_4125) begin
      _T_4126 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4122 <= 3'h0;
    end else if (_T_4121) begin
      _T_4122 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4118 <= 3'h0;
    end else if (_T_4117) begin
      _T_4118 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4114 <= 3'h0;
    end else if (_T_4113) begin
      _T_4114 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4110 <= 3'h0;
    end else if (_T_4109) begin
      _T_4110 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4106 <= 3'h0;
    end else if (_T_4105) begin
      _T_4106 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4102 <= 3'h0;
    end else if (_T_4101) begin
      _T_4102 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4098 <= 3'h0;
    end else if (_T_4097) begin
      _T_4098 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4094 <= 3'h0;
    end else if (_T_4093) begin
      _T_4094 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4090 <= 3'h0;
    end else if (_T_4089) begin
      _T_4090 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4086 <= 3'h0;
    end else if (_T_4085) begin
      _T_4086 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4082 <= 3'h0;
    end else if (_T_4081) begin
      _T_4082 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4078 <= 3'h0;
    end else if (_T_4077) begin
      _T_4078 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4074 <= 3'h0;
    end else if (_T_4073) begin
      _T_4074 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4070 <= 3'h0;
    end else if (_T_4069) begin
      _T_4070 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4066 <= 3'h0;
    end else if (_T_4065) begin
      _T_4066 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4062 <= 3'h0;
    end else if (_T_4061) begin
      _T_4062 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4058 <= 3'h0;
    end else if (_T_4057) begin
      _T_4058 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4054 <= 3'h0;
    end else if (_T_4053) begin
      _T_4054 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4050 <= 3'h0;
    end else if (_T_4049) begin
      _T_4050 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4046 <= 3'h0;
    end else if (_T_4045) begin
      _T_4046 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4042 <= 3'h0;
    end else if (_T_4041) begin
      _T_4042 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4038 <= 3'h0;
    end else if (_T_4037) begin
      _T_4038 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4034 <= 3'h0;
    end else if (_T_4033) begin
      _T_4034 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4030 <= 3'h0;
    end else if (_T_4029) begin
      _T_4030 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4026 <= 3'h0;
    end else if (_T_4025) begin
      _T_4026 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4022 <= 3'h0;
    end else if (_T_4021) begin
      _T_4022 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4018 <= 3'h0;
    end else if (_T_4017) begin
      _T_4018 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4014 <= 3'h0;
    end else if (_T_4013) begin
      _T_4014 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_289;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2615) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2611;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5807) begin
      ic_tag_valid_out_1_0 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5824) begin
      ic_tag_valid_out_1_1 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5841) begin
      ic_tag_valid_out_1_2 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5858) begin
      ic_tag_valid_out_1_3 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5875) begin
      ic_tag_valid_out_1_4 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5892) begin
      ic_tag_valid_out_1_5 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5909) begin
      ic_tag_valid_out_1_6 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5926) begin
      ic_tag_valid_out_1_7 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5943) begin
      ic_tag_valid_out_1_8 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5960) begin
      ic_tag_valid_out_1_9 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5977) begin
      ic_tag_valid_out_1_10 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5994) begin
      ic_tag_valid_out_1_11 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_6011) begin
      ic_tag_valid_out_1_12 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_6028) begin
      ic_tag_valid_out_1_13 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_6045) begin
      ic_tag_valid_out_1_14 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_6062) begin
      ic_tag_valid_out_1_15 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_6079) begin
      ic_tag_valid_out_1_16 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_6096) begin
      ic_tag_valid_out_1_17 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6113) begin
      ic_tag_valid_out_1_18 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6130) begin
      ic_tag_valid_out_1_19 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6147) begin
      ic_tag_valid_out_1_20 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6164) begin
      ic_tag_valid_out_1_21 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6181) begin
      ic_tag_valid_out_1_22 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6198) begin
      ic_tag_valid_out_1_23 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6215) begin
      ic_tag_valid_out_1_24 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6232) begin
      ic_tag_valid_out_1_25 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6249) begin
      ic_tag_valid_out_1_26 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6266) begin
      ic_tag_valid_out_1_27 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6283) begin
      ic_tag_valid_out_1_28 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6300) begin
      ic_tag_valid_out_1_29 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6317) begin
      ic_tag_valid_out_1_30 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6334) begin
      ic_tag_valid_out_1_31 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6895) begin
      ic_tag_valid_out_1_32 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6912) begin
      ic_tag_valid_out_1_33 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6929) begin
      ic_tag_valid_out_1_34 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6946) begin
      ic_tag_valid_out_1_35 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6963) begin
      ic_tag_valid_out_1_36 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6980) begin
      ic_tag_valid_out_1_37 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6997) begin
      ic_tag_valid_out_1_38 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_7014) begin
      ic_tag_valid_out_1_39 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_7031) begin
      ic_tag_valid_out_1_40 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_7048) begin
      ic_tag_valid_out_1_41 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_7065) begin
      ic_tag_valid_out_1_42 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_7082) begin
      ic_tag_valid_out_1_43 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_7099) begin
      ic_tag_valid_out_1_44 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_7116) begin
      ic_tag_valid_out_1_45 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_7133) begin
      ic_tag_valid_out_1_46 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_7150) begin
      ic_tag_valid_out_1_47 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7167) begin
      ic_tag_valid_out_1_48 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7184) begin
      ic_tag_valid_out_1_49 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7201) begin
      ic_tag_valid_out_1_50 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7218) begin
      ic_tag_valid_out_1_51 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7235) begin
      ic_tag_valid_out_1_52 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7252) begin
      ic_tag_valid_out_1_53 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7269) begin
      ic_tag_valid_out_1_54 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7286) begin
      ic_tag_valid_out_1_55 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7303) begin
      ic_tag_valid_out_1_56 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7320) begin
      ic_tag_valid_out_1_57 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7337) begin
      ic_tag_valid_out_1_58 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7354) begin
      ic_tag_valid_out_1_59 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7371) begin
      ic_tag_valid_out_1_60 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7388) begin
      ic_tag_valid_out_1_61 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7405) begin
      ic_tag_valid_out_1_62 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7422) begin
      ic_tag_valid_out_1_63 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7983) begin
      ic_tag_valid_out_1_64 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_8000) begin
      ic_tag_valid_out_1_65 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_8017) begin
      ic_tag_valid_out_1_66 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_8034) begin
      ic_tag_valid_out_1_67 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_8051) begin
      ic_tag_valid_out_1_68 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_8068) begin
      ic_tag_valid_out_1_69 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_8085) begin
      ic_tag_valid_out_1_70 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_8102) begin
      ic_tag_valid_out_1_71 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_8119) begin
      ic_tag_valid_out_1_72 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_8136) begin
      ic_tag_valid_out_1_73 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_8153) begin
      ic_tag_valid_out_1_74 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_8170) begin
      ic_tag_valid_out_1_75 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_8187) begin
      ic_tag_valid_out_1_76 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_8204) begin
      ic_tag_valid_out_1_77 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_8221) begin
      ic_tag_valid_out_1_78 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8238) begin
      ic_tag_valid_out_1_79 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8255) begin
      ic_tag_valid_out_1_80 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8272) begin
      ic_tag_valid_out_1_81 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8289) begin
      ic_tag_valid_out_1_82 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8306) begin
      ic_tag_valid_out_1_83 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8323) begin
      ic_tag_valid_out_1_84 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8340) begin
      ic_tag_valid_out_1_85 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8357) begin
      ic_tag_valid_out_1_86 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8374) begin
      ic_tag_valid_out_1_87 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8391) begin
      ic_tag_valid_out_1_88 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8408) begin
      ic_tag_valid_out_1_89 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8425) begin
      ic_tag_valid_out_1_90 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8442) begin
      ic_tag_valid_out_1_91 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8459) begin
      ic_tag_valid_out_1_92 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8476) begin
      ic_tag_valid_out_1_93 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8493) begin
      ic_tag_valid_out_1_94 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8510) begin
      ic_tag_valid_out_1_95 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_9071) begin
      ic_tag_valid_out_1_96 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_9088) begin
      ic_tag_valid_out_1_97 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_9105) begin
      ic_tag_valid_out_1_98 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_9122) begin
      ic_tag_valid_out_1_99 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_9139) begin
      ic_tag_valid_out_1_100 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_9156) begin
      ic_tag_valid_out_1_101 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_9173) begin
      ic_tag_valid_out_1_102 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_9190) begin
      ic_tag_valid_out_1_103 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_9207) begin
      ic_tag_valid_out_1_104 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_9224) begin
      ic_tag_valid_out_1_105 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_9241) begin
      ic_tag_valid_out_1_106 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_9258) begin
      ic_tag_valid_out_1_107 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_9275) begin
      ic_tag_valid_out_1_108 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9292) begin
      ic_tag_valid_out_1_109 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9309) begin
      ic_tag_valid_out_1_110 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9326) begin
      ic_tag_valid_out_1_111 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9343) begin
      ic_tag_valid_out_1_112 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9360) begin
      ic_tag_valid_out_1_113 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9377) begin
      ic_tag_valid_out_1_114 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9394) begin
      ic_tag_valid_out_1_115 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9411) begin
      ic_tag_valid_out_1_116 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9428) begin
      ic_tag_valid_out_1_117 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9445) begin
      ic_tag_valid_out_1_118 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9462) begin
      ic_tag_valid_out_1_119 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9479) begin
      ic_tag_valid_out_1_120 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9496) begin
      ic_tag_valid_out_1_121 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9513) begin
      ic_tag_valid_out_1_122 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9530) begin
      ic_tag_valid_out_1_123 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9547) begin
      ic_tag_valid_out_1_124 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9564) begin
      ic_tag_valid_out_1_125 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9581) begin
      ic_tag_valid_out_1_126 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9598) begin
      ic_tag_valid_out_1_127 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5263) begin
      ic_tag_valid_out_0_0 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5280) begin
      ic_tag_valid_out_0_1 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5297) begin
      ic_tag_valid_out_0_2 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5314) begin
      ic_tag_valid_out_0_3 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5331) begin
      ic_tag_valid_out_0_4 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5348) begin
      ic_tag_valid_out_0_5 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5365) begin
      ic_tag_valid_out_0_6 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5382) begin
      ic_tag_valid_out_0_7 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5399) begin
      ic_tag_valid_out_0_8 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5416) begin
      ic_tag_valid_out_0_9 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5433) begin
      ic_tag_valid_out_0_10 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5450) begin
      ic_tag_valid_out_0_11 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5467) begin
      ic_tag_valid_out_0_12 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5484) begin
      ic_tag_valid_out_0_13 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5501) begin
      ic_tag_valid_out_0_14 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5518) begin
      ic_tag_valid_out_0_15 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5535) begin
      ic_tag_valid_out_0_16 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5552) begin
      ic_tag_valid_out_0_17 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5569) begin
      ic_tag_valid_out_0_18 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5586) begin
      ic_tag_valid_out_0_19 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5603) begin
      ic_tag_valid_out_0_20 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5620) begin
      ic_tag_valid_out_0_21 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5637) begin
      ic_tag_valid_out_0_22 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5654) begin
      ic_tag_valid_out_0_23 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5671) begin
      ic_tag_valid_out_0_24 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5688) begin
      ic_tag_valid_out_0_25 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5705) begin
      ic_tag_valid_out_0_26 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5722) begin
      ic_tag_valid_out_0_27 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5739) begin
      ic_tag_valid_out_0_28 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5756) begin
      ic_tag_valid_out_0_29 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5773) begin
      ic_tag_valid_out_0_30 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5790) begin
      ic_tag_valid_out_0_31 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6351) begin
      ic_tag_valid_out_0_32 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6368) begin
      ic_tag_valid_out_0_33 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6385) begin
      ic_tag_valid_out_0_34 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6402) begin
      ic_tag_valid_out_0_35 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6419) begin
      ic_tag_valid_out_0_36 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6436) begin
      ic_tag_valid_out_0_37 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6453) begin
      ic_tag_valid_out_0_38 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6470) begin
      ic_tag_valid_out_0_39 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6487) begin
      ic_tag_valid_out_0_40 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6504) begin
      ic_tag_valid_out_0_41 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6521) begin
      ic_tag_valid_out_0_42 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6538) begin
      ic_tag_valid_out_0_43 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6555) begin
      ic_tag_valid_out_0_44 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6572) begin
      ic_tag_valid_out_0_45 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6589) begin
      ic_tag_valid_out_0_46 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6606) begin
      ic_tag_valid_out_0_47 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6623) begin
      ic_tag_valid_out_0_48 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6640) begin
      ic_tag_valid_out_0_49 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6657) begin
      ic_tag_valid_out_0_50 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6674) begin
      ic_tag_valid_out_0_51 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6691) begin
      ic_tag_valid_out_0_52 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6708) begin
      ic_tag_valid_out_0_53 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6725) begin
      ic_tag_valid_out_0_54 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6742) begin
      ic_tag_valid_out_0_55 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6759) begin
      ic_tag_valid_out_0_56 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6776) begin
      ic_tag_valid_out_0_57 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6793) begin
      ic_tag_valid_out_0_58 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6810) begin
      ic_tag_valid_out_0_59 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6827) begin
      ic_tag_valid_out_0_60 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6844) begin
      ic_tag_valid_out_0_61 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6861) begin
      ic_tag_valid_out_0_62 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6878) begin
      ic_tag_valid_out_0_63 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7439) begin
      ic_tag_valid_out_0_64 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7456) begin
      ic_tag_valid_out_0_65 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7473) begin
      ic_tag_valid_out_0_66 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7490) begin
      ic_tag_valid_out_0_67 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7507) begin
      ic_tag_valid_out_0_68 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7524) begin
      ic_tag_valid_out_0_69 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7541) begin
      ic_tag_valid_out_0_70 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7558) begin
      ic_tag_valid_out_0_71 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7575) begin
      ic_tag_valid_out_0_72 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7592) begin
      ic_tag_valid_out_0_73 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7609) begin
      ic_tag_valid_out_0_74 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7626) begin
      ic_tag_valid_out_0_75 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7643) begin
      ic_tag_valid_out_0_76 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7660) begin
      ic_tag_valid_out_0_77 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7677) begin
      ic_tag_valid_out_0_78 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7694) begin
      ic_tag_valid_out_0_79 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7711) begin
      ic_tag_valid_out_0_80 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7728) begin
      ic_tag_valid_out_0_81 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7745) begin
      ic_tag_valid_out_0_82 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7762) begin
      ic_tag_valid_out_0_83 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7779) begin
      ic_tag_valid_out_0_84 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7796) begin
      ic_tag_valid_out_0_85 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7813) begin
      ic_tag_valid_out_0_86 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7830) begin
      ic_tag_valid_out_0_87 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7847) begin
      ic_tag_valid_out_0_88 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7864) begin
      ic_tag_valid_out_0_89 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7881) begin
      ic_tag_valid_out_0_90 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7898) begin
      ic_tag_valid_out_0_91 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7915) begin
      ic_tag_valid_out_0_92 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7932) begin
      ic_tag_valid_out_0_93 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7949) begin
      ic_tag_valid_out_0_94 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7966) begin
      ic_tag_valid_out_0_95 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8527) begin
      ic_tag_valid_out_0_96 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8544) begin
      ic_tag_valid_out_0_97 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8561) begin
      ic_tag_valid_out_0_98 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8578) begin
      ic_tag_valid_out_0_99 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8595) begin
      ic_tag_valid_out_0_100 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8612) begin
      ic_tag_valid_out_0_101 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8629) begin
      ic_tag_valid_out_0_102 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8646) begin
      ic_tag_valid_out_0_103 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8663) begin
      ic_tag_valid_out_0_104 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8680) begin
      ic_tag_valid_out_0_105 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8697) begin
      ic_tag_valid_out_0_106 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8714) begin
      ic_tag_valid_out_0_107 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8731) begin
      ic_tag_valid_out_0_108 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8748) begin
      ic_tag_valid_out_0_109 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8765) begin
      ic_tag_valid_out_0_110 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8782) begin
      ic_tag_valid_out_0_111 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8799) begin
      ic_tag_valid_out_0_112 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8816) begin
      ic_tag_valid_out_0_113 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8833) begin
      ic_tag_valid_out_0_114 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8850) begin
      ic_tag_valid_out_0_115 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8867) begin
      ic_tag_valid_out_0_116 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8884) begin
      ic_tag_valid_out_0_117 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8901) begin
      ic_tag_valid_out_0_118 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8918) begin
      ic_tag_valid_out_0_119 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8935) begin
      ic_tag_valid_out_0_120 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8952) begin
      ic_tag_valid_out_0_121 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8969) begin
      ic_tag_valid_out_0_122 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8986) begin
      ic_tag_valid_out_0_123 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_9003) begin
      ic_tag_valid_out_0_124 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_9020) begin
      ic_tag_valid_out_0_125 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_9037) begin
      ic_tag_valid_out_0_126 <= _T_5253;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_9054) begin
      ic_tag_valid_out_0_127 <= _T_5253;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1209 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_1209 <= {{5'd0}, _T_1208};
      end else begin
        _T_1209 <= io_ic_debug_rd_data;
      end
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2564) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2639) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2683;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2465) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2467) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2477) begin
        perr_state <= 3'h0;
      end else if (_T_2480) begin
        if (_T_2482) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2486) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2490) begin
        err_stop_state <= 2'h1;
      end else if (_T_2495) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (_T_2518) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2522) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2539) begin
        if (_T_2543) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1368;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_5166 <= 7'h0;
    end else if (_T_3987) begin
      _T_5166 <= io_ic_debug_addr[9:3];
    end else begin
      _T_5166 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1408;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3922;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3097;
    end else begin
      iccm_dma_rdata <= _T_3098;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3918;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3987) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3990) begin
      way_status_new_ff <= _T_3994;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3990) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10440 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10440 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10410 <= 1'h0;
    end else begin
      _T_10410 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10411 <= 1'h0;
    end else begin
      _T_10411 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10412 <= 1'h0;
    end else begin
      _T_10412 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10416 <= 1'h0;
    end else begin
      _T_10416 <= _T_10415;
    end
    if (reset) begin
      _T_10417 <= 1'h0;
    end else begin
      _T_10417 <= bus_cmd_sent;
    end
  end
endmodule
