module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[el2_lib.scala 408:26]
  wire  clkhdr_CK; // @[el2_lib.scala 408:26]
  wire  clkhdr_EN; // @[el2_lib.scala 408:26]
  wire  clkhdr_SE; // @[el2_lib.scala 408:26]
  TEC_RV_ICG clkhdr ( // @[el2_lib.scala 408:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[el2_lib.scala 409:14]
  assign clkhdr_CK = io_clk; // @[el2_lib.scala 410:18]
  assign clkhdr_EN = io_en; // @[el2_lib.scala 411:18]
  assign clkhdr_SE = io_scan_mode; // @[el2_lib.scala 412:18]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  input         io_ifu_axi_arready,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  input         io_ifu_axi_rvalid,
  output        io_ifu_axi_rready,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [95:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [63:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_1_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_2_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_3_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_4_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_5_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_6_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_7_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_8_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_9_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_10_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_11_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_12_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_13_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_14_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_15_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_16_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_17_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_18_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_19_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_20_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_21_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_22_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_23_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_24_io_scan_mode; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_l1clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_clk; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_en; // @[el2_lib.scala 417:22]
  wire  rvclkhdr_25_io_scan_mode; // @[el2_lib.scala 417:22]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 234:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 367:36]
  wire  _T_309 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 368:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_309; // @[el2_ifu_mem_ctl.scala 368:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 235:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 300:30]
  wire  _T_1 = _T | miss_pending; // @[el2_ifu_mem_ctl.scala 235:71]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 236:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 355:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 705:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 705:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_309}; // @[el2_ifu_mem_ctl.scala 708:91]
  wire [1:0] _T_3059 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 708:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 369:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 322:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 708:113]
  wire [1:0] _T_3060 = _T_3059 & _GEN_465; // @[el2_ifu_mem_ctl.scala 708:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 694:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 708:130]
  wire [1:0] _T_3061 = _T_3060 | _GEN_466; // @[el2_ifu_mem_ctl.scala 708:130]
  wire  _T_3062 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 708:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_3062}; // @[el2_ifu_mem_ctl.scala 708:152]
  wire [1:0] _T_3063 = _T_3061 & _GEN_467; // @[el2_ifu_mem_ctl.scala 708:152]
  wire [1:0] _T_3052 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 708:91]
  wire [1:0] _T_3053 = _T_3052 & _GEN_465; // @[el2_ifu_mem_ctl.scala 708:113]
  wire [1:0] _T_3054 = _T_3053 | _GEN_466; // @[el2_ifu_mem_ctl.scala 708:130]
  wire [1:0] _T_3056 = _T_3054 & _GEN_467; // @[el2_ifu_mem_ctl.scala 708:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3063,_T_3056}; // @[Cat.scala 29:58]
  wire  _T_3163 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3164 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3165 = _T_3163 ^ _T_3164; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3173 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3174 = ^_T_3173; // @[el2_lib.scala 301:83]
  wire  _T_3175 = io_iccm_rd_data_ecc[37] ^ _T_3174; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3182 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3190 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3182}; // @[el2_lib.scala 301:103]
  wire  _T_3191 = ^_T_3190; // @[el2_lib.scala 301:110]
  wire  _T_3192 = io_iccm_rd_data_ecc[36] ^ _T_3191; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3199 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3207 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3199}; // @[el2_lib.scala 301:130]
  wire  _T_3208 = ^_T_3207; // @[el2_lib.scala 301:137]
  wire  _T_3209 = io_iccm_rd_data_ecc[35] ^ _T_3208; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3218 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3227 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3218}; // @[el2_lib.scala 301:157]
  wire  _T_3228 = ^_T_3227; // @[el2_lib.scala 301:164]
  wire  _T_3229 = io_iccm_rd_data_ecc[34] ^ _T_3228; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3238 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3247 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3238}; // @[el2_lib.scala 301:184]
  wire  _T_3248 = ^_T_3247; // @[el2_lib.scala 301:191]
  wire  _T_3249 = io_iccm_rd_data_ecc[33] ^ _T_3248; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3258 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3267 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3258}; // @[el2_lib.scala 301:211]
  wire  _T_3268 = ^_T_3267; // @[el2_lib.scala 301:218]
  wire  _T_3269 = io_iccm_rd_data_ecc[32] ^ _T_3268; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3275 = {_T_3165,_T_3175,_T_3192,_T_3209,_T_3229,_T_3249,_T_3269}; // @[Cat.scala 29:58]
  wire  _T_3276 = _T_3275 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3277 = iccm_ecc_word_enable[0] & _T_3276; // @[el2_lib.scala 302:32]
  wire  _T_3279 = _T_3277 & _T_3275[6]; // @[el2_lib.scala 302:53]
  wire  _T_3548 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3549 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3550 = _T_3548 ^ _T_3549; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3558 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3559 = ^_T_3558; // @[el2_lib.scala 301:83]
  wire  _T_3560 = io_iccm_rd_data_ecc[76] ^ _T_3559; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3567 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3575 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3567}; // @[el2_lib.scala 301:103]
  wire  _T_3576 = ^_T_3575; // @[el2_lib.scala 301:110]
  wire  _T_3577 = io_iccm_rd_data_ecc[75] ^ _T_3576; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3584 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3592 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3584}; // @[el2_lib.scala 301:130]
  wire  _T_3593 = ^_T_3592; // @[el2_lib.scala 301:137]
  wire  _T_3594 = io_iccm_rd_data_ecc[74] ^ _T_3593; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3603 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3612 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3603}; // @[el2_lib.scala 301:157]
  wire  _T_3613 = ^_T_3612; // @[el2_lib.scala 301:164]
  wire  _T_3614 = io_iccm_rd_data_ecc[73] ^ _T_3613; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3623 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3632 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3623}; // @[el2_lib.scala 301:184]
  wire  _T_3633 = ^_T_3632; // @[el2_lib.scala 301:191]
  wire  _T_3634 = io_iccm_rd_data_ecc[72] ^ _T_3633; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3643 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3652 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3643}; // @[el2_lib.scala 301:211]
  wire  _T_3653 = ^_T_3652; // @[el2_lib.scala 301:218]
  wire  _T_3654 = io_iccm_rd_data_ecc[71] ^ _T_3653; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3660 = {_T_3550,_T_3560,_T_3577,_T_3594,_T_3614,_T_3634,_T_3654}; // @[Cat.scala 29:58]
  wire  _T_3661 = _T_3660 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3662 = iccm_ecc_word_enable[1] & _T_3661; // @[el2_lib.scala 302:32]
  wire  _T_3664 = _T_3662 & _T_3660[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3279,_T_3664}; // @[Cat.scala 29:58]
  wire  _T_4 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 239:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 672:51]
  wire  _T_7 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 240:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_8 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 241:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 520:34]
  wire  _T_9 = iccm_correct_ecc | _T_8; // @[el2_ifu_mem_ctl.scala 241:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_10 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 241:90]
  wire  _T_11 = _T_9 | _T_10; // @[el2_ifu_mem_ctl.scala 241:72]
  wire  _T_2430 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2435 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2455 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 568:48]
  wire  two_byte_instr = io_ic_rd_data[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 436:39]
  wire  _T_2457 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 568:79]
  wire  _T_2458 = _T_2455 | _T_2457; // @[el2_ifu_mem_ctl.scala 568:56]
  wire  _T_2459 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 568:122]
  wire  _T_2460 = ~_T_2459; // @[el2_ifu_mem_ctl.scala 568:101]
  wire  _T_2461 = _T_2458 & _T_2460; // @[el2_ifu_mem_ctl.scala 568:99]
  wire  _T_2462 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2476 = io_ifu_fetch_val[0] & _T_309; // @[el2_ifu_mem_ctl.scala 575:45]
  wire  _T_2477 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 575:69]
  wire  _T_2478 = _T_2476 & _T_2477; // @[el2_ifu_mem_ctl.scala 575:67]
  wire  _T_2479 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_2462 ? _T_2478 : _T_2479; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2435 ? _T_2461 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2430 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_12 = _T_11 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 241:112]
  wire  _T_14 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 242:44]
  wire  _T_15 = _T_14 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 242:65]
  wire  _T_219 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 330:37]
  wire  _T_220 = ~_T_219; // @[el2_ifu_mem_ctl.scala 330:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 740:53]
  wire  _T_221 = _T_220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 330:41]
  wire  _T_199 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 321:48]
  wire  _T_200 = ifc_fetch_req_f & _T_199; // @[el2_ifu_mem_ctl.scala 321:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 371:42]
  wire  _T_201 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 321:69]
  wire  fetch_req_icache_f = _T_200 & _T_201; // @[el2_ifu_mem_ctl.scala 321:67]
  wire  _T_222 = _T_221 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 330:59]
  wire  _T_223 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 330:82]
  wire  _T_224 = _T_222 & _T_223; // @[el2_ifu_mem_ctl.scala 330:80]
  wire  ic_act_miss_f = _T_224 & _T_201; // @[el2_ifu_mem_ctl.scala 330:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 588:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 629:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 656:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 357:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 637:56]
  wire  _T_2579 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 654:69]
  wire  _T_2580 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 654:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2579 : _T_2580; // @[el2_ifu_mem_ctl.scala 654:28]
  wire  _T_2526 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 633:68]
  wire  _T_2527 = ic_act_miss_f | _T_2526; // @[el2_ifu_mem_ctl.scala 633:48]
  wire  bus_reset_data_beat_cnt = _T_2527 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 633:91]
  wire  _T_2523 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 632:50]
  wire  _T_2524 = bus_ifu_wr_en_ff & _T_2523; // @[el2_ifu_mem_ctl.scala 632:48]
  wire  _T_2525 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 632:72]
  wire  bus_inc_data_beat_cnt = _T_2524 & _T_2525; // @[el2_ifu_mem_ctl.scala 632:70]
  wire [2:0] _T_2531 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 636:115]
  wire [2:0] _T_2533 = bus_inc_data_beat_cnt ? _T_2531 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2528 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 634:32]
  wire  _T_2529 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 634:57]
  wire  bus_hold_data_beat_cnt = _T_2528 & _T_2529; // @[el2_ifu_mem_ctl.scala 634:55]
  wire [2:0] _T_2534 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2533 | _T_2534; // @[Mux.scala 27:72]
  wire  _T_16 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 242:111]
  wire  _T_17 = _T_15 & _T_16; // @[el2_ifu_mem_ctl.scala 242:85]
  wire  _T_18 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 243:39]
  wire  _T_26 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_28 = ic_act_miss_f & _T_309; // @[el2_ifu_mem_ctl.scala 249:43]
  wire [2:0] _T_30 = _T_28 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 249:27]
  wire  _T_33 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 472:45]
  wire  _T_2098 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 493:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 449:60]
  wire  _T_2129 = _T_2098 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2102 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 493:127]
  wire  _T_2130 = _T_2102 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2137 = _T_2129 | _T_2130; // @[Mux.scala 27:72]
  wire  _T_2106 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 493:127]
  wire  _T_2131 = _T_2106 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2138 = _T_2137 | _T_2131; // @[Mux.scala 27:72]
  wire  _T_2110 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 493:127]
  wire  _T_2132 = _T_2110 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2139 = _T_2138 | _T_2132; // @[Mux.scala 27:72]
  wire  _T_2114 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 493:127]
  wire  _T_2133 = _T_2114 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2140 = _T_2139 | _T_2133; // @[Mux.scala 27:72]
  wire  _T_2118 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 493:127]
  wire  _T_2134 = _T_2118 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2141 = _T_2140 | _T_2134; // @[Mux.scala 27:72]
  wire  _T_2122 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 493:127]
  wire  _T_2135 = _T_2122 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2142 = _T_2141 | _T_2135; // @[Mux.scala 27:72]
  wire  _T_2126 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 493:127]
  wire  _T_2136 = _T_2126 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2142 | _T_2136; // @[Mux.scala 27:72]
  wire  _T_2184 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 495:69]
  wire  _T_2185 = ic_miss_buff_data_valid_bypass_index & _T_2184; // @[el2_ifu_mem_ctl.scala 495:67]
  wire  _T_2187 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 495:91]
  wire  _T_2188 = _T_2185 & _T_2187; // @[el2_ifu_mem_ctl.scala 495:89]
  wire  _T_2193 = _T_2185 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 496:65]
  wire  _T_2194 = _T_2188 | _T_2193; // @[el2_ifu_mem_ctl.scala 495:112]
  wire  _T_2196 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 497:43]
  wire  _T_2199 = _T_2196 & _T_2187; // @[el2_ifu_mem_ctl.scala 497:65]
  wire  _T_2200 = _T_2194 | _T_2199; // @[el2_ifu_mem_ctl.scala 496:88]
  wire  _T_2204 = _T_2196 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 498:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 475:75]
  wire  _T_2144 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2168 = _T_2144 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2147 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2169 = _T_2147 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2176 = _T_2168 | _T_2169; // @[Mux.scala 27:72]
  wire  _T_2150 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2170 = _T_2150 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2177 = _T_2176 | _T_2170; // @[Mux.scala 27:72]
  wire  _T_2153 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2171 = _T_2153 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2178 = _T_2177 | _T_2171; // @[Mux.scala 27:72]
  wire  _T_2156 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2172 = _T_2156 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2179 = _T_2178 | _T_2172; // @[Mux.scala 27:72]
  wire  _T_2159 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2173 = _T_2159 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2180 = _T_2179 | _T_2173; // @[Mux.scala 27:72]
  wire  _T_2162 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2174 = _T_2162 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2181 = _T_2180 | _T_2174; // @[Mux.scala 27:72]
  wire  _T_2165 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 494:110]
  wire  _T_2175 = _T_2165 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2181 | _T_2175; // @[Mux.scala 27:72]
  wire  _T_2205 = _T_2204 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 498:87]
  wire  _T_2206 = _T_2200 | _T_2205; // @[el2_ifu_mem_ctl.scala 497:88]
  wire  _T_2216 = _T_2188 & _T_2126; // @[el2_ifu_mem_ctl.scala 499:87]
  wire  miss_buff_hit_unq_f = _T_2206 | _T_2216; // @[el2_ifu_mem_ctl.scala 498:131]
  wire  _T_2231 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 504:55]
  wire  _T_2232 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 504:87]
  wire  _T_2233 = _T_2231 | _T_2232; // @[el2_ifu_mem_ctl.scala 504:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2233; // @[el2_ifu_mem_ctl.scala 504:41]
  wire  _T_2217 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 501:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 358:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 492:51]
  wire  _T_2218 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 501:68]
  wire  _T_2219 = miss_buff_hit_unq_f & _T_2218; // @[el2_ifu_mem_ctl.scala 501:66]
  wire  stream_hit_f = _T_2217 & _T_2219; // @[el2_ifu_mem_ctl.scala 501:43]
  wire  _T_207 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 325:35]
  wire  _T_208 = _T_207 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 325:52]
  wire  ic_byp_hit_f = _T_208 & miss_pending; // @[el2_ifu_mem_ctl.scala 325:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 639:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 666:35]
  wire  _T_34 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 252:112]
  wire  _T_35 = last_data_recieved_ff | _T_34; // @[el2_ifu_mem_ctl.scala 252:92]
  wire  _T_36 = ic_byp_hit_f & _T_35; // @[el2_ifu_mem_ctl.scala 252:66]
  wire  _T_37 = _T_36 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 252:126]
  wire  _T_38 = io_dec_tlu_force_halt | _T_37; // @[el2_ifu_mem_ctl.scala 252:51]
  wire  _T_40 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 253:30]
  wire  _T_41 = ic_byp_hit_f & _T_40; // @[el2_ifu_mem_ctl.scala 253:27]
  wire  _T_42 = _T_41 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 253:53]
  wire  _T_44 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 254:16]
  wire  _T_46 = _T_44 & _T_309; // @[el2_ifu_mem_ctl.scala 254:30]
  wire  _T_48 = _T_46 & _T_34; // @[el2_ifu_mem_ctl.scala 254:52]
  wire  _T_49 = _T_48 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 254:85]
  wire  _T_52 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 255:51]
  wire  _T_53 = _T_34 & _T_52; // @[el2_ifu_mem_ctl.scala 255:49]
  wire  _T_55 = ic_byp_hit_f | bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 256:34]
  wire  _T_57 = _T_55 & _T_309; // @[el2_ifu_mem_ctl.scala 256:54]
  wire  _T_59 = ~_T_34; // @[el2_ifu_mem_ctl.scala 256:78]
  wire  _T_60 = _T_57 & _T_59; // @[el2_ifu_mem_ctl.scala 256:76]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 245:52]
  wire  _T_61 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 256:112]
  wire  _T_62 = _T_60 & _T_61; // @[el2_ifu_mem_ctl.scala 256:110]
  wire  _T_64 = _T_62 & _T_52; // @[el2_ifu_mem_ctl.scala 256:134]
  wire  _T_72 = _T_48 & _T_52; // @[el2_ifu_mem_ctl.scala 257:100]
  wire  _T_74 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 258:44]
  wire  _T_77 = _T_74 & _T_59; // @[el2_ifu_mem_ctl.scala 258:68]
  wire [2:0] _T_79 = _T_77 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 258:22]
  wire [2:0] _T_80 = _T_72 ? 3'h0 : _T_79; // @[el2_ifu_mem_ctl.scala 257:20]
  wire [2:0] _T_81 = _T_64 ? 3'h6 : _T_80; // @[el2_ifu_mem_ctl.scala 256:18]
  wire [2:0] _T_82 = _T_53 ? 3'h0 : _T_81; // @[el2_ifu_mem_ctl.scala 255:16]
  wire [2:0] _T_83 = _T_49 ? 3'h1 : _T_82; // @[el2_ifu_mem_ctl.scala 254:14]
  wire [2:0] _T_84 = _T_42 ? 3'h3 : _T_83; // @[el2_ifu_mem_ctl.scala 253:12]
  wire [2:0] _T_85 = _T_38 ? 3'h0 : _T_84; // @[el2_ifu_mem_ctl.scala 252:27]
  wire  _T_94 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_98 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2228 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 503:60]
  wire  _T_2229 = _T_2228 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 503:92]
  wire  stream_eol_f = _T_2229 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 503:110]
  wire  _T_100 = _T_74 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 266:72]
  wire  _T_103 = _T_100 & _T_59; // @[el2_ifu_mem_ctl.scala 266:87]
  wire  _T_105 = _T_103 & _T_2525; // @[el2_ifu_mem_ctl.scala 266:122]
  wire [2:0] _T_107 = _T_105 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 266:27]
  wire  _T_113 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_116 = io_exu_flush_final & _T_59; // @[el2_ifu_mem_ctl.scala 270:48]
  wire  _T_118 = _T_116 & _T_2525; // @[el2_ifu_mem_ctl.scala 270:82]
  wire [2:0] _T_120 = _T_118 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 270:27]
  wire  _T_124 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_228 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 331:28]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 331:42]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 331:60]
  wire  _T_231 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 331:94]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 331:81]
  wire  _T_235 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 332:39]
  wire  _T_236 = _T_232 & _T_235; // @[el2_ifu_mem_ctl.scala 331:111]
  wire  _T_238 = _T_236 & _T_52; // @[el2_ifu_mem_ctl.scala 332:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 385:51]
  wire  _T_239 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 332:116]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 332:114]
  wire  ic_miss_under_miss_f = _T_240 & _T_201; // @[el2_ifu_mem_ctl.scala 332:132]
  wire  _T_127 = ic_miss_under_miss_f & _T_59; // @[el2_ifu_mem_ctl.scala 274:50]
  wire  _T_129 = _T_127 & _T_2525; // @[el2_ifu_mem_ctl.scala 274:84]
  wire  _T_248 = _T_222 & _T_231; // @[el2_ifu_mem_ctl.scala 333:85]
  wire  _T_251 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 334:39]
  wire  _T_252 = _T_251 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 334:91]
  wire  ic_ignore_2nd_miss_f = _T_248 & _T_252; // @[el2_ifu_mem_ctl.scala 333:117]
  wire  _T_133 = ic_ignore_2nd_miss_f & _T_59; // @[el2_ifu_mem_ctl.scala 275:35]
  wire  _T_135 = _T_133 & _T_2525; // @[el2_ifu_mem_ctl.scala 275:69]
  wire [2:0] _T_137 = _T_135 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 275:12]
  wire [2:0] _T_138 = _T_129 ? 3'h5 : _T_137; // @[el2_ifu_mem_ctl.scala 274:27]
  wire  _T_143 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_146 = _T_34 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 280:12]
  wire [2:0] _T_147 = io_exu_flush_final ? _T_146 : 3'h1; // @[el2_ifu_mem_ctl.scala 279:62]
  wire [2:0] _T_148 = io_dec_tlu_force_halt ? 3'h0 : _T_147; // @[el2_ifu_mem_ctl.scala 279:27]
  wire  _T_152 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_156 = io_exu_flush_final ? _T_146 : 3'h0; // @[el2_ifu_mem_ctl.scala 284:62]
  wire [2:0] _T_157 = io_dec_tlu_force_halt ? 3'h0 : _T_156; // @[el2_ifu_mem_ctl.scala 284:27]
  wire [2:0] _GEN_0 = _T_152 ? _T_157 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_143 ? _T_148 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_124 ? _T_138 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_113 ? _T_120 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_98 ? _T_107 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_94 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_33 ? _T_85 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_26 ? _T_30 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_19 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 243:71]
  wire  _T_20 = _T_18 | _T_19; // @[el2_ifu_mem_ctl.scala 243:55]
  wire  _T_21 = uncacheable_miss_ff >> _T_20; // @[el2_ifu_mem_ctl.scala 243:26]
  wire  _T_23 = ~_T_21; // @[el2_ifu_mem_ctl.scala 243:5]
  wire  _T_24 = _T_17 & _T_23; // @[el2_ifu_mem_ctl.scala 242:116]
  wire  scnd_miss_req_in = _T_24 & _T_309; // @[el2_ifu_mem_ctl.scala 243:89]
  wire  _T_32 = ic_act_miss_f & _T_2525; // @[el2_ifu_mem_ctl.scala 250:38]
  wire  _T_86 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 259:46]
  wire  _T_87 = _T_86 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 259:67]
  wire  _T_88 = _T_87 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 259:82]
  wire  _T_90 = _T_88 | _T_34; // @[el2_ifu_mem_ctl.scala 259:105]
  wire  _T_92 = bus_ifu_wr_en_ff & _T_52; // @[el2_ifu_mem_ctl.scala 259:158]
  wire  _T_93 = _T_90 | _T_92; // @[el2_ifu_mem_ctl.scala 259:138]
  wire  _T_95 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 263:43]
  wire  _T_96 = _T_95 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 263:59]
  wire  _T_97 = _T_96 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 263:74]
  wire  _T_111 = _T_100 | _T_34; // @[el2_ifu_mem_ctl.scala 267:84]
  wire  _T_112 = _T_111 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 267:118]
  wire  _T_122 = io_exu_flush_final | _T_34; // @[el2_ifu_mem_ctl.scala 271:43]
  wire  _T_123 = _T_122 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 271:76]
  wire  _T_140 = _T_34 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 276:55]
  wire  _T_141 = _T_140 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 276:78]
  wire  _T_142 = _T_141 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 276:101]
  wire  _T_150 = _T_34 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 281:55]
  wire  _T_151 = _T_150 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 281:76]
  wire  _GEN_1 = _T_152 & _T_151; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_143 ? _T_151 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_124 ? _T_142 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_113 ? _T_123 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_98 ? _T_112 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_94 ? _T_97 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_33 ? _T_93 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_26 ? _T_32 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_166 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 301:95]
  wire  _T_167 = _T_2231 & _T_166; // @[el2_ifu_mem_ctl.scala 301:93]
  wire  crit_wd_byp_ok_ff = _T_2232 | _T_167; // @[el2_ifu_mem_ctl.scala 301:58]
  wire  _T_170 = miss_pending & _T_59; // @[el2_ifu_mem_ctl.scala 302:36]
  wire  _T_172 = _T_2231 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 302:106]
  wire  _T_173 = ~_T_172; // @[el2_ifu_mem_ctl.scala 302:72]
  wire  _T_174 = _T_170 & _T_173; // @[el2_ifu_mem_ctl.scala 302:70]
  wire  _T_176 = _T_2231 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 303:57]
  wire  _T_177 = ~_T_176; // @[el2_ifu_mem_ctl.scala 303:23]
  wire  _T_178 = _T_174 & _T_177; // @[el2_ifu_mem_ctl.scala 302:128]
  wire  _T_179 = _T_178 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 303:77]
  wire  _T_180 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 304:36]
  wire  _T_181 = miss_pending & _T_180; // @[el2_ifu_mem_ctl.scala 304:19]
  wire  sel_hold_imb = _T_179 | _T_181; // @[el2_ifu_mem_ctl.scala 303:93]
  wire  _T_183 = _T_18 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 306:57]
  wire  sel_hold_imb_scnd = _T_183 & _T_166; // @[el2_ifu_mem_ctl.scala 306:81]
  reg [6:0] _T_4976; // @[el2_ifu_mem_ctl.scala 770:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_4976[5:0]; // @[el2_ifu_mem_ctl.scala 769:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 766:121]
  wire  _T_4841 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4843 = _T_4841 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4332; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_4332[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4844 = _T_4843 & _GEN_473; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4837 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4839 = _T_4837 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4329; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_4329[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4840 = _T_4839 & _GEN_475; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4833 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4835 = _T_4833 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4326; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_4326[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4836 = _T_4835 & _GEN_477; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4829 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4831 = _T_4829 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4323; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_4323[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4832 = _T_4831 & _GEN_479; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4825 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4827 = _T_4825 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4320; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_4320[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4828 = _T_4827 & _GEN_481; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4821 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4823 = _T_4821 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4317; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_4317[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4824 = _T_4823 & _GEN_483; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4817 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4819 = _T_4817 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4314; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_4314[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4820 = _T_4819 & _GEN_485; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4813 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4815 = _T_4813 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4311; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_4311[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4816 = _T_4815 & _GEN_487; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4809 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4811 = _T_4809 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4308; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_4308[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4812 = _T_4811 & _GEN_489; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4805 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4807 = _T_4805 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4305; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_4305[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4808 = _T_4807 & _GEN_491; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [59:0] _T_4853 = {_T_4844,_T_4840,_T_4836,_T_4832,_T_4828,_T_4824,_T_4820,_T_4816,_T_4812,_T_4808}; // @[Cat.scala 29:58]
  wire  _T_4801 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4803 = _T_4801 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4302; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_4302[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4804 = _T_4803 & _GEN_493; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4797 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4799 = _T_4797 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4299; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_4299[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4800 = _T_4799 & _GEN_495; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4793 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4795 = _T_4793 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4296; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_4296[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4796 = _T_4795 & _GEN_497; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4789 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4791 = _T_4789 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4293; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_4293[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4792 = _T_4791 & _GEN_499; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4785 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4787 = _T_4785 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4290; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_4290[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4788 = _T_4787 & _GEN_501; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4781 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4783 = _T_4781 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4287; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_4287[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4784 = _T_4783 & _GEN_503; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4777 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4779 = _T_4777 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4284; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_4284[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4780 = _T_4779 & _GEN_505; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4773 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4775 = _T_4773 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4281; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_4281[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4776 = _T_4775 & _GEN_507; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4769 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4771 = _T_4769 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4278; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_4278[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4772 = _T_4771 & _GEN_509; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [113:0] _T_4862 = {_T_4853,_T_4804,_T_4800,_T_4796,_T_4792,_T_4788,_T_4784,_T_4780,_T_4776,_T_4772}; // @[Cat.scala 29:58]
  wire  _T_4765 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4767 = _T_4765 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4275; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_4275[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4768 = _T_4767 & _GEN_511; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4761 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4763 = _T_4761 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4272; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_4272[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4764 = _T_4763 & _GEN_513; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4757 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4759 = _T_4757 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4269; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_4269[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4760 = _T_4759 & _GEN_515; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4753 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4755 = _T_4753 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4266; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_4266[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4756 = _T_4755 & _GEN_517; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4749 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4751 = _T_4749 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4263; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_4263[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4752 = _T_4751 & _GEN_519; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4745 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4747 = _T_4745 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4260; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_4260[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4748 = _T_4747 & _GEN_521; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4741 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4743 = _T_4741 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4257; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_4257[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4744 = _T_4743 & _GEN_523; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4737 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4739 = _T_4737 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4254; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_4254[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4740 = _T_4739 & _GEN_525; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4733 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4735 = _T_4733 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4251; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_4251[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4736 = _T_4735 & _GEN_527; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [167:0] _T_4871 = {_T_4862,_T_4768,_T_4764,_T_4760,_T_4756,_T_4752,_T_4748,_T_4744,_T_4740,_T_4736}; // @[Cat.scala 29:58]
  wire  _T_4729 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4731 = _T_4729 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4248; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_4248[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4732 = _T_4731 & _GEN_529; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4725 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4727 = _T_4725 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4245; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_4245[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4728 = _T_4727 & _GEN_531; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4721 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4723 = _T_4721 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4242; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_4242[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4724 = _T_4723 & _GEN_533; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4717 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4719 = _T_4717 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4239; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_4239[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4720 = _T_4719 & _GEN_535; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4713 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4715 = _T_4713 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4236; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_4236[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4716 = _T_4715 & _GEN_537; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4709 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4711 = _T_4709 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4233; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_4233[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4712 = _T_4711 & _GEN_539; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4705 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4707 = _T_4705 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4230; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_4230[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4708 = _T_4707 & _GEN_541; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4701 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4703 = _T_4701 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4227; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_4227[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4704 = _T_4703 & _GEN_543; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4697 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4699 = _T_4697 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4224; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_4224[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4700 = _T_4699 & _GEN_545; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [221:0] _T_4880 = {_T_4871,_T_4732,_T_4728,_T_4724,_T_4720,_T_4716,_T_4712,_T_4708,_T_4704,_T_4700}; // @[Cat.scala 29:58]
  wire  _T_4693 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4695 = _T_4693 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4221; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_4221[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4696 = _T_4695 & _GEN_547; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4689 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4691 = _T_4689 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4218; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_4218[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4692 = _T_4691 & _GEN_549; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4685 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4687 = _T_4685 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4215; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_4215[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4688 = _T_4687 & _GEN_551; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4681 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4683 = _T_4681 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4212; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_4212[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4684 = _T_4683 & _GEN_553; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4677 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4679 = _T_4677 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4209; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_4209[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4680 = _T_4679 & _GEN_555; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4673 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4675 = _T_4673 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4206; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_4206[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4676 = _T_4675 & _GEN_557; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4669 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4671 = _T_4669 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4203; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_4203[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4672 = _T_4671 & _GEN_559; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4665 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4667 = _T_4665 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4200; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_4200[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4668 = _T_4667 & _GEN_561; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4661 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4663 = _T_4661 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4197; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_4197[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4664 = _T_4663 & _GEN_563; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [275:0] _T_4889 = {_T_4880,_T_4696,_T_4692,_T_4688,_T_4684,_T_4680,_T_4676,_T_4672,_T_4668,_T_4664}; // @[Cat.scala 29:58]
  wire  _T_4657 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4659 = _T_4657 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4194; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_4194[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4660 = _T_4659 & _GEN_565; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4653 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4655 = _T_4653 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4191; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_4191[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4656 = _T_4655 & _GEN_567; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4649 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4651 = _T_4649 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4188; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_4188[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4652 = _T_4651 & _GEN_569; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4645 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4647 = _T_4645 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4185; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_4185[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4648 = _T_4647 & _GEN_571; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4641 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4643 = _T_4641 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4182; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_4182[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4644 = _T_4643 & _GEN_573; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4637 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4639 = _T_4637 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4179; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_4179[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4640 = _T_4639 & _GEN_575; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4633 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4635 = _T_4633 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4176; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_4176[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4636 = _T_4635 & _GEN_577; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4629 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4631 = _T_4629 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4173; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_4173[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4632 = _T_4631 & _GEN_579; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4625 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4627 = _T_4625 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4170; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_4170[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4628 = _T_4627 & _GEN_581; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [329:0] _T_4898 = {_T_4889,_T_4660,_T_4656,_T_4652,_T_4648,_T_4644,_T_4640,_T_4636,_T_4632,_T_4628}; // @[Cat.scala 29:58]
  wire  _T_4621 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4623 = _T_4621 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4167; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_4167[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4624 = _T_4623 & _GEN_583; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4617 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4619 = _T_4617 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4164; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_4164[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4620 = _T_4619 & _GEN_585; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4613 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4615 = _T_4613 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4161; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_4161[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4616 = _T_4615 & _GEN_587; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4609 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4611 = _T_4609 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4158; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_4158[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4612 = _T_4611 & _GEN_589; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4605 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4607 = _T_4605 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4155; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_4155[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4608 = _T_4607 & _GEN_591; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4601 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4603 = _T_4601 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4152; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_4152[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4604 = _T_4603 & _GEN_593; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4597 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4599 = _T_4597 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4149; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_4149[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4600 = _T_4599 & _GEN_595; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4593 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4595 = _T_4593 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4146; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_4146[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4596 = _T_4595 & _GEN_597; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4589 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4591 = _T_4589 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4143; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_4143[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4592 = _T_4591 & _GEN_599; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [383:0] _T_4907 = {_T_4898,_T_4624,_T_4620,_T_4616,_T_4612,_T_4608,_T_4604,_T_4600,_T_4596,_T_4592}; // @[Cat.scala 29:58]
  wire  _T_4585 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4587 = _T_4585 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4140; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_4140[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4588 = _T_4587 & _GEN_600; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4581 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4583 = _T_4581 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4137; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_4137[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4584 = _T_4583 & _GEN_601; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4577 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4579 = _T_4577 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4134; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_4134[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4580 = _T_4579 & _GEN_602; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4573 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4575 = _T_4573 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4131; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_4131[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4576 = _T_4575 & _GEN_603; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4569 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4571 = _T_4569 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4128; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_4128[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4572 = _T_4571 & _GEN_604; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4565 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4567 = _T_4565 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4125; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_4125[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4568 = _T_4567 & _GEN_605; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4561 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4563 = _T_4561 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4122; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_4122[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4564 = _T_4563 & _GEN_606; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4557 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4559 = _T_4557 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4119; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_4119[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4560 = _T_4559 & _GEN_607; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4553 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4555 = _T_4553 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4116; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_4116[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4556 = _T_4555 & _GEN_608; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [437:0] _T_4916 = {_T_4907,_T_4588,_T_4584,_T_4580,_T_4576,_T_4572,_T_4568,_T_4564,_T_4560,_T_4556}; // @[Cat.scala 29:58]
  wire  _T_4549 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4551 = _T_4549 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4113; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_4113[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4552 = _T_4551 & _GEN_609; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4545 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4547 = _T_4545 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4110; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_4110[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4548 = _T_4547 & _GEN_610; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4541 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4543 = _T_4541 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4107; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_4107[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4544 = _T_4543 & _GEN_611; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4537 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4539 = _T_4537 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4104; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_4104[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4540 = _T_4539 & _GEN_612; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4533 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4535 = _T_4533 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4101; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_4101[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4536 = _T_4535 & _GEN_613; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4529 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4531 = _T_4529 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4098; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_4098[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4532 = _T_4531 & _GEN_614; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4525 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4527 = _T_4525 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4095; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_4095[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4528 = _T_4527 & _GEN_615; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4521 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4523 = _T_4521 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4092; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_4092[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4524 = _T_4523 & _GEN_616; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4517 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4519 = _T_4517 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4089; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_4089[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4520 = _T_4519 & _GEN_617; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [491:0] _T_4925 = {_T_4916,_T_4552,_T_4548,_T_4544,_T_4540,_T_4536,_T_4532,_T_4528,_T_4524,_T_4520}; // @[Cat.scala 29:58]
  wire  _T_4513 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4515 = _T_4513 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4086; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_4086[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4516 = _T_4515 & _GEN_618; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4509 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4511 = _T_4509 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4083; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_4083[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4512 = _T_4511 & _GEN_619; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4505 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4507 = _T_4505 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4080; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_4080[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4508 = _T_4507 & _GEN_620; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4501 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4503 = _T_4501 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4077; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_4077[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4504 = _T_4503 & _GEN_621; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4497 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4499 = _T_4497 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4074; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_4074[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4500 = _T_4499 & _GEN_622; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4493 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4495 = _T_4493 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4071; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_4071[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4496 = _T_4495 & _GEN_623; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4489 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4491 = _T_4489 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4068; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_4068[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4492 = _T_4491 & _GEN_624; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4485 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4487 = _T_4485 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4065; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_4065[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4488 = _T_4487 & _GEN_625; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4481 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4483 = _T_4481 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4062; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_4062[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4484 = _T_4483 & _GEN_626; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [545:0] _T_4934 = {_T_4925,_T_4516,_T_4512,_T_4508,_T_4504,_T_4500,_T_4496,_T_4492,_T_4488,_T_4484}; // @[Cat.scala 29:58]
  wire  _T_4477 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4479 = _T_4477 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4059; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_4059[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4480 = _T_4479 & _GEN_627; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4473 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4475 = _T_4473 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4056; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_4056[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4476 = _T_4475 & _GEN_628; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4469 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4471 = _T_4469 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4053; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_4053[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4472 = _T_4471 & _GEN_629; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4465 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4467 = _T_4465 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4050; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_4050[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4468 = _T_4467 & _GEN_630; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4461 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4463 = _T_4461 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4047; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_4047[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4464 = _T_4463 & _GEN_631; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4457 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4459 = _T_4457 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4044; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_4044[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4460 = _T_4459 & _GEN_632; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4453 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4455 = _T_4453 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4041; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_4041[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4456 = _T_4455 & _GEN_633; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4449 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4451 = _T_4449 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4038; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_4038[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4452 = _T_4451 & _GEN_634; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4445 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4447 = _T_4445 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4035; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_4035[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4448 = _T_4447 & _GEN_635; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [599:0] _T_4943 = {_T_4934,_T_4480,_T_4476,_T_4472,_T_4468,_T_4464,_T_4460,_T_4456,_T_4452,_T_4448}; // @[Cat.scala 29:58]
  wire  _T_4441 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4443 = _T_4441 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4032; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_4032[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4444 = _T_4443 & _GEN_636; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4437 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4439 = _T_4437 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4029; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_4029[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4440 = _T_4439 & _GEN_637; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4433 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4435 = _T_4433 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4026; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_4026[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4436 = _T_4435 & _GEN_638; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4429 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4431 = _T_4429 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4023; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_4023[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4432 = _T_4431 & _GEN_639; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4425 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4427 = _T_4425 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4020; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_4020[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4428 = _T_4427 & _GEN_640; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4421 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4423 = _T_4421 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4017; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_4017[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4424 = _T_4423 & _GEN_641; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4417 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4419 = _T_4417 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4014; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_4014[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4420 = _T_4419 & _GEN_642; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4413 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4415 = _T_4413 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4011; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_4011[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4416 = _T_4415 & _GEN_643; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4409 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4411 = _T_4409 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4008; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_4008[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4412 = _T_4411 & _GEN_644; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [653:0] _T_4952 = {_T_4943,_T_4444,_T_4440,_T_4436,_T_4432,_T_4428,_T_4424,_T_4420,_T_4416,_T_4412}; // @[Cat.scala 29:58]
  wire  _T_4405 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4407 = _T_4405 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4005; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_4005[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4408 = _T_4407 & _GEN_645; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4401 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4403 = _T_4401 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4002; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_4002[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4404 = _T_4403 & _GEN_646; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4397 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4399 = _T_4397 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3999; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_3999[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4400 = _T_4399 & _GEN_647; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4393 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4395 = _T_4393 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3996; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_3996[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4396 = _T_4395 & _GEN_648; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4389 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4391 = _T_4389 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3993; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_3993[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4392 = _T_4391 & _GEN_649; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4385 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4387 = _T_4385 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3990; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_3990[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4388 = _T_4387 & _GEN_650; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4381 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4383 = _T_4381 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3987; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_3987[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4384 = _T_4383 & _GEN_651; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4377 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4379 = _T_4377 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3984; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_3984[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4380 = _T_4379 & _GEN_652; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4373 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4375 = _T_4373 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3981; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_3981[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4376 = _T_4375 & _GEN_653; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [707:0] _T_4961 = {_T_4952,_T_4408,_T_4404,_T_4400,_T_4396,_T_4392,_T_4388,_T_4384,_T_4380,_T_4376}; // @[Cat.scala 29:58]
  wire  _T_4369 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4371 = _T_4369 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3978; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3978[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4372 = _T_4371 & _GEN_654; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4365 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4367 = _T_4365 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3975; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3975[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4368 = _T_4367 & _GEN_655; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4361 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4363 = _T_4361 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3972; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3972[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4364 = _T_4363 & _GEN_656; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4357 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4359 = _T_4357 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3969; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3969[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4360 = _T_4359 & _GEN_657; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4353 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4355 = _T_4353 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3966; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3966[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4356 = _T_4355 & _GEN_658; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4349 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4351 = _T_4349 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3963; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3963[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4352 = _T_4351 & _GEN_659; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4345 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4347 = _T_4345 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3960; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3960[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4348 = _T_4347 & _GEN_660; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4341 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4343 = _T_4341 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3957; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3957[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4344 = _T_4343 & _GEN_661; // @[el2_ifu_mem_ctl.scala 766:130]
  wire  _T_4337 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4339 = _T_4337 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3954; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3954[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4340 = _T_4339 & _GEN_662; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [761:0] _T_4970 = {_T_4961,_T_4372,_T_4368,_T_4364,_T_4360,_T_4356,_T_4352,_T_4348,_T_4344,_T_4340}; // @[Cat.scala 29:58]
  wire  _T_4333 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 766:121]
  wire [5:0] _T_4335 = _T_4333 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3951; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3951[0]; // @[el2_ifu_mem_ctl.scala 761:30 el2_ifu_mem_ctl.scala 763:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [5:0] _T_4336 = _T_4335 & _GEN_663; // @[el2_ifu_mem_ctl.scala 766:130]
  wire [767:0] _T_4971 = {_T_4970,_T_4336}; // @[Cat.scala 29:58]
  wire  way_status = _T_4971[0]; // @[el2_ifu_mem_ctl.scala 766:16]
  wire  _T_187 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 309:96]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 313:25]
  wire [2:0] _T_198 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_198; // @[el2_ifu_mem_ctl.scala 318:45]
  wire  _T_204 = _T_223 | _T_231; // @[el2_ifu_mem_ctl.scala 323:59]
  wire  _T_206 = _T_204 | _T_2217; // @[el2_ifu_mem_ctl.scala 323:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_206; // @[el2_ifu_mem_ctl.scala 323:41]
  wire  _T_211 = _T_219 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 329:39]
  wire  _T_213 = _T_211 & _T_187; // @[el2_ifu_mem_ctl.scala 329:60]
  wire  _T_217 = _T_213 & _T_204; // @[el2_ifu_mem_ctl.scala 329:78]
  wire  ic_act_hit_f = _T_217 & _T_239; // @[el2_ifu_mem_ctl.scala 329:126]
  wire  _T_254 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 336:31]
  wire  _T_255 = _T_254 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 336:46]
  wire  _T_256 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 336:94]
  wire  uncacheable_miss_in = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 337:84]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2600 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 662:48]
  wire  _T_2601 = _T_2600 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 662:52]
  wire  bus_ifu_wr_data_error_ff = _T_2601 & miss_pending; // @[el2_ifu_mem_ctl.scala 662:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 412:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 411:55]
  wire  _T_268 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 340:145]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 589:52]
  wire  _T_289 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 352:36]
  wire  _T_290 = miss_pending & _T_289; // @[el2_ifu_mem_ctl.scala 352:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 353:25]
  wire  _T_291 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 352:72]
  wire  reset_ic_in = _T_290 & _T_291; // @[el2_ifu_mem_ctl.scala 352:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 354:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 362:23]
  wire  _T_305 = _T_2231 & flush_final_f; // @[el2_ifu_mem_ctl.scala 366:87]
  wire  _T_306 = ~_T_305; // @[el2_ifu_mem_ctl.scala 366:55]
  wire  _T_307 = io_ifc_fetch_req_bf & _T_306; // @[el2_ifu_mem_ctl.scala 366:53]
  wire  stream_miss_f = stream_hit_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 502:83]
  wire  _T_308 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 366:106]
  wire  ifc_fetch_req_qual_bf = _T_307 & _T_308; // @[el2_ifu_mem_ctl.scala 366:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 372:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_2237 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 507:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2237}; // @[Cat.scala 29:58]
  wire  _T_2238 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2262 = _T_2238 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2241 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2263 = _T_2241 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2270 = _T_2262 | _T_2263; // @[Mux.scala 27:72]
  wire  _T_2244 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2264 = _T_2244 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2271 = _T_2270 | _T_2264; // @[Mux.scala 27:72]
  wire  _T_2247 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2265 = _T_2247 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2272 = _T_2271 | _T_2265; // @[Mux.scala 27:72]
  wire  _T_2250 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2266 = _T_2250 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2273 = _T_2272 | _T_2266; // @[Mux.scala 27:72]
  wire  _T_2253 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2267 = _T_2253 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2274 = _T_2273 | _T_2267; // @[Mux.scala 27:72]
  wire  _T_2256 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2268 = _T_2256 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2275 = _T_2274 | _T_2268; // @[Mux.scala 27:72]
  wire  _T_2259 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2269 = _T_2259 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2275 | _T_2269; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 509:46]
  wire  _T_320 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 378:35]
  wire  _T_322 = _T_320 & _T_52; // @[el2_ifu_mem_ctl.scala 378:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 659:61]
  wire  _T_2594 = ic_act_miss_f_delayed & _T_2232; // @[el2_ifu_mem_ctl.scala 660:53]
  wire  reset_tag_valid_for_miss = _T_2594 & _T_52; // @[el2_ifu_mem_ctl.scala 660:84]
  wire  sel_mb_addr = _T_322 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 378:79]
  wire [30:0] _T_327 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_329 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 380:37]
  wire [30:0] _T_330 = sel_mb_addr ? _T_327 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_331 = _T_329 ? ifu_fetch_addr_int_f : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ic_rw_addr = _T_330 | _T_331; // @[Mux.scala 27:72]
  wire  _T_336 = _T_322 & last_beat; // @[el2_ifu_mem_ctl.scala 382:84]
  wire  _T_2588 = ~_T_2600; // @[el2_ifu_mem_ctl.scala 657:84]
  wire  _T_2589 = _T_92 & _T_2588; // @[el2_ifu_mem_ctl.scala 657:82]
  wire  bus_ifu_wr_en_ff_q = _T_2589 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 657:108]
  wire  sel_mb_status_addr = _T_336 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 382:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_327 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 383:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [7:0] _T_560 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_569 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_560}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_577 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_586 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_577}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_587 = {_T_586,_T_569}; // @[el2_lib.scala 348:27]
  wire  _T_588 = ^_T_587; // @[el2_lib.scala 348:34]
  wire [7:0] _T_595 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_604 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_595}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_612 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_621 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_612}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_622 = {_T_621,_T_604}; // @[el2_lib.scala 348:44]
  wire  _T_623 = ^_T_622; // @[el2_lib.scala 348:51]
  wire [7:0] _T_630 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_639 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_630}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_647 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_656 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_647}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_657 = {_T_656,_T_639}; // @[el2_lib.scala 348:61]
  wire  _T_658 = ^_T_657; // @[el2_lib.scala 348:68]
  wire [6:0] _T_664 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_672 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_664}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_679 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_688 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_679,_T_672}; // @[el2_lib.scala 348:78]
  wire  _T_689 = ^_T_688; // @[el2_lib.scala 348:85]
  wire [6:0] _T_695 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_703 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_695}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_710 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_719 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_710,_T_703}; // @[el2_lib.scala 348:95]
  wire  _T_720 = ^_T_719; // @[el2_lib.scala 348:102]
  wire [6:0] _T_726 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_734 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_726}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_750 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_710,_T_734}; // @[el2_lib.scala 348:112]
  wire  _T_751 = ^_T_750; // @[el2_lib.scala 348:119]
  wire [6:0] _T_757 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 348:129]
  wire  _T_758 = ^_T_757; // @[el2_lib.scala 348:136]
  wire [3:0] _T_2278 = {ifu_bus_rid_ff[2:1],_T_2237,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2279 = _T_2278 == 4'h0; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1285; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_0 = _T_1285[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2326 = _T_2279 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2282 = _T_2278 == 4'h1; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1287; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_1 = _T_1287[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2327 = _T_2282 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2342 = _T_2326 | _T_2327; // @[Mux.scala 27:72]
  wire  _T_2285 = _T_2278 == 4'h2; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1289; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_2 = _T_1289[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2328 = _T_2285 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2343 = _T_2342 | _T_2328; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2278 == 4'h3; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1291; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_3 = _T_1291[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2329 = _T_2288 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2344 = _T_2343 | _T_2329; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2278 == 4'h4; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1293; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_4 = _T_1293[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2330 = _T_2291 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2345 = _T_2344 | _T_2330; // @[Mux.scala 27:72]
  wire  _T_2294 = _T_2278 == 4'h5; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1295; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_5 = _T_1295[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2331 = _T_2294 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2346 = _T_2345 | _T_2331; // @[Mux.scala 27:72]
  wire  _T_2297 = _T_2278 == 4'h6; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1297; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_6 = _T_1297[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2332 = _T_2297 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2347 = _T_2346 | _T_2332; // @[Mux.scala 27:72]
  wire  _T_2300 = _T_2278 == 4'h7; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1299; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_7 = _T_1299[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2333 = _T_2300 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2348 = _T_2347 | _T_2333; // @[Mux.scala 27:72]
  wire  _T_2303 = _T_2278 == 4'h8; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1301; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_8 = _T_1301[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2334 = _T_2303 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2349 = _T_2348 | _T_2334; // @[Mux.scala 27:72]
  wire  _T_2306 = _T_2278 == 4'h9; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1303; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_9 = _T_1303[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2335 = _T_2306 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2350 = _T_2349 | _T_2335; // @[Mux.scala 27:72]
  wire  _T_2309 = _T_2278 == 4'ha; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1305; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_10 = _T_1305[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2336 = _T_2309 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2351 = _T_2350 | _T_2336; // @[Mux.scala 27:72]
  wire  _T_2312 = _T_2278 == 4'hb; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1307; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_11 = _T_1307[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2337 = _T_2312 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2352 = _T_2351 | _T_2337; // @[Mux.scala 27:72]
  wire  _T_2315 = _T_2278 == 4'hc; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1309; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_12 = _T_1309[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2338 = _T_2315 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2353 = _T_2352 | _T_2338; // @[Mux.scala 27:72]
  wire  _T_2318 = _T_2278 == 4'hd; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1311; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_13 = _T_1311[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2339 = _T_2318 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2354 = _T_2353 | _T_2339; // @[Mux.scala 27:72]
  wire  _T_2321 = _T_2278 == 4'he; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1313; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_14 = _T_1313[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 445:26]
  wire [31:0] _T_2340 = _T_2321 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2355 = _T_2354 | _T_2340; // @[Mux.scala 27:72]
  wire  _T_2324 = _T_2278 == 4'hf; // @[el2_ifu_mem_ctl.scala 510:89]
  reg [63:0] _T_1315; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_15 = _T_1315[31:0]; // @[el2_ifu_mem_ctl.scala 443:31 el2_ifu_mem_ctl.scala 446:28]
  wire [31:0] _T_2341 = _T_2324 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2356 = _T_2355 | _T_2341; // @[Mux.scala 27:72]
  wire [3:0] _T_2358 = {ifu_bus_rid_ff[2:1],_T_2237,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2359 = _T_2358 == 4'h0; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2382 = _T_2359 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2362 = _T_2358 == 4'h1; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2383 = _T_2362 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2390 = _T_2382 | _T_2383; // @[Mux.scala 27:72]
  wire  _T_2365 = _T_2358 == 4'h2; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2384 = _T_2365 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2391 = _T_2390 | _T_2384; // @[Mux.scala 27:72]
  wire  _T_2368 = _T_2358 == 4'h3; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2385 = _T_2368 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2392 = _T_2391 | _T_2385; // @[Mux.scala 27:72]
  wire  _T_2371 = _T_2358 == 4'h4; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2386 = _T_2371 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2393 = _T_2392 | _T_2386; // @[Mux.scala 27:72]
  wire  _T_2374 = _T_2358 == 4'h5; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2387 = _T_2374 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2394 = _T_2393 | _T_2387; // @[Mux.scala 27:72]
  wire  _T_2377 = _T_2358 == 4'h6; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2388 = _T_2377 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2395 = _T_2394 | _T_2388; // @[Mux.scala 27:72]
  wire  _T_2380 = _T_2358 == 4'h7; // @[el2_ifu_mem_ctl.scala 511:64]
  wire [31:0] _T_2389 = _T_2380 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2396 = _T_2395 | _T_2389; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2356,_T_2396}; // @[Cat.scala 29:58]
  wire [7:0] _T_982 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_991 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_982}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_999 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_1008 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_999}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_1009 = {_T_1008,_T_991}; // @[el2_lib.scala 348:27]
  wire  _T_1010 = ^_T_1009; // @[el2_lib.scala 348:34]
  wire [7:0] _T_1017 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_1026 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1017}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_1034 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_1043 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1034}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_1044 = {_T_1043,_T_1026}; // @[el2_lib.scala 348:44]
  wire  _T_1045 = ^_T_1044; // @[el2_lib.scala 348:51]
  wire [7:0] _T_1052 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_1061 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1052}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_1069 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_1078 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1069}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_1079 = {_T_1078,_T_1061}; // @[el2_lib.scala 348:61]
  wire  _T_1080 = ^_T_1079; // @[el2_lib.scala 348:68]
  wire [6:0] _T_1086 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_1094 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1086}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_1101 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_1110 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1101,_T_1094}; // @[el2_lib.scala 348:78]
  wire  _T_1111 = ^_T_1110; // @[el2_lib.scala 348:85]
  wire [6:0] _T_1117 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_1125 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1117}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_1132 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_1141 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1132,_T_1125}; // @[el2_lib.scala 348:95]
  wire  _T_1142 = ^_T_1141; // @[el2_lib.scala 348:102]
  wire [6:0] _T_1148 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_1156 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_1148}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_1172 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1132,_T_1156}; // @[el2_lib.scala 348:112]
  wire  _T_1173 = ^_T_1172; // @[el2_lib.scala 348:119]
  wire [6:0] _T_1179 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 348:129]
  wire  _T_1180 = ^_T_1179; // @[el2_lib.scala 348:136]
  wire [70:0] _T_1227 = {_T_588,_T_623,_T_658,_T_689,_T_720,_T_751,_T_758,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1226 = {_T_1010,_T_1045,_T_1080,_T_1111,_T_1142,_T_1173,_T_1180,_T_2356,_T_2396}; // @[Cat.scala 29:58]
  wire [141:0] _T_1228 = {_T_588,_T_623,_T_658,_T_689,_T_720,_T_751,_T_758,ifu_bus_rdata_ff,_T_1226}; // @[Cat.scala 29:58]
  wire [141:0] _T_1231 = {_T_1010,_T_1045,_T_1080,_T_1111,_T_1142,_T_1173,_T_1180,_T_2356,_T_2396,_T_1227}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1228 : _T_1231; // @[el2_ifu_mem_ctl.scala 404:28]
  wire  _T_1188 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 394:56]
  wire  _T_1189 = _T_1188 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 394:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 457:28]
  wire  _T_1391 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  bus_ifu_wr_en = _T_14 & miss_pending; // @[el2_ifu_mem_ctl.scala 655:35]
  wire  _T_1276 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1276; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1317 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 448:118]
  wire  _T_1318 = ic_miss_buff_data_valid[0] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1318; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1414 = _T_1391 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1394 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  _T_1277 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1277; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1321 = ic_miss_buff_data_valid[1] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1321; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1415 = _T_1394 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1422 = _T_1414 | _T_1415; // @[Mux.scala 27:72]
  wire  _T_1397 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  _T_1278 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1278; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1324 = ic_miss_buff_data_valid[2] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1324; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1416 = _T_1397 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1423 = _T_1422 | _T_1416; // @[Mux.scala 27:72]
  wire  _T_1400 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  _T_1279 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1279; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1327 = ic_miss_buff_data_valid[3] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1327; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1417 = _T_1400 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1424 = _T_1423 | _T_1417; // @[Mux.scala 27:72]
  wire  _T_1403 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  _T_1280 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1280; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1330 = ic_miss_buff_data_valid[4] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1330; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1418 = _T_1403 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1425 = _T_1424 | _T_1418; // @[Mux.scala 27:72]
  wire  _T_1406 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  _T_1281 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1281; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1333 = ic_miss_buff_data_valid[5] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1333; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1419 = _T_1406 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1426 = _T_1425 | _T_1419; // @[Mux.scala 27:72]
  wire  _T_1409 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  _T_1282 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1336 = ic_miss_buff_data_valid[6] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1336; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1420 = _T_1409 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1427 = _T_1426 | _T_1420; // @[Mux.scala 27:72]
  wire  _T_1412 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 459:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 442:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 442:73]
  wire  _T_1339 = ic_miss_buff_data_valid[7] & _T_1317; // @[el2_ifu_mem_ctl.scala 448:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1339; // @[el2_ifu_mem_ctl.scala 448:88]
  wire  _T_1421 = _T_1412 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1427 | _T_1421; // @[Mux.scala 27:72]
  wire  _T_1430 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 460:58]
  wire  _T_1431 = bypass_valid_value_check & _T_1430; // @[el2_ifu_mem_ctl.scala 460:56]
  wire  _T_1433 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 460:77]
  wire  _T_1434 = _T_1431 & _T_1433; // @[el2_ifu_mem_ctl.scala 460:75]
  wire  _T_1439 = _T_1431 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 461:75]
  wire  _T_1440 = _T_1434 | _T_1439; // @[el2_ifu_mem_ctl.scala 460:95]
  wire  _T_1442 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 462:56]
  wire  _T_1445 = _T_1442 & _T_1433; // @[el2_ifu_mem_ctl.scala 462:74]
  wire  _T_1446 = _T_1440 | _T_1445; // @[el2_ifu_mem_ctl.scala 461:94]
  wire  _T_1450 = _T_1442 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 463:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 458:70]
  wire  _T_1451 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1467 = _T_1451 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1453 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1468 = _T_1453 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1475 = _T_1467 | _T_1468; // @[Mux.scala 27:72]
  wire  _T_1455 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1469 = _T_1455 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1476 = _T_1475 | _T_1469; // @[Mux.scala 27:72]
  wire  _T_1457 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1470 = _T_1457 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1477 = _T_1476 | _T_1470; // @[Mux.scala 27:72]
  wire  _T_1459 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1471 = _T_1459 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1478 = _T_1477 | _T_1471; // @[Mux.scala 27:72]
  wire  _T_1461 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1472 = _T_1461 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1479 = _T_1478 | _T_1472; // @[Mux.scala 27:72]
  wire  _T_1463 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1473 = _T_1463 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1480 = _T_1479 | _T_1473; // @[Mux.scala 27:72]
  wire  _T_1465 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 463:132]
  wire  _T_1474 = _T_1465 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1481 = _T_1480 | _T_1474; // @[Mux.scala 27:72]
  wire  _T_1483 = _T_1450 & _T_1481; // @[el2_ifu_mem_ctl.scala 463:69]
  wire  _T_1484 = _T_1446 | _T_1483; // @[el2_ifu_mem_ctl.scala 462:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 464:95]
  wire  _T_1487 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 464:95]
  wire  _T_1488 = bypass_valid_value_check & _T_1487; // @[el2_ifu_mem_ctl.scala 464:56]
  wire  bypass_data_ready_in = _T_1484 | _T_1488; // @[el2_ifu_mem_ctl.scala 463:181]
  wire  _T_1489 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 468:53]
  wire  _T_1490 = _T_1489 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 468:73]
  wire  _T_1492 = _T_1490 & _T_309; // @[el2_ifu_mem_ctl.scala 468:96]
  wire  _T_1494 = _T_1492 & _T_61; // @[el2_ifu_mem_ctl.scala 468:118]
  wire  _T_1496 = crit_wd_byp_ok_ff & _T_52; // @[el2_ifu_mem_ctl.scala 469:73]
  wire  _T_1498 = _T_1496 & _T_309; // @[el2_ifu_mem_ctl.scala 469:96]
  wire  _T_1500 = _T_1498 & _T_61; // @[el2_ifu_mem_ctl.scala 469:118]
  wire  _T_1501 = _T_1494 | _T_1500; // @[el2_ifu_mem_ctl.scala 468:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 471:58]
  wire  _T_1502 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 470:54]
  wire  _T_1503 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 470:76]
  wire  _T_1504 = _T_1502 & _T_1503; // @[el2_ifu_mem_ctl.scala 470:74]
  wire  _T_1506 = _T_1504 & _T_309; // @[el2_ifu_mem_ctl.scala 470:96]
  wire  ic_crit_wd_rdy_new_in = _T_1501 | _T_1506; // @[el2_ifu_mem_ctl.scala 469:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 665:43]
  wire  _T_1243 = ic_crit_wd_rdy | _T_2217; // @[el2_ifu_mem_ctl.scala 416:38]
  wire  _T_1245 = _T_1243 | _T_2232; // @[el2_ifu_mem_ctl.scala 416:64]
  wire  _T_1246 = ~_T_1245; // @[el2_ifu_mem_ctl.scala 416:21]
  wire  _T_1247 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 416:98]
  wire  sel_ic_data = _T_1246 & _T_1247; // @[el2_ifu_mem_ctl.scala 416:96]
  wire  _T_2399 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 513:44]
  wire  _T_1600 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 482:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 454:60]
  wire  _T_1544 = _T_1391 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1545 = _T_1394 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1552 = _T_1544 | _T_1545; // @[Mux.scala 27:72]
  wire  _T_1546 = _T_1397 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1552 | _T_1546; // @[Mux.scala 27:72]
  wire  _T_1547 = _T_1400 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1554 = _T_1553 | _T_1547; // @[Mux.scala 27:72]
  wire  _T_1548 = _T_1403 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1554 | _T_1548; // @[Mux.scala 27:72]
  wire  _T_1549 = _T_1406 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1555 | _T_1549; // @[Mux.scala 27:72]
  wire  _T_1550 = _T_1409 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1556 | _T_1550; // @[Mux.scala 27:72]
  wire  _T_1551 = _T_1412 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1557 | _T_1551; // @[Mux.scala 27:72]
  wire  _T_1583 = _T_2144 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1584 = _T_2147 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1591 = _T_1583 | _T_1584; // @[Mux.scala 27:72]
  wire  _T_1585 = _T_2150 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1592 = _T_1591 | _T_1585; // @[Mux.scala 27:72]
  wire  _T_1586 = _T_2153 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1593 = _T_1592 | _T_1586; // @[Mux.scala 27:72]
  wire  _T_1587 = _T_2156 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1594 = _T_1593 | _T_1587; // @[Mux.scala 27:72]
  wire  _T_1588 = _T_2159 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1595 = _T_1594 | _T_1588; // @[Mux.scala 27:72]
  wire  _T_1589 = _T_2162 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1596 = _T_1595 | _T_1589; // @[Mux.scala 27:72]
  wire  _T_1590 = _T_2165 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1596 | _T_1590; // @[Mux.scala 27:72]
  wire  _T_1601 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 484:70]
  wire  ifu_byp_data_err_new = _T_1600 ? ic_miss_buff_data_error_bypass : _T_1601; // @[el2_ifu_mem_ctl.scala 482:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 426:42]
  wire  _T_2400 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 513:91]
  wire  _T_2401 = ~_T_2400; // @[el2_ifu_mem_ctl.scala 513:60]
  wire  ic_rd_parity_final_err = _T_2399 & _T_2401; // @[el2_ifu_mem_ctl.scala 513:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9035 = _T_4333 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 796:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9037 = _T_4337 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9290 = _T_9035 | _T_9037; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9039 = _T_4341 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9291 = _T_9290 | _T_9039; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9041 = _T_4345 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9292 = _T_9291 | _T_9041; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9043 = _T_4349 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9293 = _T_9292 | _T_9043; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9045 = _T_4353 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9294 = _T_9293 | _T_9045; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9047 = _T_4357 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9295 = _T_9294 | _T_9047; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9049 = _T_4361 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9296 = _T_9295 | _T_9049; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9051 = _T_4365 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9297 = _T_9296 | _T_9051; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9053 = _T_4369 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9298 = _T_9297 | _T_9053; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9055 = _T_4373 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9299 = _T_9298 | _T_9055; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9057 = _T_4377 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9300 = _T_9299 | _T_9057; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9059 = _T_4381 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9301 = _T_9300 | _T_9059; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9061 = _T_4385 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9302 = _T_9301 | _T_9061; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9063 = _T_4389 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9303 = _T_9302 | _T_9063; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9065 = _T_4393 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9304 = _T_9303 | _T_9065; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9067 = _T_4397 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9305 = _T_9304 | _T_9067; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9069 = _T_4401 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9306 = _T_9305 | _T_9069; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9071 = _T_4405 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9307 = _T_9306 | _T_9071; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9073 = _T_4409 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9308 = _T_9307 | _T_9073; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9075 = _T_4413 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9309 = _T_9308 | _T_9075; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9077 = _T_4417 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9310 = _T_9309 | _T_9077; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9079 = _T_4421 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9311 = _T_9310 | _T_9079; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9081 = _T_4425 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9312 = _T_9311 | _T_9081; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9083 = _T_4429 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9313 = _T_9312 | _T_9083; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9085 = _T_4433 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9314 = _T_9313 | _T_9085; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9087 = _T_4437 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9315 = _T_9314 | _T_9087; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9089 = _T_4441 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9316 = _T_9315 | _T_9089; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9091 = _T_4445 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9317 = _T_9316 | _T_9091; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9093 = _T_4449 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9318 = _T_9317 | _T_9093; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9095 = _T_4453 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9319 = _T_9318 | _T_9095; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9097 = _T_4457 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9320 = _T_9319 | _T_9097; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9099 = _T_4461 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9321 = _T_9320 | _T_9099; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9101 = _T_4465 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9322 = _T_9321 | _T_9101; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9103 = _T_4469 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9323 = _T_9322 | _T_9103; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9105 = _T_4473 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9324 = _T_9323 | _T_9105; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9107 = _T_4477 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9325 = _T_9324 | _T_9107; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9109 = _T_4481 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9326 = _T_9325 | _T_9109; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9111 = _T_4485 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9327 = _T_9326 | _T_9111; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9113 = _T_4489 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9328 = _T_9327 | _T_9113; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9115 = _T_4493 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9329 = _T_9328 | _T_9115; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9117 = _T_4497 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9330 = _T_9329 | _T_9117; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9119 = _T_4501 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9331 = _T_9330 | _T_9119; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9121 = _T_4505 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9332 = _T_9331 | _T_9121; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9123 = _T_4509 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9333 = _T_9332 | _T_9123; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9125 = _T_4513 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9334 = _T_9333 | _T_9125; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9127 = _T_4517 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9335 = _T_9334 | _T_9127; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9129 = _T_4521 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9336 = _T_9335 | _T_9129; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9131 = _T_4525 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9337 = _T_9336 | _T_9131; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9133 = _T_4529 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9338 = _T_9337 | _T_9133; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9135 = _T_4533 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9339 = _T_9338 | _T_9135; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9137 = _T_4537 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9340 = _T_9339 | _T_9137; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9139 = _T_4541 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9341 = _T_9340 | _T_9139; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9141 = _T_4545 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9342 = _T_9341 | _T_9141; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9143 = _T_4549 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9343 = _T_9342 | _T_9143; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9145 = _T_4553 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9344 = _T_9343 | _T_9145; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9147 = _T_4557 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9345 = _T_9344 | _T_9147; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9149 = _T_4561 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9346 = _T_9345 | _T_9149; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9151 = _T_4565 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9347 = _T_9346 | _T_9151; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9153 = _T_4569 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9348 = _T_9347 | _T_9153; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9155 = _T_4573 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9349 = _T_9348 | _T_9155; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9157 = _T_4577 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9350 = _T_9349 | _T_9157; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9159 = _T_4581 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9351 = _T_9350 | _T_9159; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9161 = _T_4585 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9352 = _T_9351 | _T_9161; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9163 = _T_4589 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9353 = _T_9352 | _T_9163; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9165 = _T_4593 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9354 = _T_9353 | _T_9165; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9167 = _T_4597 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9355 = _T_9354 | _T_9167; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9169 = _T_4601 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9356 = _T_9355 | _T_9169; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9171 = _T_4605 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9357 = _T_9356 | _T_9171; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9173 = _T_4609 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9358 = _T_9357 | _T_9173; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9175 = _T_4613 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9359 = _T_9358 | _T_9175; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9177 = _T_4617 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9360 = _T_9359 | _T_9177; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9179 = _T_4621 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9361 = _T_9360 | _T_9179; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9181 = _T_4625 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9362 = _T_9361 | _T_9181; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9183 = _T_4629 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9363 = _T_9362 | _T_9183; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9185 = _T_4633 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9364 = _T_9363 | _T_9185; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9187 = _T_4637 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9365 = _T_9364 | _T_9187; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9189 = _T_4641 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9366 = _T_9365 | _T_9189; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9191 = _T_4645 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9367 = _T_9366 | _T_9191; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9193 = _T_4649 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9368 = _T_9367 | _T_9193; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9195 = _T_4653 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9369 = _T_9368 | _T_9195; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9197 = _T_4657 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9370 = _T_9369 | _T_9197; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9199 = _T_4661 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9371 = _T_9370 | _T_9199; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9201 = _T_4665 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9372 = _T_9371 | _T_9201; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9203 = _T_4669 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9373 = _T_9372 | _T_9203; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9205 = _T_4673 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9374 = _T_9373 | _T_9205; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9207 = _T_4677 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9375 = _T_9374 | _T_9207; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9209 = _T_4681 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9376 = _T_9375 | _T_9209; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9211 = _T_4685 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9377 = _T_9376 | _T_9211; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9213 = _T_4689 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9378 = _T_9377 | _T_9213; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9215 = _T_4693 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9379 = _T_9378 | _T_9215; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9217 = _T_4697 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9380 = _T_9379 | _T_9217; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9219 = _T_4701 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9381 = _T_9380 | _T_9219; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9221 = _T_4705 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9382 = _T_9381 | _T_9221; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9223 = _T_4709 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9383 = _T_9382 | _T_9223; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9225 = _T_4713 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9384 = _T_9383 | _T_9225; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9227 = _T_4717 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9385 = _T_9384 | _T_9227; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9229 = _T_4721 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9386 = _T_9385 | _T_9229; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9231 = _T_4725 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9387 = _T_9386 | _T_9231; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9233 = _T_4729 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9388 = _T_9387 | _T_9233; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9235 = _T_4733 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9389 = _T_9388 | _T_9235; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9237 = _T_4737 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9390 = _T_9389 | _T_9237; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9239 = _T_4741 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9391 = _T_9390 | _T_9239; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9241 = _T_4745 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9392 = _T_9391 | _T_9241; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9243 = _T_4749 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9393 = _T_9392 | _T_9243; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9245 = _T_4753 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9394 = _T_9393 | _T_9245; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9247 = _T_4757 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9395 = _T_9394 | _T_9247; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9249 = _T_4761 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9396 = _T_9395 | _T_9249; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9251 = _T_4765 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9397 = _T_9396 | _T_9251; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9253 = _T_4769 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9398 = _T_9397 | _T_9253; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9255 = _T_4773 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9399 = _T_9398 | _T_9255; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9257 = _T_4777 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9400 = _T_9399 | _T_9257; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9259 = _T_4781 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9401 = _T_9400 | _T_9259; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9261 = _T_4785 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9402 = _T_9401 | _T_9261; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9263 = _T_4789 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9403 = _T_9402 | _T_9263; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9265 = _T_4793 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9404 = _T_9403 | _T_9265; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9267 = _T_4797 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9405 = _T_9404 | _T_9267; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9269 = _T_4801 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9406 = _T_9405 | _T_9269; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9271 = _T_4805 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9407 = _T_9406 | _T_9271; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9273 = _T_4809 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9408 = _T_9407 | _T_9273; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9275 = _T_4813 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9409 = _T_9408 | _T_9275; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9277 = _T_4817 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9410 = _T_9409 | _T_9277; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9279 = _T_4821 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9411 = _T_9410 | _T_9279; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9281 = _T_4825 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9412 = _T_9411 | _T_9281; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9283 = _T_4829 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9413 = _T_9412 | _T_9283; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9285 = _T_4833 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9414 = _T_9413 | _T_9285; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9287 = _T_4837 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9415 = _T_9414 | _T_9287; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9289 = _T_4841 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9416 = _T_9415 | _T_9289; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8652 = _T_4333 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 796:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8654 = _T_4337 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8907 = _T_8652 | _T_8654; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8656 = _T_4341 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8908 = _T_8907 | _T_8656; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8658 = _T_4345 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8909 = _T_8908 | _T_8658; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8660 = _T_4349 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8910 = _T_8909 | _T_8660; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8662 = _T_4353 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8911 = _T_8910 | _T_8662; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8664 = _T_4357 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8912 = _T_8911 | _T_8664; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8666 = _T_4361 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8913 = _T_8912 | _T_8666; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8668 = _T_4365 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8914 = _T_8913 | _T_8668; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8670 = _T_4369 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8915 = _T_8914 | _T_8670; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8672 = _T_4373 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8916 = _T_8915 | _T_8672; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8674 = _T_4377 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8917 = _T_8916 | _T_8674; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8676 = _T_4381 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8918 = _T_8917 | _T_8676; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8678 = _T_4385 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8919 = _T_8918 | _T_8678; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8680 = _T_4389 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8920 = _T_8919 | _T_8680; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8682 = _T_4393 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8921 = _T_8920 | _T_8682; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8684 = _T_4397 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8922 = _T_8921 | _T_8684; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8686 = _T_4401 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8923 = _T_8922 | _T_8686; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8688 = _T_4405 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8924 = _T_8923 | _T_8688; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8690 = _T_4409 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8925 = _T_8924 | _T_8690; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8692 = _T_4413 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8926 = _T_8925 | _T_8692; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8694 = _T_4417 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8927 = _T_8926 | _T_8694; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8696 = _T_4421 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8928 = _T_8927 | _T_8696; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8698 = _T_4425 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8929 = _T_8928 | _T_8698; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8700 = _T_4429 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8930 = _T_8929 | _T_8700; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8702 = _T_4433 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8931 = _T_8930 | _T_8702; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8704 = _T_4437 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8932 = _T_8931 | _T_8704; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8706 = _T_4441 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8933 = _T_8932 | _T_8706; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8708 = _T_4445 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8934 = _T_8933 | _T_8708; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8710 = _T_4449 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8935 = _T_8934 | _T_8710; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_8712 = _T_4453 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8936 = _T_8935 | _T_8712; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_8714 = _T_4457 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8937 = _T_8936 | _T_8714; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_8716 = _T_4461 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8938 = _T_8937 | _T_8716; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_8718 = _T_4465 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8939 = _T_8938 | _T_8718; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_8720 = _T_4469 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8940 = _T_8939 | _T_8720; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_8722 = _T_4473 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8941 = _T_8940 | _T_8722; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_8724 = _T_4477 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8942 = _T_8941 | _T_8724; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_8726 = _T_4481 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8943 = _T_8942 | _T_8726; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_8728 = _T_4485 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8944 = _T_8943 | _T_8728; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_8730 = _T_4489 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8945 = _T_8944 | _T_8730; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_8732 = _T_4493 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8946 = _T_8945 | _T_8732; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_8734 = _T_4497 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8947 = _T_8946 | _T_8734; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_8736 = _T_4501 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8948 = _T_8947 | _T_8736; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_8738 = _T_4505 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8949 = _T_8948 | _T_8738; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_8740 = _T_4509 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8950 = _T_8949 | _T_8740; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_8742 = _T_4513 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8951 = _T_8950 | _T_8742; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_8744 = _T_4517 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8952 = _T_8951 | _T_8744; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_8746 = _T_4521 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8953 = _T_8952 | _T_8746; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_8748 = _T_4525 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8954 = _T_8953 | _T_8748; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_8750 = _T_4529 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8955 = _T_8954 | _T_8750; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_8752 = _T_4533 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8956 = _T_8955 | _T_8752; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_8754 = _T_4537 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8957 = _T_8956 | _T_8754; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_8756 = _T_4541 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8958 = _T_8957 | _T_8756; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_8758 = _T_4545 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8959 = _T_8958 | _T_8758; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_8760 = _T_4549 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8960 = _T_8959 | _T_8760; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_8762 = _T_4553 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8961 = _T_8960 | _T_8762; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_8764 = _T_4557 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8962 = _T_8961 | _T_8764; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_8766 = _T_4561 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8963 = _T_8962 | _T_8766; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_8768 = _T_4565 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8964 = _T_8963 | _T_8768; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_8770 = _T_4569 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8965 = _T_8964 | _T_8770; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_8772 = _T_4573 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8966 = _T_8965 | _T_8772; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_8774 = _T_4577 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8967 = _T_8966 | _T_8774; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_8776 = _T_4581 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8968 = _T_8967 | _T_8776; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_8778 = _T_4585 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8969 = _T_8968 | _T_8778; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_8780 = _T_4589 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8970 = _T_8969 | _T_8780; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_8782 = _T_4593 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8971 = _T_8970 | _T_8782; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_8784 = _T_4597 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8972 = _T_8971 | _T_8784; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_8786 = _T_4601 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8973 = _T_8972 | _T_8786; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_8788 = _T_4605 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8974 = _T_8973 | _T_8788; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_8790 = _T_4609 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8975 = _T_8974 | _T_8790; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_8792 = _T_4613 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8976 = _T_8975 | _T_8792; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_8794 = _T_4617 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8977 = _T_8976 | _T_8794; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_8796 = _T_4621 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8978 = _T_8977 | _T_8796; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_8798 = _T_4625 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8979 = _T_8978 | _T_8798; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_8800 = _T_4629 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8980 = _T_8979 | _T_8800; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_8802 = _T_4633 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8981 = _T_8980 | _T_8802; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_8804 = _T_4637 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8982 = _T_8981 | _T_8804; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_8806 = _T_4641 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8983 = _T_8982 | _T_8806; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_8808 = _T_4645 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8984 = _T_8983 | _T_8808; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_8810 = _T_4649 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8985 = _T_8984 | _T_8810; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_8812 = _T_4653 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8986 = _T_8985 | _T_8812; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_8814 = _T_4657 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8987 = _T_8986 | _T_8814; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_8816 = _T_4661 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8988 = _T_8987 | _T_8816; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_8818 = _T_4665 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8989 = _T_8988 | _T_8818; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_8820 = _T_4669 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8990 = _T_8989 | _T_8820; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_8822 = _T_4673 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8991 = _T_8990 | _T_8822; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_8824 = _T_4677 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8992 = _T_8991 | _T_8824; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_8826 = _T_4681 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8993 = _T_8992 | _T_8826; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_8828 = _T_4685 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8994 = _T_8993 | _T_8828; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_8830 = _T_4689 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8995 = _T_8994 | _T_8830; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_8832 = _T_4693 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8996 = _T_8995 | _T_8832; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_8834 = _T_4697 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8997 = _T_8996 | _T_8834; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_8836 = _T_4701 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8998 = _T_8997 | _T_8836; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_8838 = _T_4705 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_8999 = _T_8998 | _T_8838; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_8840 = _T_4709 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9000 = _T_8999 | _T_8840; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_8842 = _T_4713 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9001 = _T_9000 | _T_8842; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_8844 = _T_4717 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9002 = _T_9001 | _T_8844; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_8846 = _T_4721 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9003 = _T_9002 | _T_8846; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_8848 = _T_4725 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9004 = _T_9003 | _T_8848; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_8850 = _T_4729 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9005 = _T_9004 | _T_8850; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_8852 = _T_4733 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9006 = _T_9005 | _T_8852; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_8854 = _T_4737 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9007 = _T_9006 | _T_8854; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_8856 = _T_4741 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9008 = _T_9007 | _T_8856; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_8858 = _T_4745 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9009 = _T_9008 | _T_8858; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_8860 = _T_4749 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9010 = _T_9009 | _T_8860; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_8862 = _T_4753 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9011 = _T_9010 | _T_8862; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_8864 = _T_4757 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9012 = _T_9011 | _T_8864; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_8866 = _T_4761 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9013 = _T_9012 | _T_8866; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_8868 = _T_4765 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9014 = _T_9013 | _T_8868; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_8870 = _T_4769 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9015 = _T_9014 | _T_8870; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_8872 = _T_4773 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9016 = _T_9015 | _T_8872; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_8874 = _T_4777 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9017 = _T_9016 | _T_8874; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_8876 = _T_4781 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9018 = _T_9017 | _T_8876; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_8878 = _T_4785 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9019 = _T_9018 | _T_8878; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_8880 = _T_4789 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9020 = _T_9019 | _T_8880; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_8882 = _T_4793 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9021 = _T_9020 | _T_8882; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_8884 = _T_4797 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9022 = _T_9021 | _T_8884; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_8886 = _T_4801 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9023 = _T_9022 | _T_8886; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_8888 = _T_4805 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9024 = _T_9023 | _T_8888; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_8890 = _T_4809 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9025 = _T_9024 | _T_8890; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_8892 = _T_4813 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9026 = _T_9025 | _T_8892; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_8894 = _T_4817 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9027 = _T_9026 | _T_8894; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_8896 = _T_4821 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9028 = _T_9027 | _T_8896; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_8898 = _T_4825 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9029 = _T_9028 | _T_8898; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_8900 = _T_4829 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9030 = _T_9029 | _T_8900; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_8902 = _T_4833 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9031 = _T_9030 | _T_8902; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_8904 = _T_4837 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9032 = _T_9031 | _T_8904; // @[el2_ifu_mem_ctl.scala 796:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_8906 = _T_4841 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 796:10]
  wire  _T_9033 = _T_9032 | _T_8906; // @[el2_ifu_mem_ctl.scala 796:91]
  wire [1:0] ic_tag_valid_unq = {_T_9416,_T_9033}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 867:54]
  wire [1:0] _T_9455 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9456 = ic_debug_way_ff & _T_9455; // @[el2_ifu_mem_ctl.scala 850:67]
  wire [1:0] _T_9457 = ic_tag_valid_unq & _T_9456; // @[el2_ifu_mem_ctl.scala 850:48]
  wire  ic_debug_tag_val_rd_out = |_T_9457; // @[el2_ifu_mem_ctl.scala 850:115]
  wire [65:0] _T_1200 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1201; // @[el2_ifu_mem_ctl.scala 400:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2529; // @[el2_ifu_mem_ctl.scala 410:80]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_309; // @[el2_ifu_mem_ctl.scala 428:38]
  wire [1:0] _T_1265 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 432:8]
  wire [7:0] _T_1346 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1351 = ic_miss_buff_data_error[0] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  _T_2597 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 661:47]
  wire  _T_2598 = _T_2597 & _T_14; // @[el2_ifu_mem_ctl.scala 661:50]
  wire  bus_ifu_wr_data_error = _T_2598 & miss_pending; // @[el2_ifu_mem_ctl.scala 661:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1351; // @[el2_ifu_mem_ctl.scala 452:72]
  wire  _T_1355 = ic_miss_buff_data_error[1] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1355; // @[el2_ifu_mem_ctl.scala 452:72]
  wire  _T_1359 = ic_miss_buff_data_error[2] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1359; // @[el2_ifu_mem_ctl.scala 452:72]
  wire  _T_1363 = ic_miss_buff_data_error[3] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1363; // @[el2_ifu_mem_ctl.scala 452:72]
  wire  _T_1367 = ic_miss_buff_data_error[4] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1367; // @[el2_ifu_mem_ctl.scala 452:72]
  wire  _T_1371 = ic_miss_buff_data_error[5] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1371; // @[el2_ifu_mem_ctl.scala 452:72]
  wire  _T_1375 = ic_miss_buff_data_error[6] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1375; // @[el2_ifu_mem_ctl.scala 452:72]
  wire  _T_1379 = ic_miss_buff_data_error[7] & _T_1317; // @[el2_ifu_mem_ctl.scala 453:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1379; // @[el2_ifu_mem_ctl.scala 452:72]
  wire [7:0] _T_1386 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2405 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2413 = _T_7 & _T_309; // @[el2_ifu_mem_ctl.scala 531:65]
  wire  _T_2414 = _T_2413 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 531:88]
  wire  _T_2416 = _T_2414 & _T_2525; // @[el2_ifu_mem_ctl.scala 531:112]
  wire  _T_2417 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2418 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 536:50]
  wire  _T_2420 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2426 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2428 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2426 | _T_2428; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2420 ? _T_2418 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2417 ? _T_2418 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2405 ? _T_2416 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2405 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2419 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 537:56]
  wire  _GEN_43 = _T_2417 & _T_2419; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2405 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_2407 = io_ic_error_start & _T_309; // @[el2_ifu_mem_ctl.scala 530:87]
  wire  _T_2421 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 540:54]
  wire  _T_2422 = _T_2421 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 540:84]
  wire  _T_2431 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 561:66]
  wire  _T_2432 = io_dec_tlu_flush_err_wb & _T_2431; // @[el2_ifu_mem_ctl.scala 561:52]
  wire  _T_2434 = _T_2432 & _T_2525; // @[el2_ifu_mem_ctl.scala 561:81]
  wire  _T_2436 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 564:59]
  wire  _T_2437 = _T_2436 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 564:86]
  wire  _T_2451 = _T_2436 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 567:81]
  wire  _T_2452 = _T_2451 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 567:103]
  wire  _T_2453 = _T_2452 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 567:126]
  wire  _T_2473 = _T_2451 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 574:103]
  wire  _T_2480 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 579:62]
  wire  _T_2481 = io_dec_tlu_flush_lower_wb & _T_2480; // @[el2_ifu_mem_ctl.scala 579:60]
  wire  _T_2482 = _T_2481 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 579:88]
  wire  _T_2483 = _T_2482 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 579:115]
  wire  _GEN_50 = _T_2479 & _T_2437; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_2462 ? _T_2473 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_2435 ? _T_2453 : _GEN_53; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2430 ? _T_2434 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2493 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 595:64]
  wire  _T_2495 = _T_2493 & _T_2525; // @[el2_ifu_mem_ctl.scala 595:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2497 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 595:133]
  wire  _T_2498 = _T_2497 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 595:164]
  wire  _T_2499 = _T_2498 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 595:184]
  wire  _T_2500 = _T_2499 & miss_pending; // @[el2_ifu_mem_ctl.scala 595:204]
  wire  _T_2501 = ~_T_2500; // @[el2_ifu_mem_ctl.scala 595:112]
  wire  ifc_bus_ic_req_ff_in = _T_2495 & _T_2501; // @[el2_ifu_mem_ctl.scala 595:110]
  wire  _T_2502 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 596:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 627:45]
  wire  _T_2519 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 630:35]
  wire  _T_2520 = _T_2519 & miss_pending; // @[el2_ifu_mem_ctl.scala 630:53]
  wire  bus_cmd_sent = _T_2520 & _T_2525; // @[el2_ifu_mem_ctl.scala 630:68]
  wire [2:0] _T_2510 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2512 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2514 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 628:51]
  wire  _T_2543 = last_data_recieved_ff & _T_1317; // @[el2_ifu_mem_ctl.scala 638:114]
  wire  last_data_recieved_in = _T_2526 | _T_2543; // @[el2_ifu_mem_ctl.scala 638:89]
  wire [2:0] _T_2549 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 643:45]
  wire  _T_2552 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 644:81]
  wire  _T_2553 = _T_2552 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 644:97]
  wire  _T_2555 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 646:48]
  wire  _T_2556 = _T_2555 & miss_pending; // @[el2_ifu_mem_ctl.scala 646:68]
  wire  bus_inc_cmd_beat_cnt = _T_2556 & _T_2525; // @[el2_ifu_mem_ctl.scala 646:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 648:57]
  wire  _T_2560 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 649:31]
  wire  _T_2562 = ic_act_miss_f | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 649:87]
  wire  _T_2563 = ~_T_2562; // @[el2_ifu_mem_ctl.scala 649:55]
  wire  bus_hold_cmd_beat_cnt = _T_2560 & _T_2563; // @[el2_ifu_mem_ctl.scala 649:53]
  wire  _T_2564 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 650:46]
  wire  bus_cmd_beat_en = _T_2564 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 650:62]
  wire [2:0] _T_2567 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 652:46]
  wire [2:0] _T_2569 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2570 = bus_inc_cmd_beat_cnt ? _T_2567 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2571 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2573 = _T_2569 | _T_2570; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2573 | _T_2571; // @[Mux.scala 27:72]
  wire  _T_2577 = _T_2553 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 653:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 664:62]
  wire  _T_2605 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 669:50]
  wire  _T_2606 = io_ifc_dma_access_ok & _T_2605; // @[el2_ifu_mem_ctl.scala 669:47]
  wire  _T_2607 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 669:70]
  wire  ifc_dma_access_ok_d = _T_2606 & _T_2607; // @[el2_ifu_mem_ctl.scala 669:68]
  wire  _T_2611 = _T_2606 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 670:72]
  wire  _T_2612 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 670:111]
  wire  _T_2613 = _T_2611 & _T_2612; // @[el2_ifu_mem_ctl.scala 670:97]
  wire  iccm_ready = _T_2613 & _T_2607; // @[el2_ifu_mem_ctl.scala 670:127]
  wire  _T_2616 = iccm_ready & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 673:40]
  wire  _T_2617 = _T_2616 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 673:58]
  wire  _T_2620 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 674:60]
  wire  _T_2621 = _T_2616 & _T_2620; // @[el2_ifu_mem_ctl.scala 674:58]
  wire  _T_2622 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 674:104]
  wire [2:0] _T_2627 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2733 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2742 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2733}; // @[el2_lib.scala 268:22]
  wire  _T_2743 = ^_T_2742; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2751 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2760 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2751}; // @[el2_lib.scala 268:39]
  wire  _T_2761 = ^_T_2760; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2769 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2778 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2769}; // @[el2_lib.scala 268:56]
  wire  _T_2779 = ^_T_2778; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2785 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2793 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2785}; // @[el2_lib.scala 268:73]
  wire  _T_2794 = ^_T_2793; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2808 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2785}; // @[el2_lib.scala 268:90]
  wire  _T_2809 = ^_T_2808; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2814 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2815 = ^_T_2814; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2820 = {_T_2743,_T_2761,_T_2779,_T_2794,_T_2809,_T_2815}; // @[Cat.scala 29:58]
  wire  _T_2821 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2822 = ^_T_2820; // @[el2_lib.scala 269:23]
  wire  _T_2823 = _T_2821 ^ _T_2822; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2929 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2938 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2929}; // @[el2_lib.scala 268:22]
  wire  _T_2939 = ^_T_2938; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2947 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2956 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2947}; // @[el2_lib.scala 268:39]
  wire  _T_2957 = ^_T_2956; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2965 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2974 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2965}; // @[el2_lib.scala 268:56]
  wire  _T_2975 = ^_T_2974; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2981 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2989 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2981}; // @[el2_lib.scala 268:73]
  wire  _T_2990 = ^_T_2989; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3004 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2981}; // @[el2_lib.scala 268:90]
  wire  _T_3005 = ^_T_3004; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3010 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3011 = ^_T_3010; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3016 = {_T_2939,_T_2957,_T_2975,_T_2990,_T_3005,_T_3011}; // @[Cat.scala 29:58]
  wire  _T_3017 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3018 = ^_T_3016; // @[el2_lib.scala 269:23]
  wire  _T_3019 = _T_3017 ^ _T_3018; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3020 = {_T_3019,_T_2939,_T_2957,_T_2975,_T_2990,_T_3005,_T_3011}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2823,_T_2743,_T_2761,_T_2779,_T_2794,_T_2809,_T_2815,_T_3020}; // @[Cat.scala 29:58]
  wire  _T_3022 = ~_T_2616; // @[el2_ifu_mem_ctl.scala 679:45]
  wire  _T_3023 = iccm_correct_ecc & _T_3022; // @[el2_ifu_mem_ctl.scala 679:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3024 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3031 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 693:53]
  wire  _T_3363 = _T_3275[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3361 = _T_3275[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3359 = _T_3275[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3357 = _T_3275[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3355 = _T_3275[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3353 = _T_3275[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3351 = _T_3275[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3349 = _T_3275[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3347 = _T_3275[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3345 = _T_3275[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3421 = {_T_3363,_T_3361,_T_3359,_T_3357,_T_3355,_T_3353,_T_3351,_T_3349,_T_3347,_T_3345}; // @[el2_lib.scala 310:69]
  wire  _T_3343 = _T_3275[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3341 = _T_3275[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3339 = _T_3275[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3337 = _T_3275[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3335 = _T_3275[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3333 = _T_3275[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3331 = _T_3275[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3329 = _T_3275[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3327 = _T_3275[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3325 = _T_3275[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3412 = {_T_3343,_T_3341,_T_3339,_T_3337,_T_3335,_T_3333,_T_3331,_T_3329,_T_3327,_T_3325}; // @[el2_lib.scala 310:69]
  wire  _T_3323 = _T_3275[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3321 = _T_3275[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3319 = _T_3275[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3317 = _T_3275[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3315 = _T_3275[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3313 = _T_3275[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3311 = _T_3275[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3309 = _T_3275[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3307 = _T_3275[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3305 = _T_3275[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3402 = {_T_3323,_T_3321,_T_3319,_T_3317,_T_3315,_T_3313,_T_3311,_T_3309,_T_3307,_T_3305}; // @[el2_lib.scala 310:69]
  wire  _T_3303 = _T_3275[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3301 = _T_3275[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3299 = _T_3275[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3297 = _T_3275[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3295 = _T_3275[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3293 = _T_3275[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3291 = _T_3275[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3289 = _T_3275[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3287 = _T_3275[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3403 = {_T_3402,_T_3303,_T_3301,_T_3299,_T_3297,_T_3295,_T_3293,_T_3291,_T_3289,_T_3287}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3423 = {_T_3421,_T_3412,_T_3403}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3378 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3384 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3378}; // @[Cat.scala 29:58]
  wire [38:0] _T_3424 = _T_3423 ^ _T_3384; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3425 = _T_3279 ? _T_3424 : _T_3384; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3425[37:32],_T_3425[30:16],_T_3425[14:8],_T_3425[6:4],_T_3425[2]}; // @[Cat.scala 29:58]
  wire  _T_3748 = _T_3660[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3746 = _T_3660[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3744 = _T_3660[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3742 = _T_3660[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3740 = _T_3660[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3738 = _T_3660[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3736 = _T_3660[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3734 = _T_3660[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3732 = _T_3660[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3730 = _T_3660[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3806 = {_T_3748,_T_3746,_T_3744,_T_3742,_T_3740,_T_3738,_T_3736,_T_3734,_T_3732,_T_3730}; // @[el2_lib.scala 310:69]
  wire  _T_3728 = _T_3660[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3726 = _T_3660[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3724 = _T_3660[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3722 = _T_3660[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3720 = _T_3660[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3718 = _T_3660[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3716 = _T_3660[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3714 = _T_3660[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3712 = _T_3660[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3710 = _T_3660[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3797 = {_T_3728,_T_3726,_T_3724,_T_3722,_T_3720,_T_3718,_T_3716,_T_3714,_T_3712,_T_3710}; // @[el2_lib.scala 310:69]
  wire  _T_3708 = _T_3660[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3706 = _T_3660[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3704 = _T_3660[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3702 = _T_3660[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3700 = _T_3660[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3698 = _T_3660[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3696 = _T_3660[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3694 = _T_3660[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3692 = _T_3660[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3690 = _T_3660[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3787 = {_T_3708,_T_3706,_T_3704,_T_3702,_T_3700,_T_3698,_T_3696,_T_3694,_T_3692,_T_3690}; // @[el2_lib.scala 310:69]
  wire  _T_3688 = _T_3660[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3686 = _T_3660[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3684 = _T_3660[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3682 = _T_3660[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3680 = _T_3660[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3678 = _T_3660[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3676 = _T_3660[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3674 = _T_3660[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3672 = _T_3660[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3788 = {_T_3787,_T_3688,_T_3686,_T_3684,_T_3682,_T_3680,_T_3678,_T_3676,_T_3674,_T_3672}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3808 = {_T_3806,_T_3797,_T_3788}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3763 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3769 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3763}; // @[Cat.scala 29:58]
  wire [38:0] _T_3809 = _T_3808 ^ _T_3769; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3810 = _T_3664 ? _T_3809 : _T_3769; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3810[37:32],_T_3810[30:16],_T_3810[14:8],_T_3810[6:4],_T_3810[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 685:35]
  wire  _T_3283 = ~_T_3275[6]; // @[el2_lib.scala 303:55]
  wire  _T_3284 = _T_3277 & _T_3283; // @[el2_lib.scala 303:53]
  wire  _T_3668 = ~_T_3660[6]; // @[el2_lib.scala 303:55]
  wire  _T_3669 = _T_3662 & _T_3668; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3284,_T_3669}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 687:53]
  wire [63:0] _T_3035 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3036 = {iccm_dma_rdata_1_muxed,_T_3425[37:32],_T_3425[30:16],_T_3425[14:8],_T_3425[6:4],_T_3425[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 689:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 690:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 695:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 699:70]
  wire  _T_3041 = _T_2616 & _T_2605; // @[el2_ifu_mem_ctl.scala 702:65]
  wire  _T_3044 = _T_3022 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 703:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3045 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3047 = _T_3044 ? {{1'd0}, _T_3045} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 703:8]
  wire [31:0] _T_3048 = _T_3041 ? io_dma_mem_addr : {{16'd0}, _T_3047}; // @[el2_ifu_mem_ctl.scala 702:25]
  wire  _T_3437 = _T_3275 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3438 = _T_3425[38] ^ _T_3437; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3438,_T_3425[31],_T_3425[15],_T_3425[7],_T_3425[3],_T_3425[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3822 = _T_3660 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3823 = _T_3810[38] ^ _T_3822; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3823,_T_3810[31],_T_3810[15],_T_3810[7],_T_3810[3],_T_3810[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3839 = _T_4 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 715:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 717:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 718:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 726:62]
  wire  _T_3847 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 720:76]
  wire  _T_3848 = io_iccm_rd_ecc_single_err & _T_3847; // @[el2_ifu_mem_ctl.scala 720:74]
  wire  _T_3850 = _T_3848 & _T_309; // @[el2_ifu_mem_ctl.scala 720:104]
  wire  iccm_ecc_write_status = _T_3850 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 720:127]
  wire  _T_3851 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 721:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3851 & _T_309; // @[el2_ifu_mem_ctl.scala 721:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 725:51]
  wire [13:0] _T_3856 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 724:102]
  wire [38:0] _T_3860 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3865 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 729:41]
  wire  _T_3866 = io_ifc_fetch_req_bf & _T_3865; // @[el2_ifu_mem_ctl.scala 729:39]
  wire  _T_3867 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 729:72]
  wire  _T_3868 = _T_3866 & _T_3867; // @[el2_ifu_mem_ctl.scala 729:70]
  wire  _T_3870 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 730:34]
  wire  _T_3871 = _T_2217 & _T_3870; // @[el2_ifu_mem_ctl.scala 730:32]
  wire  _T_3874 = _T_2232 & _T_3870; // @[el2_ifu_mem_ctl.scala 731:37]
  wire  _T_3875 = _T_3871 | _T_3874; // @[el2_ifu_mem_ctl.scala 730:88]
  wire  _T_3876 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 732:19]
  wire  _T_3878 = _T_3876 & _T_3870; // @[el2_ifu_mem_ctl.scala 732:41]
  wire  _T_3879 = _T_3875 | _T_3878; // @[el2_ifu_mem_ctl.scala 731:88]
  wire  _T_3880 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 733:19]
  wire  _T_3882 = _T_3880 & _T_3870; // @[el2_ifu_mem_ctl.scala 733:35]
  wire  _T_3883 = _T_3879 | _T_3882; // @[el2_ifu_mem_ctl.scala 732:88]
  wire  _T_3886 = _T_2231 & _T_3870; // @[el2_ifu_mem_ctl.scala 734:38]
  wire  _T_3887 = _T_3883 | _T_3886; // @[el2_ifu_mem_ctl.scala 733:88]
  wire  _T_3889 = _T_2232 & miss_state_en; // @[el2_ifu_mem_ctl.scala 735:37]
  wire  _T_3890 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 735:71]
  wire  _T_3891 = _T_3889 & _T_3890; // @[el2_ifu_mem_ctl.scala 735:54]
  wire  _T_3892 = _T_3887 | _T_3891; // @[el2_ifu_mem_ctl.scala 734:57]
  wire  _T_3893 = ~_T_3892; // @[el2_ifu_mem_ctl.scala 730:5]
  wire  _T_3894 = _T_3868 & _T_3893; // @[el2_ifu_mem_ctl.scala 729:96]
  wire  _T_3895 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 736:28]
  wire  _T_3897 = _T_3895 & _T_3865; // @[el2_ifu_mem_ctl.scala 736:50]
  wire  _T_3899 = _T_3897 & _T_3867; // @[el2_ifu_mem_ctl.scala 736:81]
  wire  _T_3908 = ~_T_100; // @[el2_ifu_mem_ctl.scala 739:106]
  wire  _T_3909 = _T_2217 & _T_3908; // @[el2_ifu_mem_ctl.scala 739:104]
  wire  _T_3910 = _T_2232 | _T_3909; // @[el2_ifu_mem_ctl.scala 739:77]
  wire  _T_3914 = ~_T_53; // @[el2_ifu_mem_ctl.scala 739:172]
  wire  _T_3915 = _T_3910 & _T_3914; // @[el2_ifu_mem_ctl.scala 739:170]
  wire  _T_3916 = ~_T_3915; // @[el2_ifu_mem_ctl.scala 739:44]
  wire  _T_3920 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 742:64]
  wire  _T_3921 = ~_T_3920; // @[el2_ifu_mem_ctl.scala 742:50]
  wire  _T_3922 = _T_268 & _T_3921; // @[el2_ifu_mem_ctl.scala 742:48]
  wire  _T_3923 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 742:81]
  wire  ic_valid = _T_3922 & _T_3923; // @[el2_ifu_mem_ctl.scala 742:79]
  wire  _T_3925 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 743:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 746:14]
  wire  _T_3928 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 749:74]
  wire  _T_9438 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 827:45]
  wire  way_status_wr_en = _T_9438 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 827:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3928; // @[el2_ifu_mem_ctl.scala 749:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 751:14]
  wire [2:0] _T_3932 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 755:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 823:41]
  wire  way_status_new = _T_9438 | way_status_hit_new; // @[el2_ifu_mem_ctl.scala 826:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 757:14]
  wire  _T_3949 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3950 = _T_3949 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_3952 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3953 = _T_3952 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_3955 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3956 = _T_3955 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_3958 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3959 = _T_3958 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_3961 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3962 = _T_3961 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_3964 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3965 = _T_3964 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_3967 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3968 = _T_3967 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_3970 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 764:65]
  wire  _T_3971 = _T_3970 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 764:73]
  wire  _T_9443 = _T_92 & miss_pending; // @[el2_ifu_mem_ctl.scala 830:108]
  wire  bus_wren_last_0 = _T_9443 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 830:123]
  wire  _T_9446 = bus_wren_last_0 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 832:73]
  wire [1:0] ifu_tag_wren = {1'h0,_T_9446}; // @[Cat.scala 29:58]
  wire [1:0] _T_9481 = _T_3928 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9481 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 863:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 774:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 776:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 780:14]
  wire  _T_4980 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 784:82]
  wire  _T_4982 = _T_4980 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_4984 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 785:74]
  wire  _T_4986 = _T_4984 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_4987 = _T_4982 | _T_4986; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_4988 = _T_4987 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire  _T_4992 = _T_4980 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_4996 = _T_4984 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_4997 = _T_4992 | _T_4996; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_4998 = _T_4997 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire [1:0] tag_valid_clken_0 = {_T_4988,_T_4998}; // @[Cat.scala 29:58]
  wire  _T_5000 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 784:82]
  wire  _T_5002 = _T_5000 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_5004 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 785:74]
  wire  _T_5006 = _T_5004 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_5007 = _T_5002 | _T_5006; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_5008 = _T_5007 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire  _T_5012 = _T_5000 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_5016 = _T_5004 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_5017 = _T_5012 | _T_5016; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_5018 = _T_5017 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire [1:0] tag_valid_clken_1 = {_T_5008,_T_5018}; // @[Cat.scala 29:58]
  wire  _T_5020 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 784:82]
  wire  _T_5022 = _T_5020 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_5024 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 785:74]
  wire  _T_5026 = _T_5024 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_5027 = _T_5022 | _T_5026; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_5028 = _T_5027 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire  _T_5032 = _T_5020 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_5036 = _T_5024 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_5037 = _T_5032 | _T_5036; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_5038 = _T_5037 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire [1:0] tag_valid_clken_2 = {_T_5028,_T_5038}; // @[Cat.scala 29:58]
  wire  _T_5040 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 784:82]
  wire  _T_5042 = _T_5040 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_5044 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 785:74]
  wire  _T_5046 = _T_5044 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_5047 = _T_5042 | _T_5046; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_5048 = _T_5047 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire  _T_5052 = _T_5040 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 784:91]
  wire  _T_5056 = _T_5044 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 785:83]
  wire  _T_5057 = _T_5052 | _T_5056; // @[el2_ifu_mem_ctl.scala 784:113]
  wire  _T_5058 = _T_5057 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 785:106]
  wire [1:0] tag_valid_clken_3 = {_T_5048,_T_5058}; // @[Cat.scala 29:58]
  wire  _T_5069 = ic_valid_ff & _T_187; // @[el2_ifu_mem_ctl.scala 791:31]
  wire  _T_5070 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 791:58]
  wire  _T_5071 = _T_5069 & _T_5070; // @[el2_ifu_mem_ctl.scala 791:56]
  wire  _T_5074 = _T_4333 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5075 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5077 = _T_5075 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5078 = _T_5074 | _T_5077; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5088 = _T_4337 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5089 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5091 = _T_5089 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5092 = _T_5088 | _T_5091; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5102 = _T_4341 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5103 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5105 = _T_5103 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5106 = _T_5102 | _T_5105; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5116 = _T_4345 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5117 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5119 = _T_5117 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5120 = _T_5116 | _T_5119; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5130 = _T_4349 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5131 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5133 = _T_5131 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5134 = _T_5130 | _T_5133; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5144 = _T_4353 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5145 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5147 = _T_5145 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5148 = _T_5144 | _T_5147; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5158 = _T_4357 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5159 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5161 = _T_5159 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5162 = _T_5158 | _T_5161; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5172 = _T_4361 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5173 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5175 = _T_5173 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5176 = _T_5172 | _T_5175; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5186 = _T_4365 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5187 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5189 = _T_5187 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5190 = _T_5186 | _T_5189; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5200 = _T_4369 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5201 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5203 = _T_5201 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5204 = _T_5200 | _T_5203; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5214 = _T_4373 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5215 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5217 = _T_5215 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5218 = _T_5214 | _T_5217; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5228 = _T_4377 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5229 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5231 = _T_5229 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5232 = _T_5228 | _T_5231; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5242 = _T_4381 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5243 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5245 = _T_5243 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5246 = _T_5242 | _T_5245; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5256 = _T_4385 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5257 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5259 = _T_5257 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5260 = _T_5256 | _T_5259; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5270 = _T_4389 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5271 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5273 = _T_5271 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5274 = _T_5270 | _T_5273; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5284 = _T_4393 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5285 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5287 = _T_5285 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5288 = _T_5284 | _T_5287; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5298 = _T_4397 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5299 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5301 = _T_5299 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5302 = _T_5298 | _T_5301; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5312 = _T_4401 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5313 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5315 = _T_5313 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5316 = _T_5312 | _T_5315; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5326 = _T_4405 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5327 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5329 = _T_5327 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5330 = _T_5326 | _T_5329; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5340 = _T_4409 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5341 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5343 = _T_5341 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5344 = _T_5340 | _T_5343; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5354 = _T_4413 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5355 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5357 = _T_5355 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5358 = _T_5354 | _T_5357; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5368 = _T_4417 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5369 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5371 = _T_5369 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5372 = _T_5368 | _T_5371; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5382 = _T_4421 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5383 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5385 = _T_5383 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5386 = _T_5382 | _T_5385; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5396 = _T_4425 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5397 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5399 = _T_5397 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5400 = _T_5396 | _T_5399; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5410 = _T_4429 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5411 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5413 = _T_5411 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5414 = _T_5410 | _T_5413; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5424 = _T_4433 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5425 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5427 = _T_5425 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5428 = _T_5424 | _T_5427; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5438 = _T_4437 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5439 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5441 = _T_5439 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5442 = _T_5438 | _T_5441; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5452 = _T_4441 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5453 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5455 = _T_5453 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5456 = _T_5452 | _T_5455; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5466 = _T_4445 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5467 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5469 = _T_5467 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5470 = _T_5466 | _T_5469; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5480 = _T_4449 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5481 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5483 = _T_5481 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5484 = _T_5480 | _T_5483; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5494 = _T_4453 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5495 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5497 = _T_5495 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5498 = _T_5494 | _T_5497; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5508 = _T_4457 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5509 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5511 = _T_5509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5512 = _T_5508 | _T_5511; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5522 = _T_4333 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5525 = _T_5075 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5526 = _T_5522 | _T_5525; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5536 = _T_4337 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5539 = _T_5089 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5540 = _T_5536 | _T_5539; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5550 = _T_4341 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5553 = _T_5103 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5554 = _T_5550 | _T_5553; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5564 = _T_4345 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5567 = _T_5117 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5568 = _T_5564 | _T_5567; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5578 = _T_4349 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5581 = _T_5131 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5582 = _T_5578 | _T_5581; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5592 = _T_4353 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5595 = _T_5145 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5596 = _T_5592 | _T_5595; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5606 = _T_4357 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5609 = _T_5159 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5610 = _T_5606 | _T_5609; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5620 = _T_4361 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5623 = _T_5173 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5624 = _T_5620 | _T_5623; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5634 = _T_4365 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5637 = _T_5187 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5638 = _T_5634 | _T_5637; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5648 = _T_4369 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5651 = _T_5201 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5652 = _T_5648 | _T_5651; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5662 = _T_4373 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5665 = _T_5215 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5666 = _T_5662 | _T_5665; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5676 = _T_4377 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5679 = _T_5229 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5680 = _T_5676 | _T_5679; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5690 = _T_4381 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5693 = _T_5243 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5694 = _T_5690 | _T_5693; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5704 = _T_4385 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5707 = _T_5257 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5708 = _T_5704 | _T_5707; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5718 = _T_4389 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5721 = _T_5271 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5722 = _T_5718 | _T_5721; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5732 = _T_4393 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5735 = _T_5285 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5736 = _T_5732 | _T_5735; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5746 = _T_4397 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5749 = _T_5299 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5750 = _T_5746 | _T_5749; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5760 = _T_4401 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5763 = _T_5313 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5764 = _T_5760 | _T_5763; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5774 = _T_4405 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5777 = _T_5327 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5778 = _T_5774 | _T_5777; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5788 = _T_4409 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5791 = _T_5341 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5792 = _T_5788 | _T_5791; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5802 = _T_4413 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5805 = _T_5355 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5806 = _T_5802 | _T_5805; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5816 = _T_4417 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5819 = _T_5369 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5820 = _T_5816 | _T_5819; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5830 = _T_4421 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5833 = _T_5383 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5834 = _T_5830 | _T_5833; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5844 = _T_4425 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5847 = _T_5397 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5848 = _T_5844 | _T_5847; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5858 = _T_4429 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5861 = _T_5411 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5862 = _T_5858 | _T_5861; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5872 = _T_4433 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5875 = _T_5425 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5876 = _T_5872 | _T_5875; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5886 = _T_4437 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5889 = _T_5439 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5890 = _T_5886 | _T_5889; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5900 = _T_4441 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5903 = _T_5453 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5904 = _T_5900 | _T_5903; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5914 = _T_4445 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5917 = _T_5467 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5918 = _T_5914 | _T_5917; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5928 = _T_4449 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5931 = _T_5481 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5932 = _T_5928 | _T_5931; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5942 = _T_4453 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5945 = _T_5495 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5946 = _T_5942 | _T_5945; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5956 = _T_4457 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5959 = _T_5509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5960 = _T_5956 | _T_5959; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5970 = _T_4461 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5971 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5973 = _T_5971 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5974 = _T_5970 | _T_5973; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5984 = _T_4465 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5985 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_5987 = _T_5985 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_5988 = _T_5984 | _T_5987; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_5998 = _T_4469 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_5999 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6001 = _T_5999 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6002 = _T_5998 | _T_6001; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6012 = _T_4473 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6013 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6015 = _T_6013 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6016 = _T_6012 | _T_6015; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6026 = _T_4477 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6027 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6029 = _T_6027 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6030 = _T_6026 | _T_6029; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6040 = _T_4481 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6041 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6043 = _T_6041 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6044 = _T_6040 | _T_6043; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6054 = _T_4485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6055 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6057 = _T_6055 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6058 = _T_6054 | _T_6057; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6068 = _T_4489 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6069 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6071 = _T_6069 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6072 = _T_6068 | _T_6071; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6082 = _T_4493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6083 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6085 = _T_6083 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6086 = _T_6082 | _T_6085; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6096 = _T_4497 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6097 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6099 = _T_6097 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6100 = _T_6096 | _T_6099; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6110 = _T_4501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6111 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6113 = _T_6111 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6114 = _T_6110 | _T_6113; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6124 = _T_4505 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6125 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6127 = _T_6125 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6128 = _T_6124 | _T_6127; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6138 = _T_4509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6139 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6141 = _T_6139 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6142 = _T_6138 | _T_6141; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6152 = _T_4513 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6153 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6155 = _T_6153 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6156 = _T_6152 | _T_6155; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6166 = _T_4517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6167 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6169 = _T_6167 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6170 = _T_6166 | _T_6169; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6180 = _T_4521 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6181 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6183 = _T_6181 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6184 = _T_6180 | _T_6183; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6194 = _T_4525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6195 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6197 = _T_6195 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6198 = _T_6194 | _T_6197; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6208 = _T_4529 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6209 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6211 = _T_6209 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6212 = _T_6208 | _T_6211; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6222 = _T_4533 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6223 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6225 = _T_6223 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6226 = _T_6222 | _T_6225; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6236 = _T_4537 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6237 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6239 = _T_6237 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6240 = _T_6236 | _T_6239; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6250 = _T_4541 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6251 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6253 = _T_6251 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6254 = _T_6250 | _T_6253; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6264 = _T_4545 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6265 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6267 = _T_6265 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6268 = _T_6264 | _T_6267; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6278 = _T_4549 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6279 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6281 = _T_6279 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6282 = _T_6278 | _T_6281; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6292 = _T_4553 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6293 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6295 = _T_6293 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6296 = _T_6292 | _T_6295; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6306 = _T_4557 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6307 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6309 = _T_6307 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6310 = _T_6306 | _T_6309; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6320 = _T_4561 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6321 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6323 = _T_6321 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6324 = _T_6320 | _T_6323; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6334 = _T_4565 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6335 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6337 = _T_6335 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6338 = _T_6334 | _T_6337; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6348 = _T_4569 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6349 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6351 = _T_6349 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6352 = _T_6348 | _T_6351; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6362 = _T_4573 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6363 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6365 = _T_6363 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6366 = _T_6362 | _T_6365; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6376 = _T_4577 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6377 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6379 = _T_6377 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6380 = _T_6376 | _T_6379; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6390 = _T_4581 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6391 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6393 = _T_6391 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6394 = _T_6390 | _T_6393; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6404 = _T_4585 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6405 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6407 = _T_6405 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6408 = _T_6404 | _T_6407; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6418 = _T_4461 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6421 = _T_5971 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6422 = _T_6418 | _T_6421; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6432 = _T_4465 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6435 = _T_5985 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6436 = _T_6432 | _T_6435; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6446 = _T_4469 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6449 = _T_5999 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6450 = _T_6446 | _T_6449; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6460 = _T_4473 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6463 = _T_6013 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6464 = _T_6460 | _T_6463; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6474 = _T_4477 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6477 = _T_6027 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6478 = _T_6474 | _T_6477; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6488 = _T_4481 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6491 = _T_6041 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6492 = _T_6488 | _T_6491; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6502 = _T_4485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6505 = _T_6055 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6506 = _T_6502 | _T_6505; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6516 = _T_4489 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6519 = _T_6069 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6520 = _T_6516 | _T_6519; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6530 = _T_4493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6533 = _T_6083 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6534 = _T_6530 | _T_6533; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6544 = _T_4497 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6547 = _T_6097 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6548 = _T_6544 | _T_6547; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6558 = _T_4501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6561 = _T_6111 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6562 = _T_6558 | _T_6561; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6572 = _T_4505 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6575 = _T_6125 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6576 = _T_6572 | _T_6575; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6586 = _T_4509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6589 = _T_6139 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6590 = _T_6586 | _T_6589; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6600 = _T_4513 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6603 = _T_6153 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6604 = _T_6600 | _T_6603; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6614 = _T_4517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6617 = _T_6167 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6618 = _T_6614 | _T_6617; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6628 = _T_4521 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6631 = _T_6181 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6632 = _T_6628 | _T_6631; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6642 = _T_4525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6645 = _T_6195 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6646 = _T_6642 | _T_6645; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6656 = _T_4529 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6659 = _T_6209 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6660 = _T_6656 | _T_6659; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6670 = _T_4533 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6673 = _T_6223 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6674 = _T_6670 | _T_6673; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6684 = _T_4537 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6687 = _T_6237 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6688 = _T_6684 | _T_6687; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6698 = _T_4541 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6701 = _T_6251 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6702 = _T_6698 | _T_6701; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6712 = _T_4545 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6715 = _T_6265 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6716 = _T_6712 | _T_6715; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6726 = _T_4549 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6729 = _T_6279 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6730 = _T_6726 | _T_6729; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6740 = _T_4553 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6743 = _T_6293 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6744 = _T_6740 | _T_6743; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6754 = _T_4557 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6757 = _T_6307 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6758 = _T_6754 | _T_6757; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6768 = _T_4561 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6771 = _T_6321 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6772 = _T_6768 | _T_6771; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6782 = _T_4565 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6785 = _T_6335 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6786 = _T_6782 | _T_6785; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6796 = _T_4569 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6799 = _T_6349 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6800 = _T_6796 | _T_6799; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6810 = _T_4573 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6813 = _T_6363 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6814 = _T_6810 | _T_6813; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6824 = _T_4577 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6827 = _T_6377 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6828 = _T_6824 | _T_6827; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6838 = _T_4581 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6841 = _T_6391 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6842 = _T_6838 | _T_6841; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6852 = _T_4585 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6855 = _T_6405 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6856 = _T_6852 | _T_6855; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6866 = _T_4589 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6867 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6869 = _T_6867 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6870 = _T_6866 | _T_6869; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6880 = _T_4593 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6881 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6883 = _T_6881 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6884 = _T_6880 | _T_6883; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6894 = _T_4597 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6895 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6897 = _T_6895 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6898 = _T_6894 | _T_6897; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6908 = _T_4601 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6909 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6911 = _T_6909 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6912 = _T_6908 | _T_6911; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6922 = _T_4605 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6923 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6925 = _T_6923 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6926 = _T_6922 | _T_6925; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6936 = _T_4609 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6937 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6939 = _T_6937 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6940 = _T_6936 | _T_6939; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6950 = _T_4613 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6951 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6953 = _T_6951 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6954 = _T_6950 | _T_6953; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6964 = _T_4617 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6965 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6967 = _T_6965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6968 = _T_6964 | _T_6967; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6978 = _T_4621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6979 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6981 = _T_6979 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6982 = _T_6978 | _T_6981; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_6992 = _T_4625 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_6993 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_6995 = _T_6993 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_6996 = _T_6992 | _T_6995; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7006 = _T_4629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7007 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7009 = _T_7007 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7010 = _T_7006 | _T_7009; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7020 = _T_4633 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7021 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7023 = _T_7021 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7024 = _T_7020 | _T_7023; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7034 = _T_4637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7035 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7037 = _T_7035 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7038 = _T_7034 | _T_7037; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7048 = _T_4641 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7049 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7051 = _T_7049 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7052 = _T_7048 | _T_7051; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7062 = _T_4645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7063 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7065 = _T_7063 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7066 = _T_7062 | _T_7065; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7076 = _T_4649 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7077 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7079 = _T_7077 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7080 = _T_7076 | _T_7079; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7090 = _T_4653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7091 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7093 = _T_7091 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7094 = _T_7090 | _T_7093; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7104 = _T_4657 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7105 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7107 = _T_7105 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7108 = _T_7104 | _T_7107; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7118 = _T_4661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7119 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7121 = _T_7119 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7122 = _T_7118 | _T_7121; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7132 = _T_4665 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7133 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7135 = _T_7133 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7136 = _T_7132 | _T_7135; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7146 = _T_4669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7147 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7149 = _T_7147 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7150 = _T_7146 | _T_7149; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7160 = _T_4673 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7161 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7163 = _T_7161 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7164 = _T_7160 | _T_7163; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7174 = _T_4677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7175 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7177 = _T_7175 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7178 = _T_7174 | _T_7177; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7188 = _T_4681 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7189 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7191 = _T_7189 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7192 = _T_7188 | _T_7191; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7202 = _T_4685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7203 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7205 = _T_7203 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7206 = _T_7202 | _T_7205; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7216 = _T_4689 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7217 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7219 = _T_7217 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7220 = _T_7216 | _T_7219; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7230 = _T_4693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7231 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7233 = _T_7231 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7234 = _T_7230 | _T_7233; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7244 = _T_4697 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7245 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7247 = _T_7245 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7248 = _T_7244 | _T_7247; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7258 = _T_4701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7259 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7261 = _T_7259 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7262 = _T_7258 | _T_7261; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7272 = _T_4705 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7273 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7275 = _T_7273 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7276 = _T_7272 | _T_7275; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7286 = _T_4709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7287 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7289 = _T_7287 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7290 = _T_7286 | _T_7289; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7300 = _T_4713 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7301 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7303 = _T_7301 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7304 = _T_7300 | _T_7303; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7314 = _T_4589 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7317 = _T_6867 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7318 = _T_7314 | _T_7317; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7328 = _T_4593 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7331 = _T_6881 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7332 = _T_7328 | _T_7331; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7342 = _T_4597 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7345 = _T_6895 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7346 = _T_7342 | _T_7345; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7356 = _T_4601 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7359 = _T_6909 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7360 = _T_7356 | _T_7359; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7370 = _T_4605 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7373 = _T_6923 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7374 = _T_7370 | _T_7373; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7384 = _T_4609 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7387 = _T_6937 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7388 = _T_7384 | _T_7387; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7398 = _T_4613 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7401 = _T_6951 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7402 = _T_7398 | _T_7401; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7412 = _T_4617 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7415 = _T_6965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7416 = _T_7412 | _T_7415; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7426 = _T_4621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7429 = _T_6979 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7430 = _T_7426 | _T_7429; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7440 = _T_4625 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7443 = _T_6993 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7444 = _T_7440 | _T_7443; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7454 = _T_4629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7457 = _T_7007 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7458 = _T_7454 | _T_7457; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7468 = _T_4633 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7471 = _T_7021 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7472 = _T_7468 | _T_7471; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7482 = _T_4637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7485 = _T_7035 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7486 = _T_7482 | _T_7485; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7496 = _T_4641 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7499 = _T_7049 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7500 = _T_7496 | _T_7499; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7510 = _T_4645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7513 = _T_7063 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7514 = _T_7510 | _T_7513; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7524 = _T_4649 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7527 = _T_7077 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7528 = _T_7524 | _T_7527; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7538 = _T_4653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7541 = _T_7091 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7542 = _T_7538 | _T_7541; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7552 = _T_4657 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7555 = _T_7105 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7556 = _T_7552 | _T_7555; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7566 = _T_4661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7569 = _T_7119 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7570 = _T_7566 | _T_7569; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7580 = _T_4665 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7583 = _T_7133 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7584 = _T_7580 | _T_7583; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7594 = _T_4669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7597 = _T_7147 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7598 = _T_7594 | _T_7597; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7608 = _T_4673 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7611 = _T_7161 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7612 = _T_7608 | _T_7611; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7622 = _T_4677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7625 = _T_7175 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7626 = _T_7622 | _T_7625; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7636 = _T_4681 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7639 = _T_7189 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7640 = _T_7636 | _T_7639; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7650 = _T_4685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7653 = _T_7203 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7654 = _T_7650 | _T_7653; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7664 = _T_4689 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7667 = _T_7217 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7668 = _T_7664 | _T_7667; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7678 = _T_4693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7681 = _T_7231 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7682 = _T_7678 | _T_7681; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7692 = _T_4697 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7695 = _T_7245 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7696 = _T_7692 | _T_7695; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7706 = _T_4701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7709 = _T_7259 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7710 = _T_7706 | _T_7709; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7720 = _T_4705 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7723 = _T_7273 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7724 = _T_7720 | _T_7723; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7734 = _T_4709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7737 = _T_7287 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7738 = _T_7734 | _T_7737; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7748 = _T_4713 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7751 = _T_7301 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7752 = _T_7748 | _T_7751; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7762 = _T_4717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7763 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7765 = _T_7763 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7766 = _T_7762 | _T_7765; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7776 = _T_4721 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7777 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7779 = _T_7777 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7780 = _T_7776 | _T_7779; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7790 = _T_4725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7791 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7793 = _T_7791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7794 = _T_7790 | _T_7793; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7804 = _T_4729 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7805 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7807 = _T_7805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7808 = _T_7804 | _T_7807; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7818 = _T_4733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7819 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7821 = _T_7819 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7822 = _T_7818 | _T_7821; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7832 = _T_4737 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7833 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7835 = _T_7833 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7836 = _T_7832 | _T_7835; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7846 = _T_4741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7847 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7849 = _T_7847 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7850 = _T_7846 | _T_7849; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7860 = _T_4745 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7861 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7863 = _T_7861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7864 = _T_7860 | _T_7863; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7874 = _T_4749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7875 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7877 = _T_7875 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7878 = _T_7874 | _T_7877; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7888 = _T_4753 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7889 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7891 = _T_7889 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7892 = _T_7888 | _T_7891; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7902 = _T_4757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7903 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7905 = _T_7903 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7906 = _T_7902 | _T_7905; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7916 = _T_4761 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7917 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7919 = _T_7917 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7920 = _T_7916 | _T_7919; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7930 = _T_4765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7931 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7933 = _T_7931 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7934 = _T_7930 | _T_7933; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7944 = _T_4769 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7945 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7947 = _T_7945 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7948 = _T_7944 | _T_7947; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7958 = _T_4773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7959 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7961 = _T_7959 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7962 = _T_7958 | _T_7961; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7972 = _T_4777 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7973 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7975 = _T_7973 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7976 = _T_7972 | _T_7975; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_7986 = _T_4781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_7987 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_7989 = _T_7987 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_7990 = _T_7986 | _T_7989; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8000 = _T_4785 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8001 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8003 = _T_8001 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8004 = _T_8000 | _T_8003; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8014 = _T_4789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8015 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8017 = _T_8015 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8018 = _T_8014 | _T_8017; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8028 = _T_4793 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8029 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8031 = _T_8029 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8032 = _T_8028 | _T_8031; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8042 = _T_4797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8043 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8045 = _T_8043 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8046 = _T_8042 | _T_8045; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8056 = _T_4801 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8057 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8059 = _T_8057 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8060 = _T_8056 | _T_8059; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8070 = _T_4805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8071 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8073 = _T_8071 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8074 = _T_8070 | _T_8073; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8084 = _T_4809 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8085 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8087 = _T_8085 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8088 = _T_8084 | _T_8087; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8098 = _T_4813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8099 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8101 = _T_8099 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8102 = _T_8098 | _T_8101; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8112 = _T_4817 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8113 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8115 = _T_8113 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8116 = _T_8112 | _T_8115; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8126 = _T_4821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8127 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8129 = _T_8127 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8130 = _T_8126 | _T_8129; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8140 = _T_4825 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8141 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8143 = _T_8141 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8144 = _T_8140 | _T_8143; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8154 = _T_4829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8155 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8157 = _T_8155 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8158 = _T_8154 | _T_8157; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8168 = _T_4833 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8169 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8171 = _T_8169 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8172 = _T_8168 | _T_8171; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8182 = _T_4837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8183 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8185 = _T_8183 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8186 = _T_8182 | _T_8185; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8196 = _T_4841 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8197 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 792:101]
  wire  _T_8199 = _T_8197 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8200 = _T_8196 | _T_8199; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8210 = _T_4717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8213 = _T_7763 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8214 = _T_8210 | _T_8213; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8224 = _T_4721 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8227 = _T_7777 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8228 = _T_8224 | _T_8227; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8238 = _T_4725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8241 = _T_7791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8242 = _T_8238 | _T_8241; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8252 = _T_4729 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8255 = _T_7805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8256 = _T_8252 | _T_8255; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8266 = _T_4733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8269 = _T_7819 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8270 = _T_8266 | _T_8269; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8280 = _T_4737 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8283 = _T_7833 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8284 = _T_8280 | _T_8283; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8294 = _T_4741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8297 = _T_7847 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8298 = _T_8294 | _T_8297; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8308 = _T_4745 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8311 = _T_7861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8312 = _T_8308 | _T_8311; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8322 = _T_4749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8325 = _T_7875 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8326 = _T_8322 | _T_8325; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8336 = _T_4753 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8339 = _T_7889 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8340 = _T_8336 | _T_8339; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8350 = _T_4757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8353 = _T_7903 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8354 = _T_8350 | _T_8353; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8364 = _T_4761 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8367 = _T_7917 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8368 = _T_8364 | _T_8367; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8378 = _T_4765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8381 = _T_7931 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8382 = _T_8378 | _T_8381; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8392 = _T_4769 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8395 = _T_7945 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8396 = _T_8392 | _T_8395; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8406 = _T_4773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8409 = _T_7959 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8410 = _T_8406 | _T_8409; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8420 = _T_4777 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8423 = _T_7973 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8424 = _T_8420 | _T_8423; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8434 = _T_4781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8437 = _T_7987 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8438 = _T_8434 | _T_8437; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8448 = _T_4785 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8451 = _T_8001 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8452 = _T_8448 | _T_8451; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8462 = _T_4789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8465 = _T_8015 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8466 = _T_8462 | _T_8465; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8476 = _T_4793 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8479 = _T_8029 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8480 = _T_8476 | _T_8479; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8490 = _T_4797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8493 = _T_8043 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8494 = _T_8490 | _T_8493; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8504 = _T_4801 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8507 = _T_8057 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8508 = _T_8504 | _T_8507; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8518 = _T_4805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8521 = _T_8071 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8522 = _T_8518 | _T_8521; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8532 = _T_4809 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8535 = _T_8085 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8536 = _T_8532 | _T_8535; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8546 = _T_4813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8549 = _T_8099 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8550 = _T_8546 | _T_8549; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8560 = _T_4817 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8563 = _T_8113 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8564 = _T_8560 | _T_8563; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8574 = _T_4821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8577 = _T_8127 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8578 = _T_8574 | _T_8577; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8588 = _T_4825 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8591 = _T_8141 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8592 = _T_8588 | _T_8591; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8602 = _T_4829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8605 = _T_8155 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8606 = _T_8602 | _T_8605; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8616 = _T_4833 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8619 = _T_8169 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8620 = _T_8616 | _T_8619; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8630 = _T_4837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8633 = _T_8183 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8634 = _T_8630 | _T_8633; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_8644 = _T_4841 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  _T_8647 = _T_8197 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 792:123]
  wire  _T_8648 = _T_8644 | _T_8647; // @[el2_ifu_mem_ctl.scala 792:80]
  wire  _T_9449 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 847:63]
  wire  _T_9450 = _T_9449 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 847:85]
  wire [1:0] _T_9452 = _T_9450 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9459; // @[el2_ifu_mem_ctl.scala 852:58]
  reg  _T_9460; // @[el2_ifu_mem_ctl.scala 853:58]
  reg  _T_9461; // @[el2_ifu_mem_ctl.scala 854:59]
  wire  _T_9462 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 855:78]
  wire  _T_9463 = ifu_bus_arvalid_ff & _T_9462; // @[el2_ifu_mem_ctl.scala 855:76]
  wire  _T_9464 = _T_9463 & miss_pending; // @[el2_ifu_mem_ctl.scala 855:98]
  reg  _T_9465; // @[el2_ifu_mem_ctl.scala 855:56]
  reg  _T_9466; // @[el2_ifu_mem_ctl.scala 856:57]
  wire  _T_9469 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 861:71]
  wire  _T_9471 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 861:124]
  wire  _T_9473 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 862:50]
  wire  _T_9475 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 862:103]
  wire [3:0] _T_9478 = {_T_9469,_T_9471,_T_9473,_T_9475}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 864:53]
  reg  _T_9489; // @[Reg.scala 27:20]
  rvclkhdr rvclkhdr ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  rvclkhdr rvclkhdr_4 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_4_io_l1clk),
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en),
    .io_scan_mode(rvclkhdr_4_io_scan_mode)
  );
  rvclkhdr rvclkhdr_5 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_5_io_l1clk),
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en),
    .io_scan_mode(rvclkhdr_5_io_scan_mode)
  );
  rvclkhdr rvclkhdr_6 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_6_io_l1clk),
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en),
    .io_scan_mode(rvclkhdr_6_io_scan_mode)
  );
  rvclkhdr rvclkhdr_7 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_7_io_l1clk),
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en),
    .io_scan_mode(rvclkhdr_7_io_scan_mode)
  );
  rvclkhdr rvclkhdr_8 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_8_io_l1clk),
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en),
    .io_scan_mode(rvclkhdr_8_io_scan_mode)
  );
  rvclkhdr rvclkhdr_9 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_9_io_l1clk),
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en),
    .io_scan_mode(rvclkhdr_9_io_scan_mode)
  );
  rvclkhdr rvclkhdr_10 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_10_io_l1clk),
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en),
    .io_scan_mode(rvclkhdr_10_io_scan_mode)
  );
  rvclkhdr rvclkhdr_11 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_11_io_l1clk),
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en),
    .io_scan_mode(rvclkhdr_11_io_scan_mode)
  );
  rvclkhdr rvclkhdr_12 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_12_io_l1clk),
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en),
    .io_scan_mode(rvclkhdr_12_io_scan_mode)
  );
  rvclkhdr rvclkhdr_13 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_13_io_l1clk),
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en),
    .io_scan_mode(rvclkhdr_13_io_scan_mode)
  );
  rvclkhdr rvclkhdr_14 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_14_io_l1clk),
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en),
    .io_scan_mode(rvclkhdr_14_io_scan_mode)
  );
  rvclkhdr rvclkhdr_15 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_15_io_l1clk),
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en),
    .io_scan_mode(rvclkhdr_15_io_scan_mode)
  );
  rvclkhdr rvclkhdr_16 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_16_io_l1clk),
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en),
    .io_scan_mode(rvclkhdr_16_io_scan_mode)
  );
  rvclkhdr rvclkhdr_17 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_17_io_l1clk),
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en),
    .io_scan_mode(rvclkhdr_17_io_scan_mode)
  );
  rvclkhdr rvclkhdr_18 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_18_io_l1clk),
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en),
    .io_scan_mode(rvclkhdr_18_io_scan_mode)
  );
  rvclkhdr rvclkhdr_19 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_19_io_l1clk),
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en),
    .io_scan_mode(rvclkhdr_19_io_scan_mode)
  );
  rvclkhdr rvclkhdr_20 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_20_io_l1clk),
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en),
    .io_scan_mode(rvclkhdr_20_io_scan_mode)
  );
  rvclkhdr rvclkhdr_21 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_21_io_l1clk),
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en),
    .io_scan_mode(rvclkhdr_21_io_scan_mode)
  );
  rvclkhdr rvclkhdr_22 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_22_io_l1clk),
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en),
    .io_scan_mode(rvclkhdr_22_io_scan_mode)
  );
  rvclkhdr rvclkhdr_23 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_23_io_l1clk),
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en),
    .io_scan_mode(rvclkhdr_23_io_scan_mode)
  );
  rvclkhdr rvclkhdr_24 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_24_io_l1clk),
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en),
    .io_scan_mode(rvclkhdr_24_io_scan_mode)
  );
  rvclkhdr rvclkhdr_25 ( // @[el2_lib.scala 417:22]
    .io_l1clk(rvclkhdr_25_io_l1clk),
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en),
    .io_scan_mode(rvclkhdr_25_io_scan_mode)
  );
  assign io_ifu_miss_state_idle = 1'h0; // @[el2_ifu_mem_ctl.scala 131:25]
  assign io_ifu_ic_mb_empty = 1'h0; // @[el2_ifu_mem_ctl.scala 132:21]
  assign io_ic_dma_active = _T_12 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 133:19 el2_ifu_mem_ctl.scala 241:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3916; // @[el2_ifu_mem_ctl.scala 134:20 el2_ifu_mem_ctl.scala 739:21]
  assign io_ifu_pmu_ic_miss = _T_9466; // @[el2_ifu_mem_ctl.scala 135:21 el2_ifu_mem_ctl.scala 856:22]
  assign io_ifu_pmu_ic_hit = _T_9465; // @[el2_ifu_mem_ctl.scala 136:20 el2_ifu_mem_ctl.scala 855:21]
  assign io_ifu_pmu_bus_error = _T_9461; // @[el2_ifu_mem_ctl.scala 137:23 el2_ifu_mem_ctl.scala 854:24]
  assign io_ifu_pmu_bus_busy = _T_9460; // @[el2_ifu_mem_ctl.scala 138:22 el2_ifu_mem_ctl.scala 853:23]
  assign io_ifu_pmu_bus_trxn = _T_9459; // @[el2_ifu_mem_ctl.scala 139:22 el2_ifu_mem_ctl.scala 852:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 141:18]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 142:20]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 201:22]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 143:19]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 145:21]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 146:20]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 149:19]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 150:20]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 151:19]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 152:19]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 153:19]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 154:20]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 155:21 el2_ifu_mem_ctl.scala 601:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2510; // @[el2_ifu_mem_ctl.scala 157:18 el2_ifu_mem_ctl.scala 602:19]
  assign io_ifu_axi_araddr = _T_2512 & _T_2514; // @[el2_ifu_mem_ctl.scala 158:20 el2_ifu_mem_ctl.scala 603:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 159:22 el2_ifu_mem_ctl.scala 606:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 160:19]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 161:20 el2_ifu_mem_ctl.scala 604:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 162:21 el2_ifu_mem_ctl.scala 607:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 163:20]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 164:21 el2_ifu_mem_ctl.scala 605:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 165:20]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 166:19]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 167:20 el2_ifu_mem_ctl.scala 608:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 168:24 el2_ifu_mem_ctl.scala 698:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 169:21 el2_ifu_mem_ctl.scala 696:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 170:20 el2_ifu_mem_ctl.scala 700:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 171:19 el2_ifu_mem_ctl.scala 691:20]
  assign io_iccm_ready = 1'h0; // @[el2_ifu_mem_ctl.scala 172:16]
  assign io_ic_rw_addr = 31'h0; // @[el2_ifu_mem_ctl.scala 173:16]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 174:14 el2_ifu_mem_ctl.scala 738:15]
  assign io_ic_rd_en = _T_3894 | _T_3899; // @[el2_ifu_mem_ctl.scala 175:14 el2_ifu_mem_ctl.scala 729:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 176:16 el2_ifu_mem_ctl.scala 391:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 176:16 el2_ifu_mem_ctl.scala 391:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 177:22 el2_ifu_mem_ctl.scala 392:23]
  assign io_ifu_ic_debug_rd_data = _T_1201; // @[el2_ifu_mem_ctl.scala 178:26 el2_ifu_mem_ctl.scala 400:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 156:19 el2_ifu_mem_ctl.scala 857:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 128:20 el2_ifu_mem_ctl.scala 859:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 129:20 el2_ifu_mem_ctl.scala 860:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 130:24 el2_ifu_mem_ctl.scala 858:25]
  assign io_ic_debug_way = _T_9478[1:0]; // @[el2_ifu_mem_ctl.scala 200:18 el2_ifu_mem_ctl.scala 861:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9452; // @[el2_ifu_mem_ctl.scala 179:18 el2_ifu_mem_ctl.scala 847:19]
  assign io_iccm_rw_addr = _T_3048[14:0]; // @[el2_ifu_mem_ctl.scala 180:18 el2_ifu_mem_ctl.scala 702:19]
  assign io_iccm_wren = _T_2617 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 181:15 el2_ifu_mem_ctl.scala 673:16]
  assign io_iccm_rden = _T_2621 | _T_2622; // @[el2_ifu_mem_ctl.scala 182:15 el2_ifu_mem_ctl.scala 674:16]
  assign io_iccm_wr_data = _T_3023 ? _T_3024 : _T_3031; // @[el2_ifu_mem_ctl.scala 183:18 el2_ifu_mem_ctl.scala 679:19]
  assign io_iccm_wr_size = _T_2627 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 184:18 el2_ifu_mem_ctl.scala 676:19]
  assign io_ic_hit_f = _T_255 | _T_256; // @[el2_ifu_mem_ctl.scala 185:14 el2_ifu_mem_ctl.scala 336:15]
  assign io_ic_access_fault_f = _T_2400 & _T_309; // @[el2_ifu_mem_ctl.scala 186:23 el2_ifu_mem_ctl.scala 430:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1265; // @[el2_ifu_mem_ctl.scala 187:28 el2_ifu_mem_ctl.scala 431:29]
  assign io_iccm_rd_ecc_single_err = _T_3839 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 188:28 el2_ifu_mem_ctl.scala 715:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 189:28 el2_ifu_mem_ctl.scala 716:29]
  assign io_ic_error_start = _T_1189 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 190:20 el2_ifu_mem_ctl.scala 394:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:27 el2_ifu_mem_ctl.scala 240:28]
  assign io_iccm_dma_sb_error = _T_4 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 192:23 el2_ifu_mem_ctl.scala 239:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 193:20 el2_ifu_mem_ctl.scala 435:21]
  assign io_ic_data_f = 32'h0; // @[el2_ifu_mem_ctl.scala 194:15]
  assign io_ic_premux_data = 64'h0; // @[el2_ifu_mem_ctl.scala 195:20]
  assign io_ic_sel_premux_data = 1'h0; // @[el2_ifu_mem_ctl.scala 196:24]
  assign io_ifu_ic_debug_rd_data_valid = _T_9489; // @[el2_ifu_mem_ctl.scala 197:32 el2_ifu_mem_ctl.scala 868:33]
  assign io_iccm_buf_correct_ecc = 1'h0; // @[el2_ifu_mem_ctl.scala 198:26]
  assign io_iccm_correction_state = 1'h0; // @[el2_ifu_mem_ctl.scala 199:27]
  assign rvclkhdr_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_lib.scala 419:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_1_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_1_io_en = _T_1 | io_exu_flush_final; // @[el2_lib.scala 419:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_2_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_2_io_en = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_lib.scala 419:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_3_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_3_io_en = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_lib.scala 419:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_4_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_4_io_en = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_lib.scala 419:16]
  assign rvclkhdr_4_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_5_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_5_io_en = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_lib.scala 419:16]
  assign rvclkhdr_5_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_6_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_6_io_en = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_lib.scala 419:16]
  assign rvclkhdr_6_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_7_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_7_io_en = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_lib.scala 419:16]
  assign rvclkhdr_7_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_8_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_8_io_en = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_lib.scala 419:16]
  assign rvclkhdr_8_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_9_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_9_io_en = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_lib.scala 419:16]
  assign rvclkhdr_9_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_10_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_10_io_en = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_lib.scala 419:16]
  assign rvclkhdr_10_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_11_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_11_io_en = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_lib.scala 419:16]
  assign rvclkhdr_11_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_12_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_12_io_en = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_lib.scala 419:16]
  assign rvclkhdr_12_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_13_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_13_io_en = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_lib.scala 419:16]
  assign rvclkhdr_13_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_14_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_14_io_en = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_lib.scala 419:16]
  assign rvclkhdr_14_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_15_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_15_io_en = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_lib.scala 419:16]
  assign rvclkhdr_15_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_16_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_16_io_en = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_lib.scala 419:16]
  assign rvclkhdr_16_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_17_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_17_io_en = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_lib.scala 419:16]
  assign rvclkhdr_17_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_18_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_18_io_en = tag_valid_clken_0[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_18_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_19_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_19_io_en = tag_valid_clken_0[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_19_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_20_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_20_io_en = tag_valid_clken_1[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_20_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_21_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_21_io_en = tag_valid_clken_1[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_21_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_22_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_22_io_en = tag_valid_clken_2[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_22_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_23_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_23_io_en = tag_valid_clken_2[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_23_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_24_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_24_io_en = tag_valid_clken_3[0]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_24_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
  assign rvclkhdr_25_io_clk = clock; // @[el2_lib.scala 418:17]
  assign rvclkhdr_25_io_en = tag_valid_clken_3[1]; // @[el2_lib.scala 419:16]
  assign rvclkhdr_25_io_scan_mode = io_scan_mode; // @[el2_lib.scala 420:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  perr_state = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  err_stop_state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reset_all_tags = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  imb_ff = _RAND_16[30:0];
  _RAND_17 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_4976 = _RAND_19[6:0];
  _RAND_20 = {1{`RANDOM}};
  _T_4332 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4329 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4326 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4323 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4320 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4317 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4314 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4311 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4308 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4305 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4302 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4299 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4296 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4293 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4290 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4287 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4284 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4281 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4278 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4275 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4272 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4269 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4266 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4263 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4260 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4257 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4254 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4251 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4248 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4245 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4242 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4239 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4236 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4233 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4230 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4227 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4224 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4221 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4218 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4215 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4212 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4209 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4206 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4203 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4200 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4197 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4194 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4191 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4188 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4185 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_4182 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_4179 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_4176 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_4173 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_4170 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_4167 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_4164 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_4161 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_4158 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_4155 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4152 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4149 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4146 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4143 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_4140 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_4137 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_4134 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_4131 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4128 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4125 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4122 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4119 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4116 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4113 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4110 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4107 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_4104 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4101 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_4098 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_4095 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_4092 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_4089 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_4086 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_4083 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_4080 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_4077 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_4074 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_4071 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_4068 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_4065 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_4062 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_4059 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_4056 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_4053 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_4050 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_4047 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_4044 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_4041 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_4038 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_4035 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_4032 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_4029 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_4026 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_4023 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_4020 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_4017 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_4014 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_4011 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_4008 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4005 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4002 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_3999 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_3996 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_3993 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_3990 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3987 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3984 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3981 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3978 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3975 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3972 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3969 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3966 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3963 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3960 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3957 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3954 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3951 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_148[30:0];
  _RAND_149 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  reset_ic_ff = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  miss_addr = _RAND_155[25:0];
  _RAND_156 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_157[2:0];
  _RAND_158 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_158[0:0];
  _RAND_159 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  _T_1285 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  _T_1287 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  _T_1289 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  _T_1291 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  _T_1293 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  _T_1295 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  _T_1297 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  _T_1299 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  _T_1301 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  _T_1303 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  _T_1305 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  _T_1307 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  _T_1309 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  _T_1311 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  _T_1313 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  _T_1315 = _RAND_175[63:0];
  _RAND_176 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_436[0:0];
  _RAND_437 = {3{`RANDOM}};
  _T_1201 = _RAND_437[70:0];
  _RAND_438 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_438[5:0];
  _RAND_439 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_440[2:0];
  _RAND_441 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_441[0:0];
  _RAND_442 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_443[0:0];
  _RAND_444 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_444[38:0];
  _RAND_445 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_445[1:0];
  _RAND_446 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_446[2:0];
  _RAND_447 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_447[2:0];
  _RAND_448 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_449[63:0];
  _RAND_450 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_450[13:0];
  _RAND_451 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_451[0:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_452[13:0];
  _RAND_453 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_453[6:0];
  _RAND_454 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_454[0:0];
  _RAND_455 = {1{`RANDOM}};
  way_status_new_ff = _RAND_455[2:0];
  _RAND_456 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_456[1:0];
  _RAND_457 = {1{`RANDOM}};
  ic_valid_ff = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  _T_9459 = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  _T_9460 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  _T_9461 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  _T_9465 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  _T_9466 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_9489 = _RAND_463[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_26) begin
        if (_T_28) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_33) begin
        if (_T_38) begin
          miss_state <= 3'h0;
        end else if (_T_42) begin
          miss_state <= 3'h3;
        end else if (_T_49) begin
          miss_state <= 3'h1;
        end else if (_T_53) begin
          miss_state <= 3'h0;
        end else if (_T_64) begin
          miss_state <= 3'h6;
        end else if (_T_72) begin
          miss_state <= 3'h0;
        end else if (_T_77) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_94) begin
        miss_state <= 3'h0;
      end else if (_T_98) begin
        if (_T_105) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_113) begin
        if (_T_118) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_124) begin
        if (_T_129) begin
          miss_state <= 3'h5;
        end else if (_T_135) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_143) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_34) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_152) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_34) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    reset_ic_ff <= _T_290 & _T_291;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_223) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2553) begin
      if (_T_223) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2549;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1285 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1285 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1287 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1287 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1289 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1289 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1291 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1291 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1293 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1293 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1295 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1295 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1297 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1297 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1299 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1299 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1301 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1301 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1303 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1303 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1305 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1305 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1307 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1307 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1309 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1309 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1311 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1311 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1313 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1313 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1315 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1315 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1201 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1201 <= {{5'd0}, _T_1200};
    end else begin
      _T_1201 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2502) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2577) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2621;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2405) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2407) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2417) begin
        perr_state <= 3'h0;
      end else if (_T_2420) begin
        if (_T_2422) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2426) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2430) begin
        err_stop_state <= 2'h1;
      end else if (_T_2435) begin
        if (_T_2437) begin
          err_stop_state <= 2'h0;
        end else if (_T_2458) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2462) begin
        if (_T_2437) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2479) begin
        if (_T_2483) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1346;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_4976 <= 7'h0;
    end else if (_T_3925) begin
      _T_4976 <= io_ic_debug_addr[9:3];
    end else begin
      _T_4976 <= ic_rw_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1386;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3860;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3035;
    end else begin
      iccm_dma_rdata <= _T_3036;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3856;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3925) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3928) begin
      way_status_new_ff <= _T_3932;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3928) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_9489 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9489 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      _T_9459 <= 1'h0;
    end else begin
      _T_9459 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_9460 <= 1'h0;
    end else begin
      _T_9460 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_9461 <= 1'h0;
    end else begin
      _T_9461 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_9465 <= 1'h0;
    end else begin
      _T_9465 <= _T_9464;
    end
    if (reset) begin
      _T_9466 <= 1'h0;
    end else begin
      _T_9466 <= bus_cmd_sent;
    end
  end
  always @(posedge rvclkhdr_17_io_l1clk) begin
    if (reset) begin
      _T_4332 <= 3'h0;
    end else if (_T_3971) begin
      _T_4332 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4329 <= 3'h0;
    end else if (_T_3968) begin
      _T_4329 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4326 <= 3'h0;
    end else if (_T_3965) begin
      _T_4326 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4323 <= 3'h0;
    end else if (_T_3962) begin
      _T_4323 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4320 <= 3'h0;
    end else if (_T_3959) begin
      _T_4320 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4317 <= 3'h0;
    end else if (_T_3956) begin
      _T_4317 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4314 <= 3'h0;
    end else if (_T_3953) begin
      _T_4314 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4311 <= 3'h0;
    end else if (_T_3950) begin
      _T_4311 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_16_io_l1clk) begin
    if (reset) begin
      _T_4308 <= 3'h0;
    end else if (_T_3971) begin
      _T_4308 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4305 <= 3'h0;
    end else if (_T_3968) begin
      _T_4305 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4302 <= 3'h0;
    end else if (_T_3965) begin
      _T_4302 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4299 <= 3'h0;
    end else if (_T_3962) begin
      _T_4299 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4296 <= 3'h0;
    end else if (_T_3959) begin
      _T_4296 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4293 <= 3'h0;
    end else if (_T_3956) begin
      _T_4293 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4290 <= 3'h0;
    end else if (_T_3953) begin
      _T_4290 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4287 <= 3'h0;
    end else if (_T_3950) begin
      _T_4287 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_15_io_l1clk) begin
    if (reset) begin
      _T_4284 <= 3'h0;
    end else if (_T_3971) begin
      _T_4284 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4281 <= 3'h0;
    end else if (_T_3968) begin
      _T_4281 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4278 <= 3'h0;
    end else if (_T_3965) begin
      _T_4278 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4275 <= 3'h0;
    end else if (_T_3962) begin
      _T_4275 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4272 <= 3'h0;
    end else if (_T_3959) begin
      _T_4272 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4269 <= 3'h0;
    end else if (_T_3956) begin
      _T_4269 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4266 <= 3'h0;
    end else if (_T_3953) begin
      _T_4266 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4263 <= 3'h0;
    end else if (_T_3950) begin
      _T_4263 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_14_io_l1clk) begin
    if (reset) begin
      _T_4260 <= 3'h0;
    end else if (_T_3971) begin
      _T_4260 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4257 <= 3'h0;
    end else if (_T_3968) begin
      _T_4257 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4254 <= 3'h0;
    end else if (_T_3965) begin
      _T_4254 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4251 <= 3'h0;
    end else if (_T_3962) begin
      _T_4251 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4248 <= 3'h0;
    end else if (_T_3959) begin
      _T_4248 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4245 <= 3'h0;
    end else if (_T_3956) begin
      _T_4245 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4242 <= 3'h0;
    end else if (_T_3953) begin
      _T_4242 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4239 <= 3'h0;
    end else if (_T_3950) begin
      _T_4239 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_13_io_l1clk) begin
    if (reset) begin
      _T_4236 <= 3'h0;
    end else if (_T_3971) begin
      _T_4236 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4233 <= 3'h0;
    end else if (_T_3968) begin
      _T_4233 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4230 <= 3'h0;
    end else if (_T_3965) begin
      _T_4230 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4227 <= 3'h0;
    end else if (_T_3962) begin
      _T_4227 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4224 <= 3'h0;
    end else if (_T_3959) begin
      _T_4224 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4221 <= 3'h0;
    end else if (_T_3956) begin
      _T_4221 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4218 <= 3'h0;
    end else if (_T_3953) begin
      _T_4218 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4215 <= 3'h0;
    end else if (_T_3950) begin
      _T_4215 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_12_io_l1clk) begin
    if (reset) begin
      _T_4212 <= 3'h0;
    end else if (_T_3971) begin
      _T_4212 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4209 <= 3'h0;
    end else if (_T_3968) begin
      _T_4209 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4206 <= 3'h0;
    end else if (_T_3965) begin
      _T_4206 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4203 <= 3'h0;
    end else if (_T_3962) begin
      _T_4203 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4200 <= 3'h0;
    end else if (_T_3959) begin
      _T_4200 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4197 <= 3'h0;
    end else if (_T_3956) begin
      _T_4197 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4194 <= 3'h0;
    end else if (_T_3953) begin
      _T_4194 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4191 <= 3'h0;
    end else if (_T_3950) begin
      _T_4191 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_11_io_l1clk) begin
    if (reset) begin
      _T_4188 <= 3'h0;
    end else if (_T_3971) begin
      _T_4188 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4185 <= 3'h0;
    end else if (_T_3968) begin
      _T_4185 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4182 <= 3'h0;
    end else if (_T_3965) begin
      _T_4182 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4179 <= 3'h0;
    end else if (_T_3962) begin
      _T_4179 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4176 <= 3'h0;
    end else if (_T_3959) begin
      _T_4176 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4173 <= 3'h0;
    end else if (_T_3956) begin
      _T_4173 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4170 <= 3'h0;
    end else if (_T_3953) begin
      _T_4170 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4167 <= 3'h0;
    end else if (_T_3950) begin
      _T_4167 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_10_io_l1clk) begin
    if (reset) begin
      _T_4164 <= 3'h0;
    end else if (_T_3971) begin
      _T_4164 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4161 <= 3'h0;
    end else if (_T_3968) begin
      _T_4161 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4158 <= 3'h0;
    end else if (_T_3965) begin
      _T_4158 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4155 <= 3'h0;
    end else if (_T_3962) begin
      _T_4155 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4152 <= 3'h0;
    end else if (_T_3959) begin
      _T_4152 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4149 <= 3'h0;
    end else if (_T_3956) begin
      _T_4149 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4146 <= 3'h0;
    end else if (_T_3953) begin
      _T_4146 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4143 <= 3'h0;
    end else if (_T_3950) begin
      _T_4143 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_9_io_l1clk) begin
    if (reset) begin
      _T_4140 <= 3'h0;
    end else if (_T_3971) begin
      _T_4140 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4137 <= 3'h0;
    end else if (_T_3968) begin
      _T_4137 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4134 <= 3'h0;
    end else if (_T_3965) begin
      _T_4134 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4131 <= 3'h0;
    end else if (_T_3962) begin
      _T_4131 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4128 <= 3'h0;
    end else if (_T_3959) begin
      _T_4128 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4125 <= 3'h0;
    end else if (_T_3956) begin
      _T_4125 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4122 <= 3'h0;
    end else if (_T_3953) begin
      _T_4122 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4119 <= 3'h0;
    end else if (_T_3950) begin
      _T_4119 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_8_io_l1clk) begin
    if (reset) begin
      _T_4116 <= 3'h0;
    end else if (_T_3971) begin
      _T_4116 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4113 <= 3'h0;
    end else if (_T_3968) begin
      _T_4113 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4110 <= 3'h0;
    end else if (_T_3965) begin
      _T_4110 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4107 <= 3'h0;
    end else if (_T_3962) begin
      _T_4107 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4104 <= 3'h0;
    end else if (_T_3959) begin
      _T_4104 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4101 <= 3'h0;
    end else if (_T_3956) begin
      _T_4101 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4098 <= 3'h0;
    end else if (_T_3953) begin
      _T_4098 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4095 <= 3'h0;
    end else if (_T_3950) begin
      _T_4095 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_7_io_l1clk) begin
    if (reset) begin
      _T_4092 <= 3'h0;
    end else if (_T_3971) begin
      _T_4092 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4089 <= 3'h0;
    end else if (_T_3968) begin
      _T_4089 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4086 <= 3'h0;
    end else if (_T_3965) begin
      _T_4086 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4083 <= 3'h0;
    end else if (_T_3962) begin
      _T_4083 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4080 <= 3'h0;
    end else if (_T_3959) begin
      _T_4080 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4077 <= 3'h0;
    end else if (_T_3956) begin
      _T_4077 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4074 <= 3'h0;
    end else if (_T_3953) begin
      _T_4074 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4071 <= 3'h0;
    end else if (_T_3950) begin
      _T_4071 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_6_io_l1clk) begin
    if (reset) begin
      _T_4068 <= 3'h0;
    end else if (_T_3971) begin
      _T_4068 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4065 <= 3'h0;
    end else if (_T_3968) begin
      _T_4065 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4062 <= 3'h0;
    end else if (_T_3965) begin
      _T_4062 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4059 <= 3'h0;
    end else if (_T_3962) begin
      _T_4059 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4056 <= 3'h0;
    end else if (_T_3959) begin
      _T_4056 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4053 <= 3'h0;
    end else if (_T_3956) begin
      _T_4053 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4050 <= 3'h0;
    end else if (_T_3953) begin
      _T_4050 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4047 <= 3'h0;
    end else if (_T_3950) begin
      _T_4047 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_5_io_l1clk) begin
    if (reset) begin
      _T_4044 <= 3'h0;
    end else if (_T_3971) begin
      _T_4044 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4041 <= 3'h0;
    end else if (_T_3968) begin
      _T_4041 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4038 <= 3'h0;
    end else if (_T_3965) begin
      _T_4038 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4035 <= 3'h0;
    end else if (_T_3962) begin
      _T_4035 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4032 <= 3'h0;
    end else if (_T_3959) begin
      _T_4032 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4029 <= 3'h0;
    end else if (_T_3956) begin
      _T_4029 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4026 <= 3'h0;
    end else if (_T_3953) begin
      _T_4026 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4023 <= 3'h0;
    end else if (_T_3950) begin
      _T_4023 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_4_io_l1clk) begin
    if (reset) begin
      _T_4020 <= 3'h0;
    end else if (_T_3971) begin
      _T_4020 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4017 <= 3'h0;
    end else if (_T_3968) begin
      _T_4017 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4014 <= 3'h0;
    end else if (_T_3965) begin
      _T_4014 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4011 <= 3'h0;
    end else if (_T_3962) begin
      _T_4011 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4008 <= 3'h0;
    end else if (_T_3959) begin
      _T_4008 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4005 <= 3'h0;
    end else if (_T_3956) begin
      _T_4005 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4002 <= 3'h0;
    end else if (_T_3953) begin
      _T_4002 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3999 <= 3'h0;
    end else if (_T_3950) begin
      _T_3999 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk) begin
    if (reset) begin
      _T_3996 <= 3'h0;
    end else if (_T_3971) begin
      _T_3996 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3993 <= 3'h0;
    end else if (_T_3968) begin
      _T_3993 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3990 <= 3'h0;
    end else if (_T_3965) begin
      _T_3990 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3987 <= 3'h0;
    end else if (_T_3962) begin
      _T_3987 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3984 <= 3'h0;
    end else if (_T_3959) begin
      _T_3984 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3981 <= 3'h0;
    end else if (_T_3956) begin
      _T_3981 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3978 <= 3'h0;
    end else if (_T_3953) begin
      _T_3978 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3975 <= 3'h0;
    end else if (_T_3950) begin
      _T_3975 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk) begin
    if (reset) begin
      _T_3972 <= 3'h0;
    end else if (_T_3971) begin
      _T_3972 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3969 <= 3'h0;
    end else if (_T_3968) begin
      _T_3969 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3966 <= 3'h0;
    end else if (_T_3965) begin
      _T_3966 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3963 <= 3'h0;
    end else if (_T_3962) begin
      _T_3963 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3960 <= 3'h0;
    end else if (_T_3959) begin
      _T_3960 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3957 <= 3'h0;
    end else if (_T_3956) begin
      _T_3957 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3954 <= 3'h0;
    end else if (_T_3953) begin
      _T_3954 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3951 <= 3'h0;
    end else if (_T_3950) begin
      _T_3951 <= way_status_new_ff;
    end
  end
  always @(posedge rvclkhdr_19_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5526) begin
      ic_tag_valid_out_1_0 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5540) begin
      ic_tag_valid_out_1_1 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5554) begin
      ic_tag_valid_out_1_2 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5568) begin
      ic_tag_valid_out_1_3 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5582) begin
      ic_tag_valid_out_1_4 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5596) begin
      ic_tag_valid_out_1_5 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5610) begin
      ic_tag_valid_out_1_6 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5624) begin
      ic_tag_valid_out_1_7 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5638) begin
      ic_tag_valid_out_1_8 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5652) begin
      ic_tag_valid_out_1_9 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5666) begin
      ic_tag_valid_out_1_10 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5680) begin
      ic_tag_valid_out_1_11 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5694) begin
      ic_tag_valid_out_1_12 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5708) begin
      ic_tag_valid_out_1_13 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5722) begin
      ic_tag_valid_out_1_14 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5736) begin
      ic_tag_valid_out_1_15 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5750) begin
      ic_tag_valid_out_1_16 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5764) begin
      ic_tag_valid_out_1_17 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5778) begin
      ic_tag_valid_out_1_18 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5792) begin
      ic_tag_valid_out_1_19 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5806) begin
      ic_tag_valid_out_1_20 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5820) begin
      ic_tag_valid_out_1_21 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5834) begin
      ic_tag_valid_out_1_22 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5848) begin
      ic_tag_valid_out_1_23 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5862) begin
      ic_tag_valid_out_1_24 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5876) begin
      ic_tag_valid_out_1_25 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5890) begin
      ic_tag_valid_out_1_26 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5904) begin
      ic_tag_valid_out_1_27 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_5918) begin
      ic_tag_valid_out_1_28 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_5932) begin
      ic_tag_valid_out_1_29 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_5946) begin
      ic_tag_valid_out_1_30 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_5960) begin
      ic_tag_valid_out_1_31 <= _T_5071;
    end
  end
  always @(posedge rvclkhdr_21_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6422) begin
      ic_tag_valid_out_1_32 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6436) begin
      ic_tag_valid_out_1_33 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6450) begin
      ic_tag_valid_out_1_34 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6464) begin
      ic_tag_valid_out_1_35 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6478) begin
      ic_tag_valid_out_1_36 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6492) begin
      ic_tag_valid_out_1_37 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6506) begin
      ic_tag_valid_out_1_38 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6520) begin
      ic_tag_valid_out_1_39 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6534) begin
      ic_tag_valid_out_1_40 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6548) begin
      ic_tag_valid_out_1_41 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6562) begin
      ic_tag_valid_out_1_42 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6576) begin
      ic_tag_valid_out_1_43 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6590) begin
      ic_tag_valid_out_1_44 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6604) begin
      ic_tag_valid_out_1_45 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6618) begin
      ic_tag_valid_out_1_46 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6632) begin
      ic_tag_valid_out_1_47 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6646) begin
      ic_tag_valid_out_1_48 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6660) begin
      ic_tag_valid_out_1_49 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6674) begin
      ic_tag_valid_out_1_50 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6688) begin
      ic_tag_valid_out_1_51 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6702) begin
      ic_tag_valid_out_1_52 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6716) begin
      ic_tag_valid_out_1_53 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6730) begin
      ic_tag_valid_out_1_54 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6744) begin
      ic_tag_valid_out_1_55 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6758) begin
      ic_tag_valid_out_1_56 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6772) begin
      ic_tag_valid_out_1_57 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6786) begin
      ic_tag_valid_out_1_58 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6800) begin
      ic_tag_valid_out_1_59 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6814) begin
      ic_tag_valid_out_1_60 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6828) begin
      ic_tag_valid_out_1_61 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_6842) begin
      ic_tag_valid_out_1_62 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_6856) begin
      ic_tag_valid_out_1_63 <= _T_5071;
    end
  end
  always @(posedge rvclkhdr_23_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7318) begin
      ic_tag_valid_out_1_64 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7332) begin
      ic_tag_valid_out_1_65 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7346) begin
      ic_tag_valid_out_1_66 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7360) begin
      ic_tag_valid_out_1_67 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7374) begin
      ic_tag_valid_out_1_68 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7388) begin
      ic_tag_valid_out_1_69 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7402) begin
      ic_tag_valid_out_1_70 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7416) begin
      ic_tag_valid_out_1_71 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7430) begin
      ic_tag_valid_out_1_72 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7444) begin
      ic_tag_valid_out_1_73 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7458) begin
      ic_tag_valid_out_1_74 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7472) begin
      ic_tag_valid_out_1_75 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7486) begin
      ic_tag_valid_out_1_76 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7500) begin
      ic_tag_valid_out_1_77 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7514) begin
      ic_tag_valid_out_1_78 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7528) begin
      ic_tag_valid_out_1_79 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7542) begin
      ic_tag_valid_out_1_80 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7556) begin
      ic_tag_valid_out_1_81 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7570) begin
      ic_tag_valid_out_1_82 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7584) begin
      ic_tag_valid_out_1_83 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7598) begin
      ic_tag_valid_out_1_84 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7612) begin
      ic_tag_valid_out_1_85 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7626) begin
      ic_tag_valid_out_1_86 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7640) begin
      ic_tag_valid_out_1_87 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7654) begin
      ic_tag_valid_out_1_88 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7668) begin
      ic_tag_valid_out_1_89 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7682) begin
      ic_tag_valid_out_1_90 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7696) begin
      ic_tag_valid_out_1_91 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7710) begin
      ic_tag_valid_out_1_92 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7724) begin
      ic_tag_valid_out_1_93 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7738) begin
      ic_tag_valid_out_1_94 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7752) begin
      ic_tag_valid_out_1_95 <= _T_5071;
    end
  end
  always @(posedge rvclkhdr_25_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8214) begin
      ic_tag_valid_out_1_96 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8228) begin
      ic_tag_valid_out_1_97 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8242) begin
      ic_tag_valid_out_1_98 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8256) begin
      ic_tag_valid_out_1_99 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8270) begin
      ic_tag_valid_out_1_100 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8284) begin
      ic_tag_valid_out_1_101 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8298) begin
      ic_tag_valid_out_1_102 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8312) begin
      ic_tag_valid_out_1_103 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8326) begin
      ic_tag_valid_out_1_104 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8340) begin
      ic_tag_valid_out_1_105 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8354) begin
      ic_tag_valid_out_1_106 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8368) begin
      ic_tag_valid_out_1_107 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8382) begin
      ic_tag_valid_out_1_108 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8396) begin
      ic_tag_valid_out_1_109 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8410) begin
      ic_tag_valid_out_1_110 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8424) begin
      ic_tag_valid_out_1_111 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8438) begin
      ic_tag_valid_out_1_112 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8452) begin
      ic_tag_valid_out_1_113 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8466) begin
      ic_tag_valid_out_1_114 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8480) begin
      ic_tag_valid_out_1_115 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8494) begin
      ic_tag_valid_out_1_116 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8508) begin
      ic_tag_valid_out_1_117 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8522) begin
      ic_tag_valid_out_1_118 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8536) begin
      ic_tag_valid_out_1_119 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8550) begin
      ic_tag_valid_out_1_120 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8564) begin
      ic_tag_valid_out_1_121 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8578) begin
      ic_tag_valid_out_1_122 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8592) begin
      ic_tag_valid_out_1_123 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8606) begin
      ic_tag_valid_out_1_124 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8620) begin
      ic_tag_valid_out_1_125 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8634) begin
      ic_tag_valid_out_1_126 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8648) begin
      ic_tag_valid_out_1_127 <= _T_5071;
    end
  end
  always @(posedge rvclkhdr_18_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5078) begin
      ic_tag_valid_out_0_0 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5092) begin
      ic_tag_valid_out_0_1 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5106) begin
      ic_tag_valid_out_0_2 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5120) begin
      ic_tag_valid_out_0_3 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5134) begin
      ic_tag_valid_out_0_4 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5148) begin
      ic_tag_valid_out_0_5 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5162) begin
      ic_tag_valid_out_0_6 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5176) begin
      ic_tag_valid_out_0_7 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5190) begin
      ic_tag_valid_out_0_8 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5204) begin
      ic_tag_valid_out_0_9 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5218) begin
      ic_tag_valid_out_0_10 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5232) begin
      ic_tag_valid_out_0_11 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5246) begin
      ic_tag_valid_out_0_12 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5260) begin
      ic_tag_valid_out_0_13 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5274) begin
      ic_tag_valid_out_0_14 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5288) begin
      ic_tag_valid_out_0_15 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5302) begin
      ic_tag_valid_out_0_16 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5316) begin
      ic_tag_valid_out_0_17 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5330) begin
      ic_tag_valid_out_0_18 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5344) begin
      ic_tag_valid_out_0_19 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5358) begin
      ic_tag_valid_out_0_20 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5372) begin
      ic_tag_valid_out_0_21 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5386) begin
      ic_tag_valid_out_0_22 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5400) begin
      ic_tag_valid_out_0_23 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5414) begin
      ic_tag_valid_out_0_24 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5428) begin
      ic_tag_valid_out_0_25 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5442) begin
      ic_tag_valid_out_0_26 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5456) begin
      ic_tag_valid_out_0_27 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5470) begin
      ic_tag_valid_out_0_28 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5484) begin
      ic_tag_valid_out_0_29 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5498) begin
      ic_tag_valid_out_0_30 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5512) begin
      ic_tag_valid_out_0_31 <= _T_5071;
    end
  end
  always @(posedge rvclkhdr_20_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_5974) begin
      ic_tag_valid_out_0_32 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_5988) begin
      ic_tag_valid_out_0_33 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6002) begin
      ic_tag_valid_out_0_34 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6016) begin
      ic_tag_valid_out_0_35 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6030) begin
      ic_tag_valid_out_0_36 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6044) begin
      ic_tag_valid_out_0_37 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6058) begin
      ic_tag_valid_out_0_38 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6072) begin
      ic_tag_valid_out_0_39 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6086) begin
      ic_tag_valid_out_0_40 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6100) begin
      ic_tag_valid_out_0_41 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6114) begin
      ic_tag_valid_out_0_42 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6128) begin
      ic_tag_valid_out_0_43 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6142) begin
      ic_tag_valid_out_0_44 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6156) begin
      ic_tag_valid_out_0_45 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6170) begin
      ic_tag_valid_out_0_46 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6184) begin
      ic_tag_valid_out_0_47 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6198) begin
      ic_tag_valid_out_0_48 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6212) begin
      ic_tag_valid_out_0_49 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6226) begin
      ic_tag_valid_out_0_50 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6240) begin
      ic_tag_valid_out_0_51 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6254) begin
      ic_tag_valid_out_0_52 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6268) begin
      ic_tag_valid_out_0_53 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6282) begin
      ic_tag_valid_out_0_54 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6296) begin
      ic_tag_valid_out_0_55 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6310) begin
      ic_tag_valid_out_0_56 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6324) begin
      ic_tag_valid_out_0_57 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6338) begin
      ic_tag_valid_out_0_58 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6352) begin
      ic_tag_valid_out_0_59 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6366) begin
      ic_tag_valid_out_0_60 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6380) begin
      ic_tag_valid_out_0_61 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6394) begin
      ic_tag_valid_out_0_62 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6408) begin
      ic_tag_valid_out_0_63 <= _T_5071;
    end
  end
  always @(posedge rvclkhdr_22_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_6870) begin
      ic_tag_valid_out_0_64 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_6884) begin
      ic_tag_valid_out_0_65 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_6898) begin
      ic_tag_valid_out_0_66 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_6912) begin
      ic_tag_valid_out_0_67 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_6926) begin
      ic_tag_valid_out_0_68 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_6940) begin
      ic_tag_valid_out_0_69 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_6954) begin
      ic_tag_valid_out_0_70 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_6968) begin
      ic_tag_valid_out_0_71 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_6982) begin
      ic_tag_valid_out_0_72 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_6996) begin
      ic_tag_valid_out_0_73 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7010) begin
      ic_tag_valid_out_0_74 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7024) begin
      ic_tag_valid_out_0_75 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7038) begin
      ic_tag_valid_out_0_76 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7052) begin
      ic_tag_valid_out_0_77 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7066) begin
      ic_tag_valid_out_0_78 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7080) begin
      ic_tag_valid_out_0_79 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7094) begin
      ic_tag_valid_out_0_80 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7108) begin
      ic_tag_valid_out_0_81 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7122) begin
      ic_tag_valid_out_0_82 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7136) begin
      ic_tag_valid_out_0_83 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7150) begin
      ic_tag_valid_out_0_84 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7164) begin
      ic_tag_valid_out_0_85 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7178) begin
      ic_tag_valid_out_0_86 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7192) begin
      ic_tag_valid_out_0_87 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7206) begin
      ic_tag_valid_out_0_88 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7220) begin
      ic_tag_valid_out_0_89 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7234) begin
      ic_tag_valid_out_0_90 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7248) begin
      ic_tag_valid_out_0_91 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7262) begin
      ic_tag_valid_out_0_92 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7276) begin
      ic_tag_valid_out_0_93 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7290) begin
      ic_tag_valid_out_0_94 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7304) begin
      ic_tag_valid_out_0_95 <= _T_5071;
    end
  end
  always @(posedge rvclkhdr_24_io_l1clk) begin
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7766) begin
      ic_tag_valid_out_0_96 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_7780) begin
      ic_tag_valid_out_0_97 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_7794) begin
      ic_tag_valid_out_0_98 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_7808) begin
      ic_tag_valid_out_0_99 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_7822) begin
      ic_tag_valid_out_0_100 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_7836) begin
      ic_tag_valid_out_0_101 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_7850) begin
      ic_tag_valid_out_0_102 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_7864) begin
      ic_tag_valid_out_0_103 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_7878) begin
      ic_tag_valid_out_0_104 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_7892) begin
      ic_tag_valid_out_0_105 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_7906) begin
      ic_tag_valid_out_0_106 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_7920) begin
      ic_tag_valid_out_0_107 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_7934) begin
      ic_tag_valid_out_0_108 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_7948) begin
      ic_tag_valid_out_0_109 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_7962) begin
      ic_tag_valid_out_0_110 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_7976) begin
      ic_tag_valid_out_0_111 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_7990) begin
      ic_tag_valid_out_0_112 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8004) begin
      ic_tag_valid_out_0_113 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8018) begin
      ic_tag_valid_out_0_114 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8032) begin
      ic_tag_valid_out_0_115 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8046) begin
      ic_tag_valid_out_0_116 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8060) begin
      ic_tag_valid_out_0_117 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8074) begin
      ic_tag_valid_out_0_118 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8088) begin
      ic_tag_valid_out_0_119 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8102) begin
      ic_tag_valid_out_0_120 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8116) begin
      ic_tag_valid_out_0_121 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8130) begin
      ic_tag_valid_out_0_122 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8144) begin
      ic_tag_valid_out_0_123 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8158) begin
      ic_tag_valid_out_0_124 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8172) begin
      ic_tag_valid_out_0_125 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8186) begin
      ic_tag_valid_out_0_126 <= _T_5071;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8200) begin
      ic_tag_valid_out_0_127 <= _T_5071;
    end
  end
endmodule
