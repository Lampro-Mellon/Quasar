module el2_ifu_bp_ctl(
  input         clock,
  input         reset,
  input         io_active_clk,
  input         io_ic_hit_f,
  input  [30:0] io_ifc_fetch_addr_f,
  input         io_ifc_fetch_req_f,
  input         io_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_dec_tlu_br0_r_pkt_hist,
  input         io_dec_tlu_br0_r_pkt_br_error,
  input         io_dec_tlu_br0_r_pkt_br_start_error,
  input         io_dec_tlu_br0_r_pkt_way,
  input         io_dec_tlu_br0_r_pkt_middle,
  input  [7:0]  io_exu_i0_br_fghr_r,
  input  [7:0]  io_exu_i0_br_index_r,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_leak_one_wb,
  input         io_dec_tlu_bpred_disable,
  input         io_exu_mp_pkt_misp,
  input         io_exu_mp_pkt_ataken,
  input         io_exu_mp_pkt_boffset,
  input         io_exu_mp_pkt_pc4,
  input  [1:0]  io_exu_mp_pkt_hist,
  input  [11:0] io_exu_mp_pkt_toffset,
  input         io_exu_mp_pkt_valid,
  input         io_exu_mp_pkt_br_error,
  input         io_exu_mp_pkt_br_start_error,
  input  [31:0] io_exu_mp_pkt_prett,
  input         io_exu_mp_pkt_pcall,
  input         io_exu_mp_pkt_pret,
  input         io_exu_mp_pkt_pja,
  input         io_exu_mp_pkt_way,
  input  [7:0]  io_exu_mp_eghr,
  input  [7:0]  io_exu_mp_fghr,
  input  [7:0]  io_exu_mp_index,
  input  [4:0]  io_exu_mp_btag,
  input         io_exu_flush_final,
  output        io_ifu_bp_hit_taken_f,
  output [30:0] io_ifu_bp_btb_target_f,
  output        io_ifu_bp_inst_mask_f,
  output [7:0]  io_ifu_bp_fghr_f,
  output [1:0]  io_ifu_bp_way_f,
  output [1:0]  io_ifu_bp_ret_f,
  output [1:0]  io_ifu_bp_hist1_f,
  output [1:0]  io_ifu_bp_hist0_f,
  output [1:0]  io_ifu_bp_pc4_f,
  output [1:0]  io_ifu_bp_valid_f,
  output [11:0] io_ifu_bp_poffset_f,
  output [7:0]  io_test_hash,
  output [7:0]  io_test_hash_p1,
  output [1:0]  io_test
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [31:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [255:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
  reg [31:0] _RAND_1038;
`endif // RANDOMIZE_REG_INIT
  wire  _T_40 = io_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_bp_ctl.scala 133:47]
  reg  leak_one_f_d1; // @[el2_ifu_bp_ctl.scala 127:30]
  wire  _T_41 = leak_one_f_d1 & io_dec_tlu_flush_lower_wb; // @[el2_ifu_bp_ctl.scala 133:93]
  wire  leak_one_f = _T_40 | _T_41; // @[el2_ifu_bp_ctl.scala 133:76]
  wire  _T = ~leak_one_f; // @[el2_ifu_bp_ctl.scala 73:46]
  wire  exu_mp_valid = io_exu_mp_pkt_misp & _T; // @[el2_ifu_bp_ctl.scala 73:44]
  wire  dec_tlu_error_wb = io_dec_tlu_br0_r_pkt_br_start_error | io_dec_tlu_br0_r_pkt_br_error; // @[el2_ifu_bp_ctl.scala 95:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[el2_lib.scala 183:46]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[el2_lib.scala 183:84]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[el2_ifu_bp_ctl.scala 103:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[el2_lib.scala 183:46]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[el2_lib.scala 183:84]
  wire  _T_143 = ~io_ifc_fetch_addr_f[0]; // @[el2_ifu_bp_ctl.scala 179:40]
  wire  _T_2108 = btb_rd_addr_f == 8'h0; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_2620 = _T_2108 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2110 = btb_rd_addr_f == 8'h1; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_2621 = _T_2110 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2876 = _T_2620 | _T_2621; // @[Mux.scala 27:72]
  wire  _T_2112 = btb_rd_addr_f == 8'h2; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_2622 = _T_2112 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2877 = _T_2876 | _T_2622; // @[Mux.scala 27:72]
  wire  _T_2114 = btb_rd_addr_f == 8'h3; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_2623 = _T_2114 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2878 = _T_2877 | _T_2623; // @[Mux.scala 27:72]
  wire  _T_2116 = btb_rd_addr_f == 8'h4; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_2624 = _T_2116 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2879 = _T_2878 | _T_2624; // @[Mux.scala 27:72]
  wire  _T_2118 = btb_rd_addr_f == 8'h5; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_2625 = _T_2118 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2880 = _T_2879 | _T_2625; // @[Mux.scala 27:72]
  wire  _T_2120 = btb_rd_addr_f == 8'h6; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_2626 = _T_2120 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2881 = _T_2880 | _T_2626; // @[Mux.scala 27:72]
  wire  _T_2122 = btb_rd_addr_f == 8'h7; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_2627 = _T_2122 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2882 = _T_2881 | _T_2627; // @[Mux.scala 27:72]
  wire  _T_2124 = btb_rd_addr_f == 8'h8; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_2628 = _T_2124 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2883 = _T_2882 | _T_2628; // @[Mux.scala 27:72]
  wire  _T_2126 = btb_rd_addr_f == 8'h9; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_2629 = _T_2126 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2884 = _T_2883 | _T_2629; // @[Mux.scala 27:72]
  wire  _T_2128 = btb_rd_addr_f == 8'ha; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_2630 = _T_2128 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2885 = _T_2884 | _T_2630; // @[Mux.scala 27:72]
  wire  _T_2130 = btb_rd_addr_f == 8'hb; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_2631 = _T_2130 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2886 = _T_2885 | _T_2631; // @[Mux.scala 27:72]
  wire  _T_2132 = btb_rd_addr_f == 8'hc; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_2632 = _T_2132 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2887 = _T_2886 | _T_2632; // @[Mux.scala 27:72]
  wire  _T_2134 = btb_rd_addr_f == 8'hd; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_2633 = _T_2134 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2888 = _T_2887 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2136 = btb_rd_addr_f == 8'he; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_2634 = _T_2136 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2889 = _T_2888 | _T_2634; // @[Mux.scala 27:72]
  wire  _T_2138 = btb_rd_addr_f == 8'hf; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_2635 = _T_2138 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2890 = _T_2889 | _T_2635; // @[Mux.scala 27:72]
  wire  _T_2140 = btb_rd_addr_f == 8'h10; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_2636 = _T_2140 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2891 = _T_2890 | _T_2636; // @[Mux.scala 27:72]
  wire  _T_2142 = btb_rd_addr_f == 8'h11; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_2637 = _T_2142 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2892 = _T_2891 | _T_2637; // @[Mux.scala 27:72]
  wire  _T_2144 = btb_rd_addr_f == 8'h12; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_2638 = _T_2144 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2893 = _T_2892 | _T_2638; // @[Mux.scala 27:72]
  wire  _T_2146 = btb_rd_addr_f == 8'h13; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_2639 = _T_2146 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2894 = _T_2893 | _T_2639; // @[Mux.scala 27:72]
  wire  _T_2148 = btb_rd_addr_f == 8'h14; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_2640 = _T_2148 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2895 = _T_2894 | _T_2640; // @[Mux.scala 27:72]
  wire  _T_2150 = btb_rd_addr_f == 8'h15; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_2641 = _T_2150 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2896 = _T_2895 | _T_2641; // @[Mux.scala 27:72]
  wire  _T_2152 = btb_rd_addr_f == 8'h16; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_2642 = _T_2152 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2897 = _T_2896 | _T_2642; // @[Mux.scala 27:72]
  wire  _T_2154 = btb_rd_addr_f == 8'h17; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_2643 = _T_2154 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2898 = _T_2897 | _T_2643; // @[Mux.scala 27:72]
  wire  _T_2156 = btb_rd_addr_f == 8'h18; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_2644 = _T_2156 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2899 = _T_2898 | _T_2644; // @[Mux.scala 27:72]
  wire  _T_2158 = btb_rd_addr_f == 8'h19; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_2645 = _T_2158 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2900 = _T_2899 | _T_2645; // @[Mux.scala 27:72]
  wire  _T_2160 = btb_rd_addr_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_2646 = _T_2160 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2901 = _T_2900 | _T_2646; // @[Mux.scala 27:72]
  wire  _T_2162 = btb_rd_addr_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_2647 = _T_2162 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2902 = _T_2901 | _T_2647; // @[Mux.scala 27:72]
  wire  _T_2164 = btb_rd_addr_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_2648 = _T_2164 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2903 = _T_2902 | _T_2648; // @[Mux.scala 27:72]
  wire  _T_2166 = btb_rd_addr_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_2649 = _T_2166 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2904 = _T_2903 | _T_2649; // @[Mux.scala 27:72]
  wire  _T_2168 = btb_rd_addr_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_2650 = _T_2168 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2905 = _T_2904 | _T_2650; // @[Mux.scala 27:72]
  wire  _T_2170 = btb_rd_addr_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_2651 = _T_2170 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2906 = _T_2905 | _T_2651; // @[Mux.scala 27:72]
  wire  _T_2172 = btb_rd_addr_f == 8'h20; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_2652 = _T_2172 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2907 = _T_2906 | _T_2652; // @[Mux.scala 27:72]
  wire  _T_2174 = btb_rd_addr_f == 8'h21; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_2653 = _T_2174 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2908 = _T_2907 | _T_2653; // @[Mux.scala 27:72]
  wire  _T_2176 = btb_rd_addr_f == 8'h22; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_2654 = _T_2176 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2909 = _T_2908 | _T_2654; // @[Mux.scala 27:72]
  wire  _T_2178 = btb_rd_addr_f == 8'h23; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_2655 = _T_2178 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2910 = _T_2909 | _T_2655; // @[Mux.scala 27:72]
  wire  _T_2180 = btb_rd_addr_f == 8'h24; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_2656 = _T_2180 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2911 = _T_2910 | _T_2656; // @[Mux.scala 27:72]
  wire  _T_2182 = btb_rd_addr_f == 8'h25; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_2657 = _T_2182 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2912 = _T_2911 | _T_2657; // @[Mux.scala 27:72]
  wire  _T_2184 = btb_rd_addr_f == 8'h26; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_2658 = _T_2184 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2913 = _T_2912 | _T_2658; // @[Mux.scala 27:72]
  wire  _T_2186 = btb_rd_addr_f == 8'h27; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_2659 = _T_2186 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2914 = _T_2913 | _T_2659; // @[Mux.scala 27:72]
  wire  _T_2188 = btb_rd_addr_f == 8'h28; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_2660 = _T_2188 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2915 = _T_2914 | _T_2660; // @[Mux.scala 27:72]
  wire  _T_2190 = btb_rd_addr_f == 8'h29; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_2661 = _T_2190 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2916 = _T_2915 | _T_2661; // @[Mux.scala 27:72]
  wire  _T_2192 = btb_rd_addr_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_2662 = _T_2192 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2917 = _T_2916 | _T_2662; // @[Mux.scala 27:72]
  wire  _T_2194 = btb_rd_addr_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_2663 = _T_2194 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2918 = _T_2917 | _T_2663; // @[Mux.scala 27:72]
  wire  _T_2196 = btb_rd_addr_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_2664 = _T_2196 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2919 = _T_2918 | _T_2664; // @[Mux.scala 27:72]
  wire  _T_2198 = btb_rd_addr_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_2665 = _T_2198 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2920 = _T_2919 | _T_2665; // @[Mux.scala 27:72]
  wire  _T_2200 = btb_rd_addr_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_2666 = _T_2200 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2921 = _T_2920 | _T_2666; // @[Mux.scala 27:72]
  wire  _T_2202 = btb_rd_addr_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_2667 = _T_2202 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2922 = _T_2921 | _T_2667; // @[Mux.scala 27:72]
  wire  _T_2204 = btb_rd_addr_f == 8'h30; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_2668 = _T_2204 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2923 = _T_2922 | _T_2668; // @[Mux.scala 27:72]
  wire  _T_2206 = btb_rd_addr_f == 8'h31; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_2669 = _T_2206 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2924 = _T_2923 | _T_2669; // @[Mux.scala 27:72]
  wire  _T_2208 = btb_rd_addr_f == 8'h32; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_2670 = _T_2208 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2925 = _T_2924 | _T_2670; // @[Mux.scala 27:72]
  wire  _T_2210 = btb_rd_addr_f == 8'h33; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_2671 = _T_2210 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2926 = _T_2925 | _T_2671; // @[Mux.scala 27:72]
  wire  _T_2212 = btb_rd_addr_f == 8'h34; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_2672 = _T_2212 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2927 = _T_2926 | _T_2672; // @[Mux.scala 27:72]
  wire  _T_2214 = btb_rd_addr_f == 8'h35; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_2673 = _T_2214 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2928 = _T_2927 | _T_2673; // @[Mux.scala 27:72]
  wire  _T_2216 = btb_rd_addr_f == 8'h36; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_2674 = _T_2216 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2929 = _T_2928 | _T_2674; // @[Mux.scala 27:72]
  wire  _T_2218 = btb_rd_addr_f == 8'h37; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_2675 = _T_2218 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2930 = _T_2929 | _T_2675; // @[Mux.scala 27:72]
  wire  _T_2220 = btb_rd_addr_f == 8'h38; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_2676 = _T_2220 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2931 = _T_2930 | _T_2676; // @[Mux.scala 27:72]
  wire  _T_2222 = btb_rd_addr_f == 8'h39; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_2677 = _T_2222 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2932 = _T_2931 | _T_2677; // @[Mux.scala 27:72]
  wire  _T_2224 = btb_rd_addr_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_2678 = _T_2224 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2933 = _T_2932 | _T_2678; // @[Mux.scala 27:72]
  wire  _T_2226 = btb_rd_addr_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_2679 = _T_2226 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2934 = _T_2933 | _T_2679; // @[Mux.scala 27:72]
  wire  _T_2228 = btb_rd_addr_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_2680 = _T_2228 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2935 = _T_2934 | _T_2680; // @[Mux.scala 27:72]
  wire  _T_2230 = btb_rd_addr_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_2681 = _T_2230 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2936 = _T_2935 | _T_2681; // @[Mux.scala 27:72]
  wire  _T_2232 = btb_rd_addr_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_2682 = _T_2232 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2937 = _T_2936 | _T_2682; // @[Mux.scala 27:72]
  wire  _T_2234 = btb_rd_addr_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_2683 = _T_2234 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2938 = _T_2937 | _T_2683; // @[Mux.scala 27:72]
  wire  _T_2236 = btb_rd_addr_f == 8'h40; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_2684 = _T_2236 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2939 = _T_2938 | _T_2684; // @[Mux.scala 27:72]
  wire  _T_2238 = btb_rd_addr_f == 8'h41; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_2685 = _T_2238 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2940 = _T_2939 | _T_2685; // @[Mux.scala 27:72]
  wire  _T_2240 = btb_rd_addr_f == 8'h42; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_2686 = _T_2240 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2941 = _T_2940 | _T_2686; // @[Mux.scala 27:72]
  wire  _T_2242 = btb_rd_addr_f == 8'h43; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_2687 = _T_2242 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2942 = _T_2941 | _T_2687; // @[Mux.scala 27:72]
  wire  _T_2244 = btb_rd_addr_f == 8'h44; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_2688 = _T_2244 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2943 = _T_2942 | _T_2688; // @[Mux.scala 27:72]
  wire  _T_2246 = btb_rd_addr_f == 8'h45; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_2689 = _T_2246 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2944 = _T_2943 | _T_2689; // @[Mux.scala 27:72]
  wire  _T_2248 = btb_rd_addr_f == 8'h46; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_2690 = _T_2248 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2945 = _T_2944 | _T_2690; // @[Mux.scala 27:72]
  wire  _T_2250 = btb_rd_addr_f == 8'h47; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_2691 = _T_2250 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2946 = _T_2945 | _T_2691; // @[Mux.scala 27:72]
  wire  _T_2252 = btb_rd_addr_f == 8'h48; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_2692 = _T_2252 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2947 = _T_2946 | _T_2692; // @[Mux.scala 27:72]
  wire  _T_2254 = btb_rd_addr_f == 8'h49; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_2693 = _T_2254 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2948 = _T_2947 | _T_2693; // @[Mux.scala 27:72]
  wire  _T_2256 = btb_rd_addr_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_2694 = _T_2256 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2949 = _T_2948 | _T_2694; // @[Mux.scala 27:72]
  wire  _T_2258 = btb_rd_addr_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_2695 = _T_2258 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2950 = _T_2949 | _T_2695; // @[Mux.scala 27:72]
  wire  _T_2260 = btb_rd_addr_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_2696 = _T_2260 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2951 = _T_2950 | _T_2696; // @[Mux.scala 27:72]
  wire  _T_2262 = btb_rd_addr_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_2697 = _T_2262 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2952 = _T_2951 | _T_2697; // @[Mux.scala 27:72]
  wire  _T_2264 = btb_rd_addr_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_2698 = _T_2264 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2953 = _T_2952 | _T_2698; // @[Mux.scala 27:72]
  wire  _T_2266 = btb_rd_addr_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_2699 = _T_2266 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2954 = _T_2953 | _T_2699; // @[Mux.scala 27:72]
  wire  _T_2268 = btb_rd_addr_f == 8'h50; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_2700 = _T_2268 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2955 = _T_2954 | _T_2700; // @[Mux.scala 27:72]
  wire  _T_2270 = btb_rd_addr_f == 8'h51; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_2701 = _T_2270 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2956 = _T_2955 | _T_2701; // @[Mux.scala 27:72]
  wire  _T_2272 = btb_rd_addr_f == 8'h52; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_2702 = _T_2272 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2957 = _T_2956 | _T_2702; // @[Mux.scala 27:72]
  wire  _T_2274 = btb_rd_addr_f == 8'h53; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_2703 = _T_2274 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2958 = _T_2957 | _T_2703; // @[Mux.scala 27:72]
  wire  _T_2276 = btb_rd_addr_f == 8'h54; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_2704 = _T_2276 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2959 = _T_2958 | _T_2704; // @[Mux.scala 27:72]
  wire  _T_2278 = btb_rd_addr_f == 8'h55; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_2705 = _T_2278 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2960 = _T_2959 | _T_2705; // @[Mux.scala 27:72]
  wire  _T_2280 = btb_rd_addr_f == 8'h56; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_2706 = _T_2280 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2961 = _T_2960 | _T_2706; // @[Mux.scala 27:72]
  wire  _T_2282 = btb_rd_addr_f == 8'h57; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_2707 = _T_2282 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2962 = _T_2961 | _T_2707; // @[Mux.scala 27:72]
  wire  _T_2284 = btb_rd_addr_f == 8'h58; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_2708 = _T_2284 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2963 = _T_2962 | _T_2708; // @[Mux.scala 27:72]
  wire  _T_2286 = btb_rd_addr_f == 8'h59; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_2709 = _T_2286 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2964 = _T_2963 | _T_2709; // @[Mux.scala 27:72]
  wire  _T_2288 = btb_rd_addr_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_2710 = _T_2288 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2965 = _T_2964 | _T_2710; // @[Mux.scala 27:72]
  wire  _T_2290 = btb_rd_addr_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_2711 = _T_2290 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2966 = _T_2965 | _T_2711; // @[Mux.scala 27:72]
  wire  _T_2292 = btb_rd_addr_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_2712 = _T_2292 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2967 = _T_2966 | _T_2712; // @[Mux.scala 27:72]
  wire  _T_2294 = btb_rd_addr_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_2713 = _T_2294 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2968 = _T_2967 | _T_2713; // @[Mux.scala 27:72]
  wire  _T_2296 = btb_rd_addr_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_2714 = _T_2296 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2969 = _T_2968 | _T_2714; // @[Mux.scala 27:72]
  wire  _T_2298 = btb_rd_addr_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_2715 = _T_2298 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2970 = _T_2969 | _T_2715; // @[Mux.scala 27:72]
  wire  _T_2300 = btb_rd_addr_f == 8'h60; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_2716 = _T_2300 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2971 = _T_2970 | _T_2716; // @[Mux.scala 27:72]
  wire  _T_2302 = btb_rd_addr_f == 8'h61; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_2717 = _T_2302 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2972 = _T_2971 | _T_2717; // @[Mux.scala 27:72]
  wire  _T_2304 = btb_rd_addr_f == 8'h62; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_2718 = _T_2304 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2973 = _T_2972 | _T_2718; // @[Mux.scala 27:72]
  wire  _T_2306 = btb_rd_addr_f == 8'h63; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_2719 = _T_2306 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2974 = _T_2973 | _T_2719; // @[Mux.scala 27:72]
  wire  _T_2308 = btb_rd_addr_f == 8'h64; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_2720 = _T_2308 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2975 = _T_2974 | _T_2720; // @[Mux.scala 27:72]
  wire  _T_2310 = btb_rd_addr_f == 8'h65; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_2721 = _T_2310 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2976 = _T_2975 | _T_2721; // @[Mux.scala 27:72]
  wire  _T_2312 = btb_rd_addr_f == 8'h66; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_2722 = _T_2312 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2977 = _T_2976 | _T_2722; // @[Mux.scala 27:72]
  wire  _T_2314 = btb_rd_addr_f == 8'h67; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_2723 = _T_2314 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2978 = _T_2977 | _T_2723; // @[Mux.scala 27:72]
  wire  _T_2316 = btb_rd_addr_f == 8'h68; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_2724 = _T_2316 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2979 = _T_2978 | _T_2724; // @[Mux.scala 27:72]
  wire  _T_2318 = btb_rd_addr_f == 8'h69; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_2725 = _T_2318 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2980 = _T_2979 | _T_2725; // @[Mux.scala 27:72]
  wire  _T_2320 = btb_rd_addr_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_2726 = _T_2320 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2981 = _T_2980 | _T_2726; // @[Mux.scala 27:72]
  wire  _T_2322 = btb_rd_addr_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_2727 = _T_2322 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2982 = _T_2981 | _T_2727; // @[Mux.scala 27:72]
  wire  _T_2324 = btb_rd_addr_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_2728 = _T_2324 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2983 = _T_2982 | _T_2728; // @[Mux.scala 27:72]
  wire  _T_2326 = btb_rd_addr_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_2729 = _T_2326 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2984 = _T_2983 | _T_2729; // @[Mux.scala 27:72]
  wire  _T_2328 = btb_rd_addr_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_2730 = _T_2328 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2985 = _T_2984 | _T_2730; // @[Mux.scala 27:72]
  wire  _T_2330 = btb_rd_addr_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_2731 = _T_2330 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2986 = _T_2985 | _T_2731; // @[Mux.scala 27:72]
  wire  _T_2332 = btb_rd_addr_f == 8'h70; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_2732 = _T_2332 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2987 = _T_2986 | _T_2732; // @[Mux.scala 27:72]
  wire  _T_2334 = btb_rd_addr_f == 8'h71; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_2733 = _T_2334 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2988 = _T_2987 | _T_2733; // @[Mux.scala 27:72]
  wire  _T_2336 = btb_rd_addr_f == 8'h72; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_2734 = _T_2336 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2989 = _T_2988 | _T_2734; // @[Mux.scala 27:72]
  wire  _T_2338 = btb_rd_addr_f == 8'h73; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_2735 = _T_2338 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2990 = _T_2989 | _T_2735; // @[Mux.scala 27:72]
  wire  _T_2340 = btb_rd_addr_f == 8'h74; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_2736 = _T_2340 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2991 = _T_2990 | _T_2736; // @[Mux.scala 27:72]
  wire  _T_2342 = btb_rd_addr_f == 8'h75; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_2737 = _T_2342 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2992 = _T_2991 | _T_2737; // @[Mux.scala 27:72]
  wire  _T_2344 = btb_rd_addr_f == 8'h76; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_2738 = _T_2344 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2993 = _T_2992 | _T_2738; // @[Mux.scala 27:72]
  wire  _T_2346 = btb_rd_addr_f == 8'h77; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_2739 = _T_2346 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2994 = _T_2993 | _T_2739; // @[Mux.scala 27:72]
  wire  _T_2348 = btb_rd_addr_f == 8'h78; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_2740 = _T_2348 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2995 = _T_2994 | _T_2740; // @[Mux.scala 27:72]
  wire  _T_2350 = btb_rd_addr_f == 8'h79; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_2741 = _T_2350 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2996 = _T_2995 | _T_2741; // @[Mux.scala 27:72]
  wire  _T_2352 = btb_rd_addr_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_2742 = _T_2352 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2997 = _T_2996 | _T_2742; // @[Mux.scala 27:72]
  wire  _T_2354 = btb_rd_addr_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_2743 = _T_2354 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2998 = _T_2997 | _T_2743; // @[Mux.scala 27:72]
  wire  _T_2356 = btb_rd_addr_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_2744 = _T_2356 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2999 = _T_2998 | _T_2744; // @[Mux.scala 27:72]
  wire  _T_2358 = btb_rd_addr_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_2745 = _T_2358 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3000 = _T_2999 | _T_2745; // @[Mux.scala 27:72]
  wire  _T_2360 = btb_rd_addr_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_2746 = _T_2360 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3001 = _T_3000 | _T_2746; // @[Mux.scala 27:72]
  wire  _T_2362 = btb_rd_addr_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_2747 = _T_2362 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3002 = _T_3001 | _T_2747; // @[Mux.scala 27:72]
  wire  _T_2364 = btb_rd_addr_f == 8'h80; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_2748 = _T_2364 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3003 = _T_3002 | _T_2748; // @[Mux.scala 27:72]
  wire  _T_2366 = btb_rd_addr_f == 8'h81; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_2749 = _T_2366 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3004 = _T_3003 | _T_2749; // @[Mux.scala 27:72]
  wire  _T_2368 = btb_rd_addr_f == 8'h82; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_2750 = _T_2368 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3005 = _T_3004 | _T_2750; // @[Mux.scala 27:72]
  wire  _T_2370 = btb_rd_addr_f == 8'h83; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_2751 = _T_2370 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3006 = _T_3005 | _T_2751; // @[Mux.scala 27:72]
  wire  _T_2372 = btb_rd_addr_f == 8'h84; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_2752 = _T_2372 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3007 = _T_3006 | _T_2752; // @[Mux.scala 27:72]
  wire  _T_2374 = btb_rd_addr_f == 8'h85; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_2753 = _T_2374 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3008 = _T_3007 | _T_2753; // @[Mux.scala 27:72]
  wire  _T_2376 = btb_rd_addr_f == 8'h86; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_2754 = _T_2376 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3009 = _T_3008 | _T_2754; // @[Mux.scala 27:72]
  wire  _T_2378 = btb_rd_addr_f == 8'h87; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_2755 = _T_2378 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3010 = _T_3009 | _T_2755; // @[Mux.scala 27:72]
  wire  _T_2380 = btb_rd_addr_f == 8'h88; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_2756 = _T_2380 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3011 = _T_3010 | _T_2756; // @[Mux.scala 27:72]
  wire  _T_2382 = btb_rd_addr_f == 8'h89; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_2757 = _T_2382 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3012 = _T_3011 | _T_2757; // @[Mux.scala 27:72]
  wire  _T_2384 = btb_rd_addr_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_2758 = _T_2384 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3013 = _T_3012 | _T_2758; // @[Mux.scala 27:72]
  wire  _T_2386 = btb_rd_addr_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_2759 = _T_2386 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3014 = _T_3013 | _T_2759; // @[Mux.scala 27:72]
  wire  _T_2388 = btb_rd_addr_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_2760 = _T_2388 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3015 = _T_3014 | _T_2760; // @[Mux.scala 27:72]
  wire  _T_2390 = btb_rd_addr_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_2761 = _T_2390 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3016 = _T_3015 | _T_2761; // @[Mux.scala 27:72]
  wire  _T_2392 = btb_rd_addr_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_2762 = _T_2392 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3017 = _T_3016 | _T_2762; // @[Mux.scala 27:72]
  wire  _T_2394 = btb_rd_addr_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_2763 = _T_2394 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3018 = _T_3017 | _T_2763; // @[Mux.scala 27:72]
  wire  _T_2396 = btb_rd_addr_f == 8'h90; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_2764 = _T_2396 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3019 = _T_3018 | _T_2764; // @[Mux.scala 27:72]
  wire  _T_2398 = btb_rd_addr_f == 8'h91; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_2765 = _T_2398 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3020 = _T_3019 | _T_2765; // @[Mux.scala 27:72]
  wire  _T_2400 = btb_rd_addr_f == 8'h92; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_2766 = _T_2400 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3021 = _T_3020 | _T_2766; // @[Mux.scala 27:72]
  wire  _T_2402 = btb_rd_addr_f == 8'h93; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_2767 = _T_2402 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3022 = _T_3021 | _T_2767; // @[Mux.scala 27:72]
  wire  _T_2404 = btb_rd_addr_f == 8'h94; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_2768 = _T_2404 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3023 = _T_3022 | _T_2768; // @[Mux.scala 27:72]
  wire  _T_2406 = btb_rd_addr_f == 8'h95; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_2769 = _T_2406 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3024 = _T_3023 | _T_2769; // @[Mux.scala 27:72]
  wire  _T_2408 = btb_rd_addr_f == 8'h96; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_2770 = _T_2408 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3025 = _T_3024 | _T_2770; // @[Mux.scala 27:72]
  wire  _T_2410 = btb_rd_addr_f == 8'h97; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_2771 = _T_2410 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3026 = _T_3025 | _T_2771; // @[Mux.scala 27:72]
  wire  _T_2412 = btb_rd_addr_f == 8'h98; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_2772 = _T_2412 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3027 = _T_3026 | _T_2772; // @[Mux.scala 27:72]
  wire  _T_2414 = btb_rd_addr_f == 8'h99; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_2773 = _T_2414 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3028 = _T_3027 | _T_2773; // @[Mux.scala 27:72]
  wire  _T_2416 = btb_rd_addr_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_2774 = _T_2416 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3029 = _T_3028 | _T_2774; // @[Mux.scala 27:72]
  wire  _T_2418 = btb_rd_addr_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_2775 = _T_2418 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3030 = _T_3029 | _T_2775; // @[Mux.scala 27:72]
  wire  _T_2420 = btb_rd_addr_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_2776 = _T_2420 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3031 = _T_3030 | _T_2776; // @[Mux.scala 27:72]
  wire  _T_2422 = btb_rd_addr_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_2777 = _T_2422 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3032 = _T_3031 | _T_2777; // @[Mux.scala 27:72]
  wire  _T_2424 = btb_rd_addr_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_2778 = _T_2424 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3033 = _T_3032 | _T_2778; // @[Mux.scala 27:72]
  wire  _T_2426 = btb_rd_addr_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_2779 = _T_2426 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3034 = _T_3033 | _T_2779; // @[Mux.scala 27:72]
  wire  _T_2428 = btb_rd_addr_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_2780 = _T_2428 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3035 = _T_3034 | _T_2780; // @[Mux.scala 27:72]
  wire  _T_2430 = btb_rd_addr_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_2781 = _T_2430 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3036 = _T_3035 | _T_2781; // @[Mux.scala 27:72]
  wire  _T_2432 = btb_rd_addr_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_2782 = _T_2432 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3037 = _T_3036 | _T_2782; // @[Mux.scala 27:72]
  wire  _T_2434 = btb_rd_addr_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_2783 = _T_2434 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3038 = _T_3037 | _T_2783; // @[Mux.scala 27:72]
  wire  _T_2436 = btb_rd_addr_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_2784 = _T_2436 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3039 = _T_3038 | _T_2784; // @[Mux.scala 27:72]
  wire  _T_2438 = btb_rd_addr_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_2785 = _T_2438 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3040 = _T_3039 | _T_2785; // @[Mux.scala 27:72]
  wire  _T_2440 = btb_rd_addr_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_2786 = _T_2440 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3041 = _T_3040 | _T_2786; // @[Mux.scala 27:72]
  wire  _T_2442 = btb_rd_addr_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_2787 = _T_2442 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3042 = _T_3041 | _T_2787; // @[Mux.scala 27:72]
  wire  _T_2444 = btb_rd_addr_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_2788 = _T_2444 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3043 = _T_3042 | _T_2788; // @[Mux.scala 27:72]
  wire  _T_2446 = btb_rd_addr_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_2789 = _T_2446 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3044 = _T_3043 | _T_2789; // @[Mux.scala 27:72]
  wire  _T_2448 = btb_rd_addr_f == 8'haa; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_2790 = _T_2448 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3045 = _T_3044 | _T_2790; // @[Mux.scala 27:72]
  wire  _T_2450 = btb_rd_addr_f == 8'hab; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_2791 = _T_2450 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3046 = _T_3045 | _T_2791; // @[Mux.scala 27:72]
  wire  _T_2452 = btb_rd_addr_f == 8'hac; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_2792 = _T_2452 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3047 = _T_3046 | _T_2792; // @[Mux.scala 27:72]
  wire  _T_2454 = btb_rd_addr_f == 8'had; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_2793 = _T_2454 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3048 = _T_3047 | _T_2793; // @[Mux.scala 27:72]
  wire  _T_2456 = btb_rd_addr_f == 8'hae; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_2794 = _T_2456 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3049 = _T_3048 | _T_2794; // @[Mux.scala 27:72]
  wire  _T_2458 = btb_rd_addr_f == 8'haf; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_2795 = _T_2458 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3050 = _T_3049 | _T_2795; // @[Mux.scala 27:72]
  wire  _T_2460 = btb_rd_addr_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_2796 = _T_2460 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3051 = _T_3050 | _T_2796; // @[Mux.scala 27:72]
  wire  _T_2462 = btb_rd_addr_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_2797 = _T_2462 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3052 = _T_3051 | _T_2797; // @[Mux.scala 27:72]
  wire  _T_2464 = btb_rd_addr_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_2798 = _T_2464 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3053 = _T_3052 | _T_2798; // @[Mux.scala 27:72]
  wire  _T_2466 = btb_rd_addr_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_2799 = _T_2466 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3054 = _T_3053 | _T_2799; // @[Mux.scala 27:72]
  wire  _T_2468 = btb_rd_addr_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_2800 = _T_2468 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3055 = _T_3054 | _T_2800; // @[Mux.scala 27:72]
  wire  _T_2470 = btb_rd_addr_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_2801 = _T_2470 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3056 = _T_3055 | _T_2801; // @[Mux.scala 27:72]
  wire  _T_2472 = btb_rd_addr_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_2802 = _T_2472 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3057 = _T_3056 | _T_2802; // @[Mux.scala 27:72]
  wire  _T_2474 = btb_rd_addr_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_2803 = _T_2474 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3058 = _T_3057 | _T_2803; // @[Mux.scala 27:72]
  wire  _T_2476 = btb_rd_addr_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_2804 = _T_2476 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3059 = _T_3058 | _T_2804; // @[Mux.scala 27:72]
  wire  _T_2478 = btb_rd_addr_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_2805 = _T_2478 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3060 = _T_3059 | _T_2805; // @[Mux.scala 27:72]
  wire  _T_2480 = btb_rd_addr_f == 8'hba; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_2806 = _T_2480 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3061 = _T_3060 | _T_2806; // @[Mux.scala 27:72]
  wire  _T_2482 = btb_rd_addr_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_2807 = _T_2482 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3062 = _T_3061 | _T_2807; // @[Mux.scala 27:72]
  wire  _T_2484 = btb_rd_addr_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_2808 = _T_2484 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3063 = _T_3062 | _T_2808; // @[Mux.scala 27:72]
  wire  _T_2486 = btb_rd_addr_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_2809 = _T_2486 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3064 = _T_3063 | _T_2809; // @[Mux.scala 27:72]
  wire  _T_2488 = btb_rd_addr_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_2810 = _T_2488 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3065 = _T_3064 | _T_2810; // @[Mux.scala 27:72]
  wire  _T_2490 = btb_rd_addr_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_2811 = _T_2490 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3066 = _T_3065 | _T_2811; // @[Mux.scala 27:72]
  wire  _T_2492 = btb_rd_addr_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_2812 = _T_2492 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3067 = _T_3066 | _T_2812; // @[Mux.scala 27:72]
  wire  _T_2494 = btb_rd_addr_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_2813 = _T_2494 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3068 = _T_3067 | _T_2813; // @[Mux.scala 27:72]
  wire  _T_2496 = btb_rd_addr_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_2814 = _T_2496 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3069 = _T_3068 | _T_2814; // @[Mux.scala 27:72]
  wire  _T_2498 = btb_rd_addr_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_2815 = _T_2498 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3070 = _T_3069 | _T_2815; // @[Mux.scala 27:72]
  wire  _T_2500 = btb_rd_addr_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_2816 = _T_2500 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3071 = _T_3070 | _T_2816; // @[Mux.scala 27:72]
  wire  _T_2502 = btb_rd_addr_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_2817 = _T_2502 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3072 = _T_3071 | _T_2817; // @[Mux.scala 27:72]
  wire  _T_2504 = btb_rd_addr_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_2818 = _T_2504 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3073 = _T_3072 | _T_2818; // @[Mux.scala 27:72]
  wire  _T_2506 = btb_rd_addr_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_2819 = _T_2506 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3074 = _T_3073 | _T_2819; // @[Mux.scala 27:72]
  wire  _T_2508 = btb_rd_addr_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_2820 = _T_2508 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3075 = _T_3074 | _T_2820; // @[Mux.scala 27:72]
  wire  _T_2510 = btb_rd_addr_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_2821 = _T_2510 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3076 = _T_3075 | _T_2821; // @[Mux.scala 27:72]
  wire  _T_2512 = btb_rd_addr_f == 8'hca; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_2822 = _T_2512 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3077 = _T_3076 | _T_2822; // @[Mux.scala 27:72]
  wire  _T_2514 = btb_rd_addr_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_2823 = _T_2514 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3078 = _T_3077 | _T_2823; // @[Mux.scala 27:72]
  wire  _T_2516 = btb_rd_addr_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_2824 = _T_2516 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3079 = _T_3078 | _T_2824; // @[Mux.scala 27:72]
  wire  _T_2518 = btb_rd_addr_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_2825 = _T_2518 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3080 = _T_3079 | _T_2825; // @[Mux.scala 27:72]
  wire  _T_2520 = btb_rd_addr_f == 8'hce; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_2826 = _T_2520 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3081 = _T_3080 | _T_2826; // @[Mux.scala 27:72]
  wire  _T_2522 = btb_rd_addr_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_2827 = _T_2522 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3082 = _T_3081 | _T_2827; // @[Mux.scala 27:72]
  wire  _T_2524 = btb_rd_addr_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_2828 = _T_2524 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3083 = _T_3082 | _T_2828; // @[Mux.scala 27:72]
  wire  _T_2526 = btb_rd_addr_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_2829 = _T_2526 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3084 = _T_3083 | _T_2829; // @[Mux.scala 27:72]
  wire  _T_2528 = btb_rd_addr_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_2830 = _T_2528 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3085 = _T_3084 | _T_2830; // @[Mux.scala 27:72]
  wire  _T_2530 = btb_rd_addr_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_2831 = _T_2530 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3086 = _T_3085 | _T_2831; // @[Mux.scala 27:72]
  wire  _T_2532 = btb_rd_addr_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_2832 = _T_2532 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3087 = _T_3086 | _T_2832; // @[Mux.scala 27:72]
  wire  _T_2534 = btb_rd_addr_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_2833 = _T_2534 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3088 = _T_3087 | _T_2833; // @[Mux.scala 27:72]
  wire  _T_2536 = btb_rd_addr_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_2834 = _T_2536 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3089 = _T_3088 | _T_2834; // @[Mux.scala 27:72]
  wire  _T_2538 = btb_rd_addr_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_2835 = _T_2538 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3090 = _T_3089 | _T_2835; // @[Mux.scala 27:72]
  wire  _T_2540 = btb_rd_addr_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_2836 = _T_2540 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3091 = _T_3090 | _T_2836; // @[Mux.scala 27:72]
  wire  _T_2542 = btb_rd_addr_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_2837 = _T_2542 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3092 = _T_3091 | _T_2837; // @[Mux.scala 27:72]
  wire  _T_2544 = btb_rd_addr_f == 8'hda; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_2838 = _T_2544 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3093 = _T_3092 | _T_2838; // @[Mux.scala 27:72]
  wire  _T_2546 = btb_rd_addr_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_2839 = _T_2546 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3094 = _T_3093 | _T_2839; // @[Mux.scala 27:72]
  wire  _T_2548 = btb_rd_addr_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_2840 = _T_2548 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3095 = _T_3094 | _T_2840; // @[Mux.scala 27:72]
  wire  _T_2550 = btb_rd_addr_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_2841 = _T_2550 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3096 = _T_3095 | _T_2841; // @[Mux.scala 27:72]
  wire  _T_2552 = btb_rd_addr_f == 8'hde; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_2842 = _T_2552 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3097 = _T_3096 | _T_2842; // @[Mux.scala 27:72]
  wire  _T_2554 = btb_rd_addr_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_2843 = _T_2554 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3098 = _T_3097 | _T_2843; // @[Mux.scala 27:72]
  wire  _T_2556 = btb_rd_addr_f == 8'he0; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_2844 = _T_2556 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3099 = _T_3098 | _T_2844; // @[Mux.scala 27:72]
  wire  _T_2558 = btb_rd_addr_f == 8'he1; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_2845 = _T_2558 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3100 = _T_3099 | _T_2845; // @[Mux.scala 27:72]
  wire  _T_2560 = btb_rd_addr_f == 8'he2; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_2846 = _T_2560 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3101 = _T_3100 | _T_2846; // @[Mux.scala 27:72]
  wire  _T_2562 = btb_rd_addr_f == 8'he3; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_2847 = _T_2562 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3102 = _T_3101 | _T_2847; // @[Mux.scala 27:72]
  wire  _T_2564 = btb_rd_addr_f == 8'he4; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_2848 = _T_2564 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3103 = _T_3102 | _T_2848; // @[Mux.scala 27:72]
  wire  _T_2566 = btb_rd_addr_f == 8'he5; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_2849 = _T_2566 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3104 = _T_3103 | _T_2849; // @[Mux.scala 27:72]
  wire  _T_2568 = btb_rd_addr_f == 8'he6; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_2850 = _T_2568 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3105 = _T_3104 | _T_2850; // @[Mux.scala 27:72]
  wire  _T_2570 = btb_rd_addr_f == 8'he7; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_2851 = _T_2570 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3106 = _T_3105 | _T_2851; // @[Mux.scala 27:72]
  wire  _T_2572 = btb_rd_addr_f == 8'he8; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_2852 = _T_2572 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3107 = _T_3106 | _T_2852; // @[Mux.scala 27:72]
  wire  _T_2574 = btb_rd_addr_f == 8'he9; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_2853 = _T_2574 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3108 = _T_3107 | _T_2853; // @[Mux.scala 27:72]
  wire  _T_2576 = btb_rd_addr_f == 8'hea; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_2854 = _T_2576 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3109 = _T_3108 | _T_2854; // @[Mux.scala 27:72]
  wire  _T_2578 = btb_rd_addr_f == 8'heb; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_2855 = _T_2578 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3110 = _T_3109 | _T_2855; // @[Mux.scala 27:72]
  wire  _T_2580 = btb_rd_addr_f == 8'hec; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_2856 = _T_2580 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3111 = _T_3110 | _T_2856; // @[Mux.scala 27:72]
  wire  _T_2582 = btb_rd_addr_f == 8'hed; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_2857 = _T_2582 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3112 = _T_3111 | _T_2857; // @[Mux.scala 27:72]
  wire  _T_2584 = btb_rd_addr_f == 8'hee; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_2858 = _T_2584 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3113 = _T_3112 | _T_2858; // @[Mux.scala 27:72]
  wire  _T_2586 = btb_rd_addr_f == 8'hef; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_2859 = _T_2586 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3114 = _T_3113 | _T_2859; // @[Mux.scala 27:72]
  wire  _T_2588 = btb_rd_addr_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_2860 = _T_2588 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3115 = _T_3114 | _T_2860; // @[Mux.scala 27:72]
  wire  _T_2590 = btb_rd_addr_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_2861 = _T_2590 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3116 = _T_3115 | _T_2861; // @[Mux.scala 27:72]
  wire  _T_2592 = btb_rd_addr_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_2862 = _T_2592 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3117 = _T_3116 | _T_2862; // @[Mux.scala 27:72]
  wire  _T_2594 = btb_rd_addr_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_2863 = _T_2594 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3118 = _T_3117 | _T_2863; // @[Mux.scala 27:72]
  wire  _T_2596 = btb_rd_addr_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_2864 = _T_2596 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3119 = _T_3118 | _T_2864; // @[Mux.scala 27:72]
  wire  _T_2598 = btb_rd_addr_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_2865 = _T_2598 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3120 = _T_3119 | _T_2865; // @[Mux.scala 27:72]
  wire  _T_2600 = btb_rd_addr_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_2866 = _T_2600 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3121 = _T_3120 | _T_2866; // @[Mux.scala 27:72]
  wire  _T_2602 = btb_rd_addr_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_2867 = _T_2602 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3122 = _T_3121 | _T_2867; // @[Mux.scala 27:72]
  wire  _T_2604 = btb_rd_addr_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_2868 = _T_2604 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3123 = _T_3122 | _T_2868; // @[Mux.scala 27:72]
  wire  _T_2606 = btb_rd_addr_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_2869 = _T_2606 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3124 = _T_3123 | _T_2869; // @[Mux.scala 27:72]
  wire  _T_2608 = btb_rd_addr_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_2870 = _T_2608 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3125 = _T_3124 | _T_2870; // @[Mux.scala 27:72]
  wire  _T_2610 = btb_rd_addr_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_2871 = _T_2610 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3126 = _T_3125 | _T_2871; // @[Mux.scala 27:72]
  wire  _T_2612 = btb_rd_addr_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_2872 = _T_2612 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3127 = _T_3126 | _T_2872; // @[Mux.scala 27:72]
  wire  _T_2614 = btb_rd_addr_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_2873 = _T_2614 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3128 = _T_3127 | _T_2873; // @[Mux.scala 27:72]
  wire  _T_2616 = btb_rd_addr_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_2874 = _T_2616 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3129 = _T_3128 | _T_2874; // @[Mux.scala 27:72]
  wire  _T_2618 = btb_rd_addr_f == 8'hff; // @[el2_ifu_bp_ctl.scala 369:77]
  reg [21:0] btb_bank0_rd_data_way0_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_2875 = _T_2618 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3129 | _T_2875; // @[Mux.scala 27:72]
  wire [4:0] _T_25 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[el2_lib.scala 174:111]
  wire [4:0] fetch_rd_tag_f = _T_25 ^ io_ifc_fetch_addr_f[23:19]; // @[el2_lib.scala 174:111]
  wire  _T_45 = btb_bank0_rd_data_way0_f[21:17] == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 136:97]
  wire  _T_46 = btb_bank0_rd_data_way0_f[0] & _T_45; // @[el2_ifu_bp_ctl.scala 136:55]
  reg  dec_tlu_way_wb_f; // @[el2_ifu_bp_ctl.scala 128:33]
  wire [6:0] btb_error_addr_wb = io_exu_i0_br_index_r[6:0]; // @[el2_ifu_bp_ctl.scala 96:21]
  wire [7:0] _GEN_1034 = {{1'd0}, btb_error_addr_wb}; // @[el2_ifu_bp_ctl.scala 114:72]
  wire  _T_19 = _GEN_1034 == btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 114:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[el2_ifu_bp_ctl.scala 114:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 118:63]
  wire  _T_47 = dec_tlu_way_wb_f & branch_error_bank_conflict_f; // @[el2_ifu_bp_ctl.scala 137:22]
  wire  _T_48 = ~_T_47; // @[el2_ifu_bp_ctl.scala 137:3]
  wire  _T_49 = _T_46 & _T_48; // @[el2_ifu_bp_ctl.scala 136:117]
  wire  _T_50 = _T_49 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 137:54]
  wire  tag_match_way0_f = _T_50 & _T; // @[el2_ifu_bp_ctl.scala 137:75]
  wire  _T_81 = btb_bank0_rd_data_way0_f[3] ^ btb_bank0_rd_data_way0_f[4]; // @[el2_ifu_bp_ctl.scala 149:91]
  wire  _T_82 = tag_match_way0_f & _T_81; // @[el2_ifu_bp_ctl.scala 149:56]
  wire  _T_86 = ~_T_81; // @[el2_ifu_bp_ctl.scala 150:58]
  wire  _T_87 = tag_match_way0_f & _T_86; // @[el2_ifu_bp_ctl.scala 150:56]
  wire [1:0] tag_match_way0_expanded_f = {_T_82,_T_87}; // @[Cat.scala 29:58]
  wire [21:0] _T_126 = tag_match_way0_expanded_f[1] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_3644 = _T_2108 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_3645 = _T_2110 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3900 = _T_3644 | _T_3645; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_3646 = _T_2112 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3901 = _T_3900 | _T_3646; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_3647 = _T_2114 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3902 = _T_3901 | _T_3647; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_3648 = _T_2116 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3903 = _T_3902 | _T_3648; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_3649 = _T_2118 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3904 = _T_3903 | _T_3649; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_3650 = _T_2120 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3905 = _T_3904 | _T_3650; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_3651 = _T_2122 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3906 = _T_3905 | _T_3651; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_3652 = _T_2124 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3907 = _T_3906 | _T_3652; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_3653 = _T_2126 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3908 = _T_3907 | _T_3653; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_3654 = _T_2128 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3909 = _T_3908 | _T_3654; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_3655 = _T_2130 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3910 = _T_3909 | _T_3655; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_3656 = _T_2132 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3911 = _T_3910 | _T_3656; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_3657 = _T_2134 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3912 = _T_3911 | _T_3657; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_3658 = _T_2136 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3913 = _T_3912 | _T_3658; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_3659 = _T_2138 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3914 = _T_3913 | _T_3659; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_3660 = _T_2140 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3915 = _T_3914 | _T_3660; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_3661 = _T_2142 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3916 = _T_3915 | _T_3661; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_3662 = _T_2144 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3917 = _T_3916 | _T_3662; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_3663 = _T_2146 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3918 = _T_3917 | _T_3663; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_3664 = _T_2148 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3919 = _T_3918 | _T_3664; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_3665 = _T_2150 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3920 = _T_3919 | _T_3665; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_3666 = _T_2152 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3921 = _T_3920 | _T_3666; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_3667 = _T_2154 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3922 = _T_3921 | _T_3667; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_3668 = _T_2156 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3923 = _T_3922 | _T_3668; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_3669 = _T_2158 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3924 = _T_3923 | _T_3669; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_3670 = _T_2160 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3925 = _T_3924 | _T_3670; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_3671 = _T_2162 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3926 = _T_3925 | _T_3671; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_3672 = _T_2164 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3927 = _T_3926 | _T_3672; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_3673 = _T_2166 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3928 = _T_3927 | _T_3673; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_3674 = _T_2168 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3929 = _T_3928 | _T_3674; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_3675 = _T_2170 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3930 = _T_3929 | _T_3675; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_3676 = _T_2172 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3931 = _T_3930 | _T_3676; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_3677 = _T_2174 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3932 = _T_3931 | _T_3677; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_3678 = _T_2176 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3933 = _T_3932 | _T_3678; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_3679 = _T_2178 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3934 = _T_3933 | _T_3679; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_3680 = _T_2180 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3935 = _T_3934 | _T_3680; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_3681 = _T_2182 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3936 = _T_3935 | _T_3681; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_3682 = _T_2184 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3937 = _T_3936 | _T_3682; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_3683 = _T_2186 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3938 = _T_3937 | _T_3683; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_3684 = _T_2188 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3939 = _T_3938 | _T_3684; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_3685 = _T_2190 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3940 = _T_3939 | _T_3685; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_3686 = _T_2192 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3941 = _T_3940 | _T_3686; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_3687 = _T_2194 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3942 = _T_3941 | _T_3687; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_3688 = _T_2196 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3943 = _T_3942 | _T_3688; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_3689 = _T_2198 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3944 = _T_3943 | _T_3689; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_3690 = _T_2200 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3945 = _T_3944 | _T_3690; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_3691 = _T_2202 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3946 = _T_3945 | _T_3691; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_3692 = _T_2204 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3947 = _T_3946 | _T_3692; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_3693 = _T_2206 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3948 = _T_3947 | _T_3693; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_3694 = _T_2208 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3949 = _T_3948 | _T_3694; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_3695 = _T_2210 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3950 = _T_3949 | _T_3695; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_3696 = _T_2212 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3951 = _T_3950 | _T_3696; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_3697 = _T_2214 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3952 = _T_3951 | _T_3697; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_3698 = _T_2216 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3953 = _T_3952 | _T_3698; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_3699 = _T_2218 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3954 = _T_3953 | _T_3699; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_3700 = _T_2220 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3955 = _T_3954 | _T_3700; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_3701 = _T_2222 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3956 = _T_3955 | _T_3701; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_3702 = _T_2224 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3957 = _T_3956 | _T_3702; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_3703 = _T_2226 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3958 = _T_3957 | _T_3703; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_3704 = _T_2228 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3959 = _T_3958 | _T_3704; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_3705 = _T_2230 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3960 = _T_3959 | _T_3705; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_3706 = _T_2232 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3961 = _T_3960 | _T_3706; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_3707 = _T_2234 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3962 = _T_3961 | _T_3707; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_3708 = _T_2236 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3963 = _T_3962 | _T_3708; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_3709 = _T_2238 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3964 = _T_3963 | _T_3709; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_3710 = _T_2240 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3965 = _T_3964 | _T_3710; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_3711 = _T_2242 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3966 = _T_3965 | _T_3711; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_3712 = _T_2244 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3967 = _T_3966 | _T_3712; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_3713 = _T_2246 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3968 = _T_3967 | _T_3713; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_3714 = _T_2248 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3969 = _T_3968 | _T_3714; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_3715 = _T_2250 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3970 = _T_3969 | _T_3715; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_3716 = _T_2252 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3971 = _T_3970 | _T_3716; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_3717 = _T_2254 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3972 = _T_3971 | _T_3717; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_3718 = _T_2256 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3973 = _T_3972 | _T_3718; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_3719 = _T_2258 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3974 = _T_3973 | _T_3719; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_3720 = _T_2260 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3975 = _T_3974 | _T_3720; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_3721 = _T_2262 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3976 = _T_3975 | _T_3721; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_3722 = _T_2264 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3977 = _T_3976 | _T_3722; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_3723 = _T_2266 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3978 = _T_3977 | _T_3723; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_3724 = _T_2268 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3979 = _T_3978 | _T_3724; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_3725 = _T_2270 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3980 = _T_3979 | _T_3725; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_3726 = _T_2272 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3981 = _T_3980 | _T_3726; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_3727 = _T_2274 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3982 = _T_3981 | _T_3727; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_3728 = _T_2276 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3983 = _T_3982 | _T_3728; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_3729 = _T_2278 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3984 = _T_3983 | _T_3729; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_3730 = _T_2280 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3985 = _T_3984 | _T_3730; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_3731 = _T_2282 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3986 = _T_3985 | _T_3731; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_3732 = _T_2284 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3987 = _T_3986 | _T_3732; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_3733 = _T_2286 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3988 = _T_3987 | _T_3733; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_3734 = _T_2288 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3989 = _T_3988 | _T_3734; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_3735 = _T_2290 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3990 = _T_3989 | _T_3735; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_3736 = _T_2292 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3991 = _T_3990 | _T_3736; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_3737 = _T_2294 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3992 = _T_3991 | _T_3737; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_3738 = _T_2296 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3993 = _T_3992 | _T_3738; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_3739 = _T_2298 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3994 = _T_3993 | _T_3739; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_3740 = _T_2300 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3995 = _T_3994 | _T_3740; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_3741 = _T_2302 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3996 = _T_3995 | _T_3741; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_3742 = _T_2304 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3997 = _T_3996 | _T_3742; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_3743 = _T_2306 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3998 = _T_3997 | _T_3743; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_3744 = _T_2308 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3999 = _T_3998 | _T_3744; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_3745 = _T_2310 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4000 = _T_3999 | _T_3745; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_3746 = _T_2312 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4001 = _T_4000 | _T_3746; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_3747 = _T_2314 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4002 = _T_4001 | _T_3747; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_3748 = _T_2316 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4003 = _T_4002 | _T_3748; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_3749 = _T_2318 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4004 = _T_4003 | _T_3749; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_3750 = _T_2320 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4005 = _T_4004 | _T_3750; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_3751 = _T_2322 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4006 = _T_4005 | _T_3751; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_3752 = _T_2324 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4007 = _T_4006 | _T_3752; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_3753 = _T_2326 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4008 = _T_4007 | _T_3753; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_3754 = _T_2328 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4009 = _T_4008 | _T_3754; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_3755 = _T_2330 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4010 = _T_4009 | _T_3755; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_3756 = _T_2332 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4011 = _T_4010 | _T_3756; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_3757 = _T_2334 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4012 = _T_4011 | _T_3757; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_3758 = _T_2336 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4013 = _T_4012 | _T_3758; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_3759 = _T_2338 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4014 = _T_4013 | _T_3759; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_3760 = _T_2340 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4015 = _T_4014 | _T_3760; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_3761 = _T_2342 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4016 = _T_4015 | _T_3761; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_3762 = _T_2344 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4017 = _T_4016 | _T_3762; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_3763 = _T_2346 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4018 = _T_4017 | _T_3763; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_3764 = _T_2348 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4019 = _T_4018 | _T_3764; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_3765 = _T_2350 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4020 = _T_4019 | _T_3765; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_3766 = _T_2352 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4021 = _T_4020 | _T_3766; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_3767 = _T_2354 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4022 = _T_4021 | _T_3767; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_3768 = _T_2356 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4023 = _T_4022 | _T_3768; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_3769 = _T_2358 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4024 = _T_4023 | _T_3769; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_3770 = _T_2360 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4025 = _T_4024 | _T_3770; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_3771 = _T_2362 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4026 = _T_4025 | _T_3771; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_3772 = _T_2364 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4027 = _T_4026 | _T_3772; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_3773 = _T_2366 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4028 = _T_4027 | _T_3773; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_3774 = _T_2368 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4029 = _T_4028 | _T_3774; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_3775 = _T_2370 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4030 = _T_4029 | _T_3775; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_3776 = _T_2372 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4031 = _T_4030 | _T_3776; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_3777 = _T_2374 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4032 = _T_4031 | _T_3777; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_3778 = _T_2376 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4033 = _T_4032 | _T_3778; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_3779 = _T_2378 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4034 = _T_4033 | _T_3779; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_3780 = _T_2380 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4035 = _T_4034 | _T_3780; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_3781 = _T_2382 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4036 = _T_4035 | _T_3781; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_3782 = _T_2384 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4037 = _T_4036 | _T_3782; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_3783 = _T_2386 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4038 = _T_4037 | _T_3783; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_3784 = _T_2388 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4039 = _T_4038 | _T_3784; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_3785 = _T_2390 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4040 = _T_4039 | _T_3785; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_3786 = _T_2392 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4041 = _T_4040 | _T_3786; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_3787 = _T_2394 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4042 = _T_4041 | _T_3787; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_3788 = _T_2396 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4043 = _T_4042 | _T_3788; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_3789 = _T_2398 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4044 = _T_4043 | _T_3789; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_3790 = _T_2400 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4045 = _T_4044 | _T_3790; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_3791 = _T_2402 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4046 = _T_4045 | _T_3791; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_3792 = _T_2404 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4047 = _T_4046 | _T_3792; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_3793 = _T_2406 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4048 = _T_4047 | _T_3793; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_3794 = _T_2408 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4049 = _T_4048 | _T_3794; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_3795 = _T_2410 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4050 = _T_4049 | _T_3795; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_3796 = _T_2412 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4051 = _T_4050 | _T_3796; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_3797 = _T_2414 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4052 = _T_4051 | _T_3797; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_3798 = _T_2416 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4053 = _T_4052 | _T_3798; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_3799 = _T_2418 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4054 = _T_4053 | _T_3799; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_3800 = _T_2420 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4055 = _T_4054 | _T_3800; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_3801 = _T_2422 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4056 = _T_4055 | _T_3801; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_3802 = _T_2424 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4057 = _T_4056 | _T_3802; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_3803 = _T_2426 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4058 = _T_4057 | _T_3803; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_3804 = _T_2428 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4059 = _T_4058 | _T_3804; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_3805 = _T_2430 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4060 = _T_4059 | _T_3805; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_3806 = _T_2432 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4061 = _T_4060 | _T_3806; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_3807 = _T_2434 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4062 = _T_4061 | _T_3807; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_3808 = _T_2436 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4063 = _T_4062 | _T_3808; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_3809 = _T_2438 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4064 = _T_4063 | _T_3809; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_3810 = _T_2440 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4065 = _T_4064 | _T_3810; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_3811 = _T_2442 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4066 = _T_4065 | _T_3811; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_3812 = _T_2444 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4067 = _T_4066 | _T_3812; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_3813 = _T_2446 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4068 = _T_4067 | _T_3813; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_3814 = _T_2448 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4069 = _T_4068 | _T_3814; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_3815 = _T_2450 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4070 = _T_4069 | _T_3815; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_3816 = _T_2452 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4071 = _T_4070 | _T_3816; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_3817 = _T_2454 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4072 = _T_4071 | _T_3817; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_3818 = _T_2456 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4073 = _T_4072 | _T_3818; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_3819 = _T_2458 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4074 = _T_4073 | _T_3819; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_3820 = _T_2460 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4075 = _T_4074 | _T_3820; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_3821 = _T_2462 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4076 = _T_4075 | _T_3821; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_3822 = _T_2464 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4077 = _T_4076 | _T_3822; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_3823 = _T_2466 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4078 = _T_4077 | _T_3823; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_3824 = _T_2468 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4079 = _T_4078 | _T_3824; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_3825 = _T_2470 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4080 = _T_4079 | _T_3825; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_3826 = _T_2472 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4081 = _T_4080 | _T_3826; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_3827 = _T_2474 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4082 = _T_4081 | _T_3827; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_3828 = _T_2476 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4083 = _T_4082 | _T_3828; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_3829 = _T_2478 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4084 = _T_4083 | _T_3829; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_3830 = _T_2480 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4085 = _T_4084 | _T_3830; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_3831 = _T_2482 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4086 = _T_4085 | _T_3831; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_3832 = _T_2484 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4087 = _T_4086 | _T_3832; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_3833 = _T_2486 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4088 = _T_4087 | _T_3833; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_3834 = _T_2488 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4089 = _T_4088 | _T_3834; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_3835 = _T_2490 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4090 = _T_4089 | _T_3835; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_3836 = _T_2492 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4091 = _T_4090 | _T_3836; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_3837 = _T_2494 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4092 = _T_4091 | _T_3837; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_3838 = _T_2496 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4093 = _T_4092 | _T_3838; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_3839 = _T_2498 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4094 = _T_4093 | _T_3839; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_3840 = _T_2500 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4095 = _T_4094 | _T_3840; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_3841 = _T_2502 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4096 = _T_4095 | _T_3841; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_3842 = _T_2504 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4097 = _T_4096 | _T_3842; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_3843 = _T_2506 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4098 = _T_4097 | _T_3843; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_3844 = _T_2508 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4099 = _T_4098 | _T_3844; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_3845 = _T_2510 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4100 = _T_4099 | _T_3845; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_3846 = _T_2512 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4101 = _T_4100 | _T_3846; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_3847 = _T_2514 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4102 = _T_4101 | _T_3847; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_3848 = _T_2516 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4103 = _T_4102 | _T_3848; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_3849 = _T_2518 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4104 = _T_4103 | _T_3849; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_3850 = _T_2520 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4105 = _T_4104 | _T_3850; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_3851 = _T_2522 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4106 = _T_4105 | _T_3851; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_3852 = _T_2524 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4107 = _T_4106 | _T_3852; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_3853 = _T_2526 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4108 = _T_4107 | _T_3853; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_3854 = _T_2528 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4109 = _T_4108 | _T_3854; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_3855 = _T_2530 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4110 = _T_4109 | _T_3855; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_3856 = _T_2532 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4111 = _T_4110 | _T_3856; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_3857 = _T_2534 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4112 = _T_4111 | _T_3857; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_3858 = _T_2536 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4113 = _T_4112 | _T_3858; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_3859 = _T_2538 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4114 = _T_4113 | _T_3859; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_3860 = _T_2540 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4115 = _T_4114 | _T_3860; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_3861 = _T_2542 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4116 = _T_4115 | _T_3861; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_3862 = _T_2544 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4117 = _T_4116 | _T_3862; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_3863 = _T_2546 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4118 = _T_4117 | _T_3863; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_3864 = _T_2548 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4119 = _T_4118 | _T_3864; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_3865 = _T_2550 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4120 = _T_4119 | _T_3865; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_3866 = _T_2552 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4121 = _T_4120 | _T_3866; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_3867 = _T_2554 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4122 = _T_4121 | _T_3867; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_3868 = _T_2556 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4123 = _T_4122 | _T_3868; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_3869 = _T_2558 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4124 = _T_4123 | _T_3869; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_3870 = _T_2560 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4125 = _T_4124 | _T_3870; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_3871 = _T_2562 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4126 = _T_4125 | _T_3871; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_3872 = _T_2564 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4127 = _T_4126 | _T_3872; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_3873 = _T_2566 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4128 = _T_4127 | _T_3873; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_3874 = _T_2568 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4129 = _T_4128 | _T_3874; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_3875 = _T_2570 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4130 = _T_4129 | _T_3875; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_3876 = _T_2572 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4131 = _T_4130 | _T_3876; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_3877 = _T_2574 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4132 = _T_4131 | _T_3877; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_3878 = _T_2576 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4133 = _T_4132 | _T_3878; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_3879 = _T_2578 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4134 = _T_4133 | _T_3879; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_3880 = _T_2580 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4135 = _T_4134 | _T_3880; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_3881 = _T_2582 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4136 = _T_4135 | _T_3881; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_3882 = _T_2584 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4137 = _T_4136 | _T_3882; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_3883 = _T_2586 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4138 = _T_4137 | _T_3883; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_3884 = _T_2588 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4139 = _T_4138 | _T_3884; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_3885 = _T_2590 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4140 = _T_4139 | _T_3885; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_3886 = _T_2592 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4141 = _T_4140 | _T_3886; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_3887 = _T_2594 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4142 = _T_4141 | _T_3887; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_3888 = _T_2596 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4143 = _T_4142 | _T_3888; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_3889 = _T_2598 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4144 = _T_4143 | _T_3889; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_3890 = _T_2600 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4145 = _T_4144 | _T_3890; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_3891 = _T_2602 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4146 = _T_4145 | _T_3891; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_3892 = _T_2604 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4147 = _T_4146 | _T_3892; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_3893 = _T_2606 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4148 = _T_4147 | _T_3893; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_3894 = _T_2608 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4149 = _T_4148 | _T_3894; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_3895 = _T_2610 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4150 = _T_4149 | _T_3895; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_3896 = _T_2612 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4151 = _T_4150 | _T_3896; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_3897 = _T_2614 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4152 = _T_4151 | _T_3897; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_3898 = _T_2616 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4153 = _T_4152 | _T_3898; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_3899 = _T_2618 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4153 | _T_3899; // @[Mux.scala 27:72]
  wire  _T_54 = btb_bank0_rd_data_way1_f[21:17] == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 139:97]
  wire  _T_55 = btb_bank0_rd_data_way1_f[0] & _T_54; // @[el2_ifu_bp_ctl.scala 139:55]
  wire  _T_58 = _T_55 & _T_48; // @[el2_ifu_bp_ctl.scala 139:117]
  wire  _T_59 = _T_58 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 140:54]
  wire  tag_match_way1_f = _T_59 & _T; // @[el2_ifu_bp_ctl.scala 140:75]
  wire  _T_90 = btb_bank0_rd_data_way1_f[3] ^ btb_bank0_rd_data_way1_f[4]; // @[el2_ifu_bp_ctl.scala 152:91]
  wire  _T_91 = tag_match_way1_f & _T_90; // @[el2_ifu_bp_ctl.scala 152:56]
  wire  _T_95 = ~_T_90; // @[el2_ifu_bp_ctl.scala 153:58]
  wire  _T_96 = tag_match_way1_f & _T_95; // @[el2_ifu_bp_ctl.scala 153:56]
  wire [1:0] tag_match_way1_expanded_f = {_T_91,_T_96}; // @[Cat.scala 29:58]
  wire [21:0] _T_127 = tag_match_way1_expanded_f[1] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0o_rd_data_f = _T_126 | _T_127; // @[Mux.scala 27:72]
  wire [21:0] _T_145 = _T_143 ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4156 = btb_rd_addr_p1_f == 8'h0; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4668 = _T_4156 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4158 = btb_rd_addr_p1_f == 8'h1; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4669 = _T_4158 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4924 = _T_4668 | _T_4669; // @[Mux.scala 27:72]
  wire  _T_4160 = btb_rd_addr_p1_f == 8'h2; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4670 = _T_4160 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4925 = _T_4924 | _T_4670; // @[Mux.scala 27:72]
  wire  _T_4162 = btb_rd_addr_p1_f == 8'h3; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4671 = _T_4162 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4926 = _T_4925 | _T_4671; // @[Mux.scala 27:72]
  wire  _T_4164 = btb_rd_addr_p1_f == 8'h4; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4672 = _T_4164 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4927 = _T_4926 | _T_4672; // @[Mux.scala 27:72]
  wire  _T_4166 = btb_rd_addr_p1_f == 8'h5; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4673 = _T_4166 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4928 = _T_4927 | _T_4673; // @[Mux.scala 27:72]
  wire  _T_4168 = btb_rd_addr_p1_f == 8'h6; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4674 = _T_4168 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4929 = _T_4928 | _T_4674; // @[Mux.scala 27:72]
  wire  _T_4170 = btb_rd_addr_p1_f == 8'h7; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4675 = _T_4170 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4930 = _T_4929 | _T_4675; // @[Mux.scala 27:72]
  wire  _T_4172 = btb_rd_addr_p1_f == 8'h8; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4676 = _T_4172 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4931 = _T_4930 | _T_4676; // @[Mux.scala 27:72]
  wire  _T_4174 = btb_rd_addr_p1_f == 8'h9; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4677 = _T_4174 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4932 = _T_4931 | _T_4677; // @[Mux.scala 27:72]
  wire  _T_4176 = btb_rd_addr_p1_f == 8'ha; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4678 = _T_4176 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4933 = _T_4932 | _T_4678; // @[Mux.scala 27:72]
  wire  _T_4178 = btb_rd_addr_p1_f == 8'hb; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4679 = _T_4178 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4934 = _T_4933 | _T_4679; // @[Mux.scala 27:72]
  wire  _T_4180 = btb_rd_addr_p1_f == 8'hc; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4680 = _T_4180 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4935 = _T_4934 | _T_4680; // @[Mux.scala 27:72]
  wire  _T_4182 = btb_rd_addr_p1_f == 8'hd; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4681 = _T_4182 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4936 = _T_4935 | _T_4681; // @[Mux.scala 27:72]
  wire  _T_4184 = btb_rd_addr_p1_f == 8'he; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4682 = _T_4184 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4937 = _T_4936 | _T_4682; // @[Mux.scala 27:72]
  wire  _T_4186 = btb_rd_addr_p1_f == 8'hf; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4683 = _T_4186 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4938 = _T_4937 | _T_4683; // @[Mux.scala 27:72]
  wire  _T_4188 = btb_rd_addr_p1_f == 8'h10; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4684 = _T_4188 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4939 = _T_4938 | _T_4684; // @[Mux.scala 27:72]
  wire  _T_4190 = btb_rd_addr_p1_f == 8'h11; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4685 = _T_4190 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4940 = _T_4939 | _T_4685; // @[Mux.scala 27:72]
  wire  _T_4192 = btb_rd_addr_p1_f == 8'h12; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4686 = _T_4192 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4941 = _T_4940 | _T_4686; // @[Mux.scala 27:72]
  wire  _T_4194 = btb_rd_addr_p1_f == 8'h13; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4687 = _T_4194 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4942 = _T_4941 | _T_4687; // @[Mux.scala 27:72]
  wire  _T_4196 = btb_rd_addr_p1_f == 8'h14; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4688 = _T_4196 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4943 = _T_4942 | _T_4688; // @[Mux.scala 27:72]
  wire  _T_4198 = btb_rd_addr_p1_f == 8'h15; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4689 = _T_4198 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4944 = _T_4943 | _T_4689; // @[Mux.scala 27:72]
  wire  _T_4200 = btb_rd_addr_p1_f == 8'h16; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4690 = _T_4200 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4945 = _T_4944 | _T_4690; // @[Mux.scala 27:72]
  wire  _T_4202 = btb_rd_addr_p1_f == 8'h17; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4691 = _T_4202 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4946 = _T_4945 | _T_4691; // @[Mux.scala 27:72]
  wire  _T_4204 = btb_rd_addr_p1_f == 8'h18; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4692 = _T_4204 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4947 = _T_4946 | _T_4692; // @[Mux.scala 27:72]
  wire  _T_4206 = btb_rd_addr_p1_f == 8'h19; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4693 = _T_4206 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4948 = _T_4947 | _T_4693; // @[Mux.scala 27:72]
  wire  _T_4208 = btb_rd_addr_p1_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4694 = _T_4208 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4949 = _T_4948 | _T_4694; // @[Mux.scala 27:72]
  wire  _T_4210 = btb_rd_addr_p1_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4695 = _T_4210 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4950 = _T_4949 | _T_4695; // @[Mux.scala 27:72]
  wire  _T_4212 = btb_rd_addr_p1_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4696 = _T_4212 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4951 = _T_4950 | _T_4696; // @[Mux.scala 27:72]
  wire  _T_4214 = btb_rd_addr_p1_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4697 = _T_4214 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4952 = _T_4951 | _T_4697; // @[Mux.scala 27:72]
  wire  _T_4216 = btb_rd_addr_p1_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4698 = _T_4216 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4953 = _T_4952 | _T_4698; // @[Mux.scala 27:72]
  wire  _T_4218 = btb_rd_addr_p1_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4699 = _T_4218 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4954 = _T_4953 | _T_4699; // @[Mux.scala 27:72]
  wire  _T_4220 = btb_rd_addr_p1_f == 8'h20; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4700 = _T_4220 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4955 = _T_4954 | _T_4700; // @[Mux.scala 27:72]
  wire  _T_4222 = btb_rd_addr_p1_f == 8'h21; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4701 = _T_4222 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4956 = _T_4955 | _T_4701; // @[Mux.scala 27:72]
  wire  _T_4224 = btb_rd_addr_p1_f == 8'h22; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4702 = _T_4224 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4957 = _T_4956 | _T_4702; // @[Mux.scala 27:72]
  wire  _T_4226 = btb_rd_addr_p1_f == 8'h23; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4703 = _T_4226 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4958 = _T_4957 | _T_4703; // @[Mux.scala 27:72]
  wire  _T_4228 = btb_rd_addr_p1_f == 8'h24; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4704 = _T_4228 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4959 = _T_4958 | _T_4704; // @[Mux.scala 27:72]
  wire  _T_4230 = btb_rd_addr_p1_f == 8'h25; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4705 = _T_4230 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4960 = _T_4959 | _T_4705; // @[Mux.scala 27:72]
  wire  _T_4232 = btb_rd_addr_p1_f == 8'h26; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4706 = _T_4232 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4961 = _T_4960 | _T_4706; // @[Mux.scala 27:72]
  wire  _T_4234 = btb_rd_addr_p1_f == 8'h27; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4707 = _T_4234 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4962 = _T_4961 | _T_4707; // @[Mux.scala 27:72]
  wire  _T_4236 = btb_rd_addr_p1_f == 8'h28; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4708 = _T_4236 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4963 = _T_4962 | _T_4708; // @[Mux.scala 27:72]
  wire  _T_4238 = btb_rd_addr_p1_f == 8'h29; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4709 = _T_4238 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4964 = _T_4963 | _T_4709; // @[Mux.scala 27:72]
  wire  _T_4240 = btb_rd_addr_p1_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4710 = _T_4240 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4965 = _T_4964 | _T_4710; // @[Mux.scala 27:72]
  wire  _T_4242 = btb_rd_addr_p1_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4711 = _T_4242 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4966 = _T_4965 | _T_4711; // @[Mux.scala 27:72]
  wire  _T_4244 = btb_rd_addr_p1_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4712 = _T_4244 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4967 = _T_4966 | _T_4712; // @[Mux.scala 27:72]
  wire  _T_4246 = btb_rd_addr_p1_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4713 = _T_4246 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4968 = _T_4967 | _T_4713; // @[Mux.scala 27:72]
  wire  _T_4248 = btb_rd_addr_p1_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4714 = _T_4248 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4969 = _T_4968 | _T_4714; // @[Mux.scala 27:72]
  wire  _T_4250 = btb_rd_addr_p1_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4715 = _T_4250 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4970 = _T_4969 | _T_4715; // @[Mux.scala 27:72]
  wire  _T_4252 = btb_rd_addr_p1_f == 8'h30; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4716 = _T_4252 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4971 = _T_4970 | _T_4716; // @[Mux.scala 27:72]
  wire  _T_4254 = btb_rd_addr_p1_f == 8'h31; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4717 = _T_4254 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4972 = _T_4971 | _T_4717; // @[Mux.scala 27:72]
  wire  _T_4256 = btb_rd_addr_p1_f == 8'h32; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4718 = _T_4256 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4973 = _T_4972 | _T_4718; // @[Mux.scala 27:72]
  wire  _T_4258 = btb_rd_addr_p1_f == 8'h33; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4719 = _T_4258 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4974 = _T_4973 | _T_4719; // @[Mux.scala 27:72]
  wire  _T_4260 = btb_rd_addr_p1_f == 8'h34; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4720 = _T_4260 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4975 = _T_4974 | _T_4720; // @[Mux.scala 27:72]
  wire  _T_4262 = btb_rd_addr_p1_f == 8'h35; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4721 = _T_4262 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4976 = _T_4975 | _T_4721; // @[Mux.scala 27:72]
  wire  _T_4264 = btb_rd_addr_p1_f == 8'h36; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4722 = _T_4264 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4977 = _T_4976 | _T_4722; // @[Mux.scala 27:72]
  wire  _T_4266 = btb_rd_addr_p1_f == 8'h37; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4723 = _T_4266 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4978 = _T_4977 | _T_4723; // @[Mux.scala 27:72]
  wire  _T_4268 = btb_rd_addr_p1_f == 8'h38; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4724 = _T_4268 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4979 = _T_4978 | _T_4724; // @[Mux.scala 27:72]
  wire  _T_4270 = btb_rd_addr_p1_f == 8'h39; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4725 = _T_4270 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4980 = _T_4979 | _T_4725; // @[Mux.scala 27:72]
  wire  _T_4272 = btb_rd_addr_p1_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4726 = _T_4272 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4981 = _T_4980 | _T_4726; // @[Mux.scala 27:72]
  wire  _T_4274 = btb_rd_addr_p1_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4727 = _T_4274 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4982 = _T_4981 | _T_4727; // @[Mux.scala 27:72]
  wire  _T_4276 = btb_rd_addr_p1_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4728 = _T_4276 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4983 = _T_4982 | _T_4728; // @[Mux.scala 27:72]
  wire  _T_4278 = btb_rd_addr_p1_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4729 = _T_4278 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4984 = _T_4983 | _T_4729; // @[Mux.scala 27:72]
  wire  _T_4280 = btb_rd_addr_p1_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4730 = _T_4280 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4985 = _T_4984 | _T_4730; // @[Mux.scala 27:72]
  wire  _T_4282 = btb_rd_addr_p1_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4731 = _T_4282 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4986 = _T_4985 | _T_4731; // @[Mux.scala 27:72]
  wire  _T_4284 = btb_rd_addr_p1_f == 8'h40; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4732 = _T_4284 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4987 = _T_4986 | _T_4732; // @[Mux.scala 27:72]
  wire  _T_4286 = btb_rd_addr_p1_f == 8'h41; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4733 = _T_4286 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4988 = _T_4987 | _T_4733; // @[Mux.scala 27:72]
  wire  _T_4288 = btb_rd_addr_p1_f == 8'h42; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4734 = _T_4288 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4989 = _T_4988 | _T_4734; // @[Mux.scala 27:72]
  wire  _T_4290 = btb_rd_addr_p1_f == 8'h43; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4735 = _T_4290 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4990 = _T_4989 | _T_4735; // @[Mux.scala 27:72]
  wire  _T_4292 = btb_rd_addr_p1_f == 8'h44; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4736 = _T_4292 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4991 = _T_4990 | _T_4736; // @[Mux.scala 27:72]
  wire  _T_4294 = btb_rd_addr_p1_f == 8'h45; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4737 = _T_4294 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4992 = _T_4991 | _T_4737; // @[Mux.scala 27:72]
  wire  _T_4296 = btb_rd_addr_p1_f == 8'h46; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4738 = _T_4296 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4993 = _T_4992 | _T_4738; // @[Mux.scala 27:72]
  wire  _T_4298 = btb_rd_addr_p1_f == 8'h47; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4739 = _T_4298 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4994 = _T_4993 | _T_4739; // @[Mux.scala 27:72]
  wire  _T_4300 = btb_rd_addr_p1_f == 8'h48; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4740 = _T_4300 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4995 = _T_4994 | _T_4740; // @[Mux.scala 27:72]
  wire  _T_4302 = btb_rd_addr_p1_f == 8'h49; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4741 = _T_4302 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4996 = _T_4995 | _T_4741; // @[Mux.scala 27:72]
  wire  _T_4304 = btb_rd_addr_p1_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4742 = _T_4304 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4997 = _T_4996 | _T_4742; // @[Mux.scala 27:72]
  wire  _T_4306 = btb_rd_addr_p1_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4743 = _T_4306 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4998 = _T_4997 | _T_4743; // @[Mux.scala 27:72]
  wire  _T_4308 = btb_rd_addr_p1_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4744 = _T_4308 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4999 = _T_4998 | _T_4744; // @[Mux.scala 27:72]
  wire  _T_4310 = btb_rd_addr_p1_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4745 = _T_4310 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5000 = _T_4999 | _T_4745; // @[Mux.scala 27:72]
  wire  _T_4312 = btb_rd_addr_p1_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4746 = _T_4312 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5001 = _T_5000 | _T_4746; // @[Mux.scala 27:72]
  wire  _T_4314 = btb_rd_addr_p1_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4747 = _T_4314 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5002 = _T_5001 | _T_4747; // @[Mux.scala 27:72]
  wire  _T_4316 = btb_rd_addr_p1_f == 8'h50; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4748 = _T_4316 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5003 = _T_5002 | _T_4748; // @[Mux.scala 27:72]
  wire  _T_4318 = btb_rd_addr_p1_f == 8'h51; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4749 = _T_4318 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5004 = _T_5003 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4320 = btb_rd_addr_p1_f == 8'h52; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4750 = _T_4320 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5005 = _T_5004 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4322 = btb_rd_addr_p1_f == 8'h53; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4751 = _T_4322 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5006 = _T_5005 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4324 = btb_rd_addr_p1_f == 8'h54; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4752 = _T_4324 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5007 = _T_5006 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4326 = btb_rd_addr_p1_f == 8'h55; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4753 = _T_4326 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5008 = _T_5007 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4328 = btb_rd_addr_p1_f == 8'h56; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4754 = _T_4328 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5009 = _T_5008 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4330 = btb_rd_addr_p1_f == 8'h57; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4755 = _T_4330 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5010 = _T_5009 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4332 = btb_rd_addr_p1_f == 8'h58; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4756 = _T_4332 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5011 = _T_5010 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4334 = btb_rd_addr_p1_f == 8'h59; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4757 = _T_4334 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5012 = _T_5011 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4336 = btb_rd_addr_p1_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4758 = _T_4336 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5013 = _T_5012 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4338 = btb_rd_addr_p1_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4759 = _T_4338 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5014 = _T_5013 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4340 = btb_rd_addr_p1_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4760 = _T_4340 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5015 = _T_5014 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4342 = btb_rd_addr_p1_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4761 = _T_4342 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5016 = _T_5015 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4344 = btb_rd_addr_p1_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4762 = _T_4344 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5017 = _T_5016 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4346 = btb_rd_addr_p1_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4763 = _T_4346 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5018 = _T_5017 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4348 = btb_rd_addr_p1_f == 8'h60; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4764 = _T_4348 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5019 = _T_5018 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4350 = btb_rd_addr_p1_f == 8'h61; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4765 = _T_4350 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5020 = _T_5019 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4352 = btb_rd_addr_p1_f == 8'h62; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4766 = _T_4352 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5021 = _T_5020 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4354 = btb_rd_addr_p1_f == 8'h63; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4767 = _T_4354 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5022 = _T_5021 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4356 = btb_rd_addr_p1_f == 8'h64; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4768 = _T_4356 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5023 = _T_5022 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4358 = btb_rd_addr_p1_f == 8'h65; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4769 = _T_4358 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5024 = _T_5023 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4360 = btb_rd_addr_p1_f == 8'h66; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4770 = _T_4360 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5025 = _T_5024 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4362 = btb_rd_addr_p1_f == 8'h67; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4771 = _T_4362 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5026 = _T_5025 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4364 = btb_rd_addr_p1_f == 8'h68; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4772 = _T_4364 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5027 = _T_5026 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4366 = btb_rd_addr_p1_f == 8'h69; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4773 = _T_4366 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5028 = _T_5027 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4368 = btb_rd_addr_p1_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4774 = _T_4368 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5029 = _T_5028 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4370 = btb_rd_addr_p1_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4775 = _T_4370 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5030 = _T_5029 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4372 = btb_rd_addr_p1_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4776 = _T_4372 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5031 = _T_5030 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4374 = btb_rd_addr_p1_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4777 = _T_4374 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5032 = _T_5031 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4376 = btb_rd_addr_p1_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4778 = _T_4376 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5033 = _T_5032 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4378 = btb_rd_addr_p1_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4779 = _T_4378 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5034 = _T_5033 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4380 = btb_rd_addr_p1_f == 8'h70; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4780 = _T_4380 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5035 = _T_5034 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4382 = btb_rd_addr_p1_f == 8'h71; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4781 = _T_4382 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5036 = _T_5035 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4384 = btb_rd_addr_p1_f == 8'h72; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4782 = _T_4384 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5037 = _T_5036 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4386 = btb_rd_addr_p1_f == 8'h73; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4783 = _T_4386 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5038 = _T_5037 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4388 = btb_rd_addr_p1_f == 8'h74; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4784 = _T_4388 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5039 = _T_5038 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4390 = btb_rd_addr_p1_f == 8'h75; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4785 = _T_4390 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5040 = _T_5039 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4392 = btb_rd_addr_p1_f == 8'h76; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4786 = _T_4392 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5041 = _T_5040 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4394 = btb_rd_addr_p1_f == 8'h77; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4787 = _T_4394 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5042 = _T_5041 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4396 = btb_rd_addr_p1_f == 8'h78; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4788 = _T_4396 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5043 = _T_5042 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4398 = btb_rd_addr_p1_f == 8'h79; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4789 = _T_4398 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5044 = _T_5043 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4400 = btb_rd_addr_p1_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4790 = _T_4400 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5045 = _T_5044 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4402 = btb_rd_addr_p1_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4791 = _T_4402 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5046 = _T_5045 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4404 = btb_rd_addr_p1_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4792 = _T_4404 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5047 = _T_5046 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4406 = btb_rd_addr_p1_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4793 = _T_4406 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5048 = _T_5047 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4408 = btb_rd_addr_p1_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4794 = _T_4408 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5049 = _T_5048 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4410 = btb_rd_addr_p1_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4795 = _T_4410 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5050 = _T_5049 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4412 = btb_rd_addr_p1_f == 8'h80; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4796 = _T_4412 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5051 = _T_5050 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4414 = btb_rd_addr_p1_f == 8'h81; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4797 = _T_4414 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5052 = _T_5051 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4416 = btb_rd_addr_p1_f == 8'h82; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4798 = _T_4416 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5053 = _T_5052 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4418 = btb_rd_addr_p1_f == 8'h83; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4799 = _T_4418 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5054 = _T_5053 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4420 = btb_rd_addr_p1_f == 8'h84; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4800 = _T_4420 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5055 = _T_5054 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4422 = btb_rd_addr_p1_f == 8'h85; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4801 = _T_4422 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5056 = _T_5055 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4424 = btb_rd_addr_p1_f == 8'h86; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4802 = _T_4424 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5057 = _T_5056 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4426 = btb_rd_addr_p1_f == 8'h87; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4803 = _T_4426 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5058 = _T_5057 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4428 = btb_rd_addr_p1_f == 8'h88; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4804 = _T_4428 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5059 = _T_5058 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4430 = btb_rd_addr_p1_f == 8'h89; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4805 = _T_4430 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5060 = _T_5059 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4432 = btb_rd_addr_p1_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4806 = _T_4432 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5061 = _T_5060 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4434 = btb_rd_addr_p1_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4807 = _T_4434 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5062 = _T_5061 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4436 = btb_rd_addr_p1_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4808 = _T_4436 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5063 = _T_5062 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4438 = btb_rd_addr_p1_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4809 = _T_4438 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5064 = _T_5063 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4440 = btb_rd_addr_p1_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4810 = _T_4440 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5065 = _T_5064 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4442 = btb_rd_addr_p1_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4811 = _T_4442 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5066 = _T_5065 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4444 = btb_rd_addr_p1_f == 8'h90; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4812 = _T_4444 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5067 = _T_5066 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4446 = btb_rd_addr_p1_f == 8'h91; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4813 = _T_4446 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5068 = _T_5067 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4448 = btb_rd_addr_p1_f == 8'h92; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4814 = _T_4448 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5069 = _T_5068 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4450 = btb_rd_addr_p1_f == 8'h93; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4815 = _T_4450 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5070 = _T_5069 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4452 = btb_rd_addr_p1_f == 8'h94; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4816 = _T_4452 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5071 = _T_5070 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4454 = btb_rd_addr_p1_f == 8'h95; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4817 = _T_4454 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5072 = _T_5071 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4456 = btb_rd_addr_p1_f == 8'h96; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4818 = _T_4456 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5073 = _T_5072 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4458 = btb_rd_addr_p1_f == 8'h97; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4819 = _T_4458 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5074 = _T_5073 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4460 = btb_rd_addr_p1_f == 8'h98; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4820 = _T_4460 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5075 = _T_5074 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4462 = btb_rd_addr_p1_f == 8'h99; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4821 = _T_4462 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5076 = _T_5075 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4464 = btb_rd_addr_p1_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4822 = _T_4464 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5077 = _T_5076 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4466 = btb_rd_addr_p1_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4823 = _T_4466 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5078 = _T_5077 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4468 = btb_rd_addr_p1_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4824 = _T_4468 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5079 = _T_5078 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4470 = btb_rd_addr_p1_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4825 = _T_4470 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5080 = _T_5079 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4472 = btb_rd_addr_p1_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4826 = _T_4472 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5081 = _T_5080 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4474 = btb_rd_addr_p1_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4827 = _T_4474 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5082 = _T_5081 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4476 = btb_rd_addr_p1_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4828 = _T_4476 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5083 = _T_5082 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4478 = btb_rd_addr_p1_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4829 = _T_4478 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5084 = _T_5083 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4480 = btb_rd_addr_p1_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4830 = _T_4480 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5085 = _T_5084 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4482 = btb_rd_addr_p1_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4831 = _T_4482 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5086 = _T_5085 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4484 = btb_rd_addr_p1_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4832 = _T_4484 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5087 = _T_5086 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4486 = btb_rd_addr_p1_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4833 = _T_4486 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5088 = _T_5087 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4488 = btb_rd_addr_p1_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4834 = _T_4488 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5089 = _T_5088 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4490 = btb_rd_addr_p1_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4835 = _T_4490 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5090 = _T_5089 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4492 = btb_rd_addr_p1_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4836 = _T_4492 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5091 = _T_5090 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4494 = btb_rd_addr_p1_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4837 = _T_4494 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5092 = _T_5091 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4496 = btb_rd_addr_p1_f == 8'haa; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4838 = _T_4496 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5093 = _T_5092 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4498 = btb_rd_addr_p1_f == 8'hab; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4839 = _T_4498 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5094 = _T_5093 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4500 = btb_rd_addr_p1_f == 8'hac; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4840 = _T_4500 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5095 = _T_5094 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4502 = btb_rd_addr_p1_f == 8'had; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4841 = _T_4502 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5096 = _T_5095 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4504 = btb_rd_addr_p1_f == 8'hae; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4842 = _T_4504 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5097 = _T_5096 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4506 = btb_rd_addr_p1_f == 8'haf; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4843 = _T_4506 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5098 = _T_5097 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4508 = btb_rd_addr_p1_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4844 = _T_4508 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5099 = _T_5098 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4510 = btb_rd_addr_p1_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4845 = _T_4510 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5100 = _T_5099 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4512 = btb_rd_addr_p1_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4846 = _T_4512 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5101 = _T_5100 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4514 = btb_rd_addr_p1_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4847 = _T_4514 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5102 = _T_5101 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4516 = btb_rd_addr_p1_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4848 = _T_4516 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5103 = _T_5102 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4518 = btb_rd_addr_p1_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4849 = _T_4518 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5104 = _T_5103 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4520 = btb_rd_addr_p1_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4850 = _T_4520 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5105 = _T_5104 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4522 = btb_rd_addr_p1_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4851 = _T_4522 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5106 = _T_5105 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4524 = btb_rd_addr_p1_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4852 = _T_4524 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5107 = _T_5106 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4526 = btb_rd_addr_p1_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4853 = _T_4526 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5108 = _T_5107 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4528 = btb_rd_addr_p1_f == 8'hba; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4854 = _T_4528 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5109 = _T_5108 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4530 = btb_rd_addr_p1_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4855 = _T_4530 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5110 = _T_5109 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4532 = btb_rd_addr_p1_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4856 = _T_4532 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5111 = _T_5110 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4534 = btb_rd_addr_p1_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4857 = _T_4534 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5112 = _T_5111 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4536 = btb_rd_addr_p1_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4858 = _T_4536 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5113 = _T_5112 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4538 = btb_rd_addr_p1_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4859 = _T_4538 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5114 = _T_5113 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4540 = btb_rd_addr_p1_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4860 = _T_4540 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5115 = _T_5114 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4542 = btb_rd_addr_p1_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4861 = _T_4542 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5116 = _T_5115 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4544 = btb_rd_addr_p1_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4862 = _T_4544 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5117 = _T_5116 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4546 = btb_rd_addr_p1_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4863 = _T_4546 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5118 = _T_5117 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4548 = btb_rd_addr_p1_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4864 = _T_4548 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5119 = _T_5118 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4550 = btb_rd_addr_p1_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4865 = _T_4550 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5120 = _T_5119 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4552 = btb_rd_addr_p1_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4866 = _T_4552 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5121 = _T_5120 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4554 = btb_rd_addr_p1_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4867 = _T_4554 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5122 = _T_5121 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4556 = btb_rd_addr_p1_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4868 = _T_4556 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5123 = _T_5122 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4558 = btb_rd_addr_p1_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4869 = _T_4558 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5124 = _T_5123 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4560 = btb_rd_addr_p1_f == 8'hca; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4870 = _T_4560 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5125 = _T_5124 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4562 = btb_rd_addr_p1_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4871 = _T_4562 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5126 = _T_5125 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4564 = btb_rd_addr_p1_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4872 = _T_4564 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5127 = _T_5126 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4566 = btb_rd_addr_p1_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4873 = _T_4566 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5128 = _T_5127 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4568 = btb_rd_addr_p1_f == 8'hce; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4874 = _T_4568 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5129 = _T_5128 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4570 = btb_rd_addr_p1_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4875 = _T_4570 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5130 = _T_5129 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4572 = btb_rd_addr_p1_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4876 = _T_4572 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5131 = _T_5130 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4574 = btb_rd_addr_p1_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4877 = _T_4574 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5132 = _T_5131 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4576 = btb_rd_addr_p1_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4878 = _T_4576 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5133 = _T_5132 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4578 = btb_rd_addr_p1_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4879 = _T_4578 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5134 = _T_5133 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4580 = btb_rd_addr_p1_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4880 = _T_4580 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5135 = _T_5134 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4582 = btb_rd_addr_p1_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4881 = _T_4582 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5136 = _T_5135 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4584 = btb_rd_addr_p1_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4882 = _T_4584 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5137 = _T_5136 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4586 = btb_rd_addr_p1_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4883 = _T_4586 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5138 = _T_5137 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4588 = btb_rd_addr_p1_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4884 = _T_4588 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5139 = _T_5138 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4590 = btb_rd_addr_p1_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4885 = _T_4590 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5140 = _T_5139 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4592 = btb_rd_addr_p1_f == 8'hda; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4886 = _T_4592 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5141 = _T_5140 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4594 = btb_rd_addr_p1_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4887 = _T_4594 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5142 = _T_5141 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4596 = btb_rd_addr_p1_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4888 = _T_4596 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5143 = _T_5142 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4598 = btb_rd_addr_p1_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4889 = _T_4598 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5144 = _T_5143 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4600 = btb_rd_addr_p1_f == 8'hde; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4890 = _T_4600 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5145 = _T_5144 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4602 = btb_rd_addr_p1_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4891 = _T_4602 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5146 = _T_5145 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4604 = btb_rd_addr_p1_f == 8'he0; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4892 = _T_4604 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5147 = _T_5146 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4606 = btb_rd_addr_p1_f == 8'he1; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4893 = _T_4606 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5148 = _T_5147 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4608 = btb_rd_addr_p1_f == 8'he2; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4894 = _T_4608 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5149 = _T_5148 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4610 = btb_rd_addr_p1_f == 8'he3; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4895 = _T_4610 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5150 = _T_5149 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4612 = btb_rd_addr_p1_f == 8'he4; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4896 = _T_4612 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5151 = _T_5150 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4614 = btb_rd_addr_p1_f == 8'he5; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4897 = _T_4614 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5152 = _T_5151 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4616 = btb_rd_addr_p1_f == 8'he6; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4898 = _T_4616 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5153 = _T_5152 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4618 = btb_rd_addr_p1_f == 8'he7; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4899 = _T_4618 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5154 = _T_5153 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4620 = btb_rd_addr_p1_f == 8'he8; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4900 = _T_4620 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5155 = _T_5154 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4622 = btb_rd_addr_p1_f == 8'he9; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4901 = _T_4622 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5156 = _T_5155 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4624 = btb_rd_addr_p1_f == 8'hea; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4902 = _T_4624 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5157 = _T_5156 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4626 = btb_rd_addr_p1_f == 8'heb; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4903 = _T_4626 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5158 = _T_5157 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4628 = btb_rd_addr_p1_f == 8'hec; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4904 = _T_4628 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5159 = _T_5158 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4630 = btb_rd_addr_p1_f == 8'hed; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4905 = _T_4630 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5160 = _T_5159 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4632 = btb_rd_addr_p1_f == 8'hee; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4906 = _T_4632 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5161 = _T_5160 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4634 = btb_rd_addr_p1_f == 8'hef; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4907 = _T_4634 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5162 = _T_5161 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4636 = btb_rd_addr_p1_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4908 = _T_4636 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5163 = _T_5162 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4638 = btb_rd_addr_p1_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4909 = _T_4638 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5164 = _T_5163 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4640 = btb_rd_addr_p1_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4910 = _T_4640 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5165 = _T_5164 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4642 = btb_rd_addr_p1_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4911 = _T_4642 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5166 = _T_5165 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4644 = btb_rd_addr_p1_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4912 = _T_4644 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5167 = _T_5166 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4646 = btb_rd_addr_p1_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4913 = _T_4646 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5168 = _T_5167 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4648 = btb_rd_addr_p1_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4914 = _T_4648 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5169 = _T_5168 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4650 = btb_rd_addr_p1_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4915 = _T_4650 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5170 = _T_5169 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4652 = btb_rd_addr_p1_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4916 = _T_4652 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5171 = _T_5170 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4654 = btb_rd_addr_p1_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4917 = _T_4654 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5172 = _T_5171 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4656 = btb_rd_addr_p1_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4918 = _T_4656 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5173 = _T_5172 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4658 = btb_rd_addr_p1_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4919 = _T_4658 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5174 = _T_5173 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4660 = btb_rd_addr_p1_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4920 = _T_4660 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5175 = _T_5174 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4662 = btb_rd_addr_p1_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4921 = _T_4662 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5176 = _T_5175 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4664 = btb_rd_addr_p1_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4922 = _T_4664 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5177 = _T_5176 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4666 = btb_rd_addr_p1_f == 8'hff; // @[el2_ifu_bp_ctl.scala 372:83]
  wire [21:0] _T_4923 = _T_4666 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5177 | _T_4923; // @[Mux.scala 27:72]
  wire [4:0] _T_31 = _T_8[13:9] ^ _T_8[18:14]; // @[el2_lib.scala 174:111]
  wire [4:0] fetch_rd_tag_p1_f = _T_31 ^ _T_8[23:19]; // @[el2_lib.scala 174:111]
  wire  _T_63 = btb_bank0_rd_data_way0_p1_f[21:17] == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 142:106]
  wire  _T_64 = btb_bank0_rd_data_way0_p1_f[0] & _T_63; // @[el2_ifu_bp_ctl.scala 142:61]
  wire  _T_67 = _T_64 & _T_48; // @[el2_ifu_bp_ctl.scala 142:129]
  wire  _T_68 = _T_67 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 143:56]
  wire  tag_match_way0_p1_f = _T_68 & _T; // @[el2_ifu_bp_ctl.scala 143:77]
  wire  _T_99 = btb_bank0_rd_data_way0_p1_f[3] ^ btb_bank0_rd_data_way0_p1_f[4]; // @[el2_ifu_bp_ctl.scala 156:100]
  wire  _T_100 = tag_match_way0_p1_f & _T_99; // @[el2_ifu_bp_ctl.scala 156:62]
  wire  _T_104 = ~_T_99; // @[el2_ifu_bp_ctl.scala 157:64]
  wire  _T_105 = tag_match_way0_p1_f & _T_104; // @[el2_ifu_bp_ctl.scala 157:62]
  wire [1:0] tag_match_way0_expanded_p1_f = {_T_100,_T_105}; // @[Cat.scala 29:58]
  wire [21:0] _T_133 = tag_match_way0_expanded_p1_f[0] ? btb_bank0_rd_data_way0_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5692 = _T_4156 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5693 = _T_4158 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5948 = _T_5692 | _T_5693; // @[Mux.scala 27:72]
  wire [21:0] _T_5694 = _T_4160 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5949 = _T_5948 | _T_5694; // @[Mux.scala 27:72]
  wire [21:0] _T_5695 = _T_4162 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5950 = _T_5949 | _T_5695; // @[Mux.scala 27:72]
  wire [21:0] _T_5696 = _T_4164 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5951 = _T_5950 | _T_5696; // @[Mux.scala 27:72]
  wire [21:0] _T_5697 = _T_4166 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5952 = _T_5951 | _T_5697; // @[Mux.scala 27:72]
  wire [21:0] _T_5698 = _T_4168 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5953 = _T_5952 | _T_5698; // @[Mux.scala 27:72]
  wire [21:0] _T_5699 = _T_4170 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5954 = _T_5953 | _T_5699; // @[Mux.scala 27:72]
  wire [21:0] _T_5700 = _T_4172 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5955 = _T_5954 | _T_5700; // @[Mux.scala 27:72]
  wire [21:0] _T_5701 = _T_4174 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5956 = _T_5955 | _T_5701; // @[Mux.scala 27:72]
  wire [21:0] _T_5702 = _T_4176 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5957 = _T_5956 | _T_5702; // @[Mux.scala 27:72]
  wire [21:0] _T_5703 = _T_4178 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5958 = _T_5957 | _T_5703; // @[Mux.scala 27:72]
  wire [21:0] _T_5704 = _T_4180 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5959 = _T_5958 | _T_5704; // @[Mux.scala 27:72]
  wire [21:0] _T_5705 = _T_4182 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5960 = _T_5959 | _T_5705; // @[Mux.scala 27:72]
  wire [21:0] _T_5706 = _T_4184 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5961 = _T_5960 | _T_5706; // @[Mux.scala 27:72]
  wire [21:0] _T_5707 = _T_4186 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5962 = _T_5961 | _T_5707; // @[Mux.scala 27:72]
  wire [21:0] _T_5708 = _T_4188 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5963 = _T_5962 | _T_5708; // @[Mux.scala 27:72]
  wire [21:0] _T_5709 = _T_4190 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5964 = _T_5963 | _T_5709; // @[Mux.scala 27:72]
  wire [21:0] _T_5710 = _T_4192 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5965 = _T_5964 | _T_5710; // @[Mux.scala 27:72]
  wire [21:0] _T_5711 = _T_4194 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5966 = _T_5965 | _T_5711; // @[Mux.scala 27:72]
  wire [21:0] _T_5712 = _T_4196 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5967 = _T_5966 | _T_5712; // @[Mux.scala 27:72]
  wire [21:0] _T_5713 = _T_4198 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5968 = _T_5967 | _T_5713; // @[Mux.scala 27:72]
  wire [21:0] _T_5714 = _T_4200 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5969 = _T_5968 | _T_5714; // @[Mux.scala 27:72]
  wire [21:0] _T_5715 = _T_4202 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5970 = _T_5969 | _T_5715; // @[Mux.scala 27:72]
  wire [21:0] _T_5716 = _T_4204 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5971 = _T_5970 | _T_5716; // @[Mux.scala 27:72]
  wire [21:0] _T_5717 = _T_4206 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5972 = _T_5971 | _T_5717; // @[Mux.scala 27:72]
  wire [21:0] _T_5718 = _T_4208 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5973 = _T_5972 | _T_5718; // @[Mux.scala 27:72]
  wire [21:0] _T_5719 = _T_4210 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5974 = _T_5973 | _T_5719; // @[Mux.scala 27:72]
  wire [21:0] _T_5720 = _T_4212 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5975 = _T_5974 | _T_5720; // @[Mux.scala 27:72]
  wire [21:0] _T_5721 = _T_4214 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5976 = _T_5975 | _T_5721; // @[Mux.scala 27:72]
  wire [21:0] _T_5722 = _T_4216 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5977 = _T_5976 | _T_5722; // @[Mux.scala 27:72]
  wire [21:0] _T_5723 = _T_4218 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5978 = _T_5977 | _T_5723; // @[Mux.scala 27:72]
  wire [21:0] _T_5724 = _T_4220 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5979 = _T_5978 | _T_5724; // @[Mux.scala 27:72]
  wire [21:0] _T_5725 = _T_4222 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5980 = _T_5979 | _T_5725; // @[Mux.scala 27:72]
  wire [21:0] _T_5726 = _T_4224 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5981 = _T_5980 | _T_5726; // @[Mux.scala 27:72]
  wire [21:0] _T_5727 = _T_4226 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5982 = _T_5981 | _T_5727; // @[Mux.scala 27:72]
  wire [21:0] _T_5728 = _T_4228 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5983 = _T_5982 | _T_5728; // @[Mux.scala 27:72]
  wire [21:0] _T_5729 = _T_4230 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5984 = _T_5983 | _T_5729; // @[Mux.scala 27:72]
  wire [21:0] _T_5730 = _T_4232 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5985 = _T_5984 | _T_5730; // @[Mux.scala 27:72]
  wire [21:0] _T_5731 = _T_4234 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5986 = _T_5985 | _T_5731; // @[Mux.scala 27:72]
  wire [21:0] _T_5732 = _T_4236 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5987 = _T_5986 | _T_5732; // @[Mux.scala 27:72]
  wire [21:0] _T_5733 = _T_4238 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5988 = _T_5987 | _T_5733; // @[Mux.scala 27:72]
  wire [21:0] _T_5734 = _T_4240 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5989 = _T_5988 | _T_5734; // @[Mux.scala 27:72]
  wire [21:0] _T_5735 = _T_4242 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5990 = _T_5989 | _T_5735; // @[Mux.scala 27:72]
  wire [21:0] _T_5736 = _T_4244 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5991 = _T_5990 | _T_5736; // @[Mux.scala 27:72]
  wire [21:0] _T_5737 = _T_4246 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5992 = _T_5991 | _T_5737; // @[Mux.scala 27:72]
  wire [21:0] _T_5738 = _T_4248 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5993 = _T_5992 | _T_5738; // @[Mux.scala 27:72]
  wire [21:0] _T_5739 = _T_4250 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5994 = _T_5993 | _T_5739; // @[Mux.scala 27:72]
  wire [21:0] _T_5740 = _T_4252 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5995 = _T_5994 | _T_5740; // @[Mux.scala 27:72]
  wire [21:0] _T_5741 = _T_4254 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5996 = _T_5995 | _T_5741; // @[Mux.scala 27:72]
  wire [21:0] _T_5742 = _T_4256 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5997 = _T_5996 | _T_5742; // @[Mux.scala 27:72]
  wire [21:0] _T_5743 = _T_4258 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5998 = _T_5997 | _T_5743; // @[Mux.scala 27:72]
  wire [21:0] _T_5744 = _T_4260 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5999 = _T_5998 | _T_5744; // @[Mux.scala 27:72]
  wire [21:0] _T_5745 = _T_4262 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6000 = _T_5999 | _T_5745; // @[Mux.scala 27:72]
  wire [21:0] _T_5746 = _T_4264 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6001 = _T_6000 | _T_5746; // @[Mux.scala 27:72]
  wire [21:0] _T_5747 = _T_4266 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6002 = _T_6001 | _T_5747; // @[Mux.scala 27:72]
  wire [21:0] _T_5748 = _T_4268 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6003 = _T_6002 | _T_5748; // @[Mux.scala 27:72]
  wire [21:0] _T_5749 = _T_4270 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6004 = _T_6003 | _T_5749; // @[Mux.scala 27:72]
  wire [21:0] _T_5750 = _T_4272 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6005 = _T_6004 | _T_5750; // @[Mux.scala 27:72]
  wire [21:0] _T_5751 = _T_4274 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6006 = _T_6005 | _T_5751; // @[Mux.scala 27:72]
  wire [21:0] _T_5752 = _T_4276 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6007 = _T_6006 | _T_5752; // @[Mux.scala 27:72]
  wire [21:0] _T_5753 = _T_4278 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6008 = _T_6007 | _T_5753; // @[Mux.scala 27:72]
  wire [21:0] _T_5754 = _T_4280 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6009 = _T_6008 | _T_5754; // @[Mux.scala 27:72]
  wire [21:0] _T_5755 = _T_4282 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6010 = _T_6009 | _T_5755; // @[Mux.scala 27:72]
  wire [21:0] _T_5756 = _T_4284 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6011 = _T_6010 | _T_5756; // @[Mux.scala 27:72]
  wire [21:0] _T_5757 = _T_4286 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6012 = _T_6011 | _T_5757; // @[Mux.scala 27:72]
  wire [21:0] _T_5758 = _T_4288 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6013 = _T_6012 | _T_5758; // @[Mux.scala 27:72]
  wire [21:0] _T_5759 = _T_4290 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6014 = _T_6013 | _T_5759; // @[Mux.scala 27:72]
  wire [21:0] _T_5760 = _T_4292 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6015 = _T_6014 | _T_5760; // @[Mux.scala 27:72]
  wire [21:0] _T_5761 = _T_4294 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6016 = _T_6015 | _T_5761; // @[Mux.scala 27:72]
  wire [21:0] _T_5762 = _T_4296 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6017 = _T_6016 | _T_5762; // @[Mux.scala 27:72]
  wire [21:0] _T_5763 = _T_4298 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6018 = _T_6017 | _T_5763; // @[Mux.scala 27:72]
  wire [21:0] _T_5764 = _T_4300 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6019 = _T_6018 | _T_5764; // @[Mux.scala 27:72]
  wire [21:0] _T_5765 = _T_4302 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6020 = _T_6019 | _T_5765; // @[Mux.scala 27:72]
  wire [21:0] _T_5766 = _T_4304 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6021 = _T_6020 | _T_5766; // @[Mux.scala 27:72]
  wire [21:0] _T_5767 = _T_4306 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6022 = _T_6021 | _T_5767; // @[Mux.scala 27:72]
  wire [21:0] _T_5768 = _T_4308 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6023 = _T_6022 | _T_5768; // @[Mux.scala 27:72]
  wire [21:0] _T_5769 = _T_4310 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6024 = _T_6023 | _T_5769; // @[Mux.scala 27:72]
  wire [21:0] _T_5770 = _T_4312 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6025 = _T_6024 | _T_5770; // @[Mux.scala 27:72]
  wire [21:0] _T_5771 = _T_4314 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6026 = _T_6025 | _T_5771; // @[Mux.scala 27:72]
  wire [21:0] _T_5772 = _T_4316 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6027 = _T_6026 | _T_5772; // @[Mux.scala 27:72]
  wire [21:0] _T_5773 = _T_4318 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6028 = _T_6027 | _T_5773; // @[Mux.scala 27:72]
  wire [21:0] _T_5774 = _T_4320 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6029 = _T_6028 | _T_5774; // @[Mux.scala 27:72]
  wire [21:0] _T_5775 = _T_4322 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6030 = _T_6029 | _T_5775; // @[Mux.scala 27:72]
  wire [21:0] _T_5776 = _T_4324 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6031 = _T_6030 | _T_5776; // @[Mux.scala 27:72]
  wire [21:0] _T_5777 = _T_4326 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6032 = _T_6031 | _T_5777; // @[Mux.scala 27:72]
  wire [21:0] _T_5778 = _T_4328 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6033 = _T_6032 | _T_5778; // @[Mux.scala 27:72]
  wire [21:0] _T_5779 = _T_4330 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6034 = _T_6033 | _T_5779; // @[Mux.scala 27:72]
  wire [21:0] _T_5780 = _T_4332 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6035 = _T_6034 | _T_5780; // @[Mux.scala 27:72]
  wire [21:0] _T_5781 = _T_4334 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6036 = _T_6035 | _T_5781; // @[Mux.scala 27:72]
  wire [21:0] _T_5782 = _T_4336 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6037 = _T_6036 | _T_5782; // @[Mux.scala 27:72]
  wire [21:0] _T_5783 = _T_4338 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6038 = _T_6037 | _T_5783; // @[Mux.scala 27:72]
  wire [21:0] _T_5784 = _T_4340 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6039 = _T_6038 | _T_5784; // @[Mux.scala 27:72]
  wire [21:0] _T_5785 = _T_4342 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6040 = _T_6039 | _T_5785; // @[Mux.scala 27:72]
  wire [21:0] _T_5786 = _T_4344 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6041 = _T_6040 | _T_5786; // @[Mux.scala 27:72]
  wire [21:0] _T_5787 = _T_4346 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6042 = _T_6041 | _T_5787; // @[Mux.scala 27:72]
  wire [21:0] _T_5788 = _T_4348 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6043 = _T_6042 | _T_5788; // @[Mux.scala 27:72]
  wire [21:0] _T_5789 = _T_4350 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6044 = _T_6043 | _T_5789; // @[Mux.scala 27:72]
  wire [21:0] _T_5790 = _T_4352 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6045 = _T_6044 | _T_5790; // @[Mux.scala 27:72]
  wire [21:0] _T_5791 = _T_4354 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6046 = _T_6045 | _T_5791; // @[Mux.scala 27:72]
  wire [21:0] _T_5792 = _T_4356 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6047 = _T_6046 | _T_5792; // @[Mux.scala 27:72]
  wire [21:0] _T_5793 = _T_4358 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6048 = _T_6047 | _T_5793; // @[Mux.scala 27:72]
  wire [21:0] _T_5794 = _T_4360 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6049 = _T_6048 | _T_5794; // @[Mux.scala 27:72]
  wire [21:0] _T_5795 = _T_4362 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6050 = _T_6049 | _T_5795; // @[Mux.scala 27:72]
  wire [21:0] _T_5796 = _T_4364 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6051 = _T_6050 | _T_5796; // @[Mux.scala 27:72]
  wire [21:0] _T_5797 = _T_4366 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6052 = _T_6051 | _T_5797; // @[Mux.scala 27:72]
  wire [21:0] _T_5798 = _T_4368 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6053 = _T_6052 | _T_5798; // @[Mux.scala 27:72]
  wire [21:0] _T_5799 = _T_4370 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6054 = _T_6053 | _T_5799; // @[Mux.scala 27:72]
  wire [21:0] _T_5800 = _T_4372 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6055 = _T_6054 | _T_5800; // @[Mux.scala 27:72]
  wire [21:0] _T_5801 = _T_4374 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6056 = _T_6055 | _T_5801; // @[Mux.scala 27:72]
  wire [21:0] _T_5802 = _T_4376 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6057 = _T_6056 | _T_5802; // @[Mux.scala 27:72]
  wire [21:0] _T_5803 = _T_4378 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6058 = _T_6057 | _T_5803; // @[Mux.scala 27:72]
  wire [21:0] _T_5804 = _T_4380 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6059 = _T_6058 | _T_5804; // @[Mux.scala 27:72]
  wire [21:0] _T_5805 = _T_4382 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6060 = _T_6059 | _T_5805; // @[Mux.scala 27:72]
  wire [21:0] _T_5806 = _T_4384 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6061 = _T_6060 | _T_5806; // @[Mux.scala 27:72]
  wire [21:0] _T_5807 = _T_4386 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6062 = _T_6061 | _T_5807; // @[Mux.scala 27:72]
  wire [21:0] _T_5808 = _T_4388 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6063 = _T_6062 | _T_5808; // @[Mux.scala 27:72]
  wire [21:0] _T_5809 = _T_4390 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6064 = _T_6063 | _T_5809; // @[Mux.scala 27:72]
  wire [21:0] _T_5810 = _T_4392 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6065 = _T_6064 | _T_5810; // @[Mux.scala 27:72]
  wire [21:0] _T_5811 = _T_4394 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6066 = _T_6065 | _T_5811; // @[Mux.scala 27:72]
  wire [21:0] _T_5812 = _T_4396 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6067 = _T_6066 | _T_5812; // @[Mux.scala 27:72]
  wire [21:0] _T_5813 = _T_4398 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6068 = _T_6067 | _T_5813; // @[Mux.scala 27:72]
  wire [21:0] _T_5814 = _T_4400 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6069 = _T_6068 | _T_5814; // @[Mux.scala 27:72]
  wire [21:0] _T_5815 = _T_4402 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6070 = _T_6069 | _T_5815; // @[Mux.scala 27:72]
  wire [21:0] _T_5816 = _T_4404 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6071 = _T_6070 | _T_5816; // @[Mux.scala 27:72]
  wire [21:0] _T_5817 = _T_4406 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6072 = _T_6071 | _T_5817; // @[Mux.scala 27:72]
  wire [21:0] _T_5818 = _T_4408 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6073 = _T_6072 | _T_5818; // @[Mux.scala 27:72]
  wire [21:0] _T_5819 = _T_4410 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6074 = _T_6073 | _T_5819; // @[Mux.scala 27:72]
  wire [21:0] _T_5820 = _T_4412 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6075 = _T_6074 | _T_5820; // @[Mux.scala 27:72]
  wire [21:0] _T_5821 = _T_4414 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6076 = _T_6075 | _T_5821; // @[Mux.scala 27:72]
  wire [21:0] _T_5822 = _T_4416 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6077 = _T_6076 | _T_5822; // @[Mux.scala 27:72]
  wire [21:0] _T_5823 = _T_4418 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6078 = _T_6077 | _T_5823; // @[Mux.scala 27:72]
  wire [21:0] _T_5824 = _T_4420 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6079 = _T_6078 | _T_5824; // @[Mux.scala 27:72]
  wire [21:0] _T_5825 = _T_4422 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6080 = _T_6079 | _T_5825; // @[Mux.scala 27:72]
  wire [21:0] _T_5826 = _T_4424 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6081 = _T_6080 | _T_5826; // @[Mux.scala 27:72]
  wire [21:0] _T_5827 = _T_4426 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6082 = _T_6081 | _T_5827; // @[Mux.scala 27:72]
  wire [21:0] _T_5828 = _T_4428 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6083 = _T_6082 | _T_5828; // @[Mux.scala 27:72]
  wire [21:0] _T_5829 = _T_4430 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6084 = _T_6083 | _T_5829; // @[Mux.scala 27:72]
  wire [21:0] _T_5830 = _T_4432 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6085 = _T_6084 | _T_5830; // @[Mux.scala 27:72]
  wire [21:0] _T_5831 = _T_4434 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6086 = _T_6085 | _T_5831; // @[Mux.scala 27:72]
  wire [21:0] _T_5832 = _T_4436 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6087 = _T_6086 | _T_5832; // @[Mux.scala 27:72]
  wire [21:0] _T_5833 = _T_4438 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6088 = _T_6087 | _T_5833; // @[Mux.scala 27:72]
  wire [21:0] _T_5834 = _T_4440 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6089 = _T_6088 | _T_5834; // @[Mux.scala 27:72]
  wire [21:0] _T_5835 = _T_4442 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6090 = _T_6089 | _T_5835; // @[Mux.scala 27:72]
  wire [21:0] _T_5836 = _T_4444 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6091 = _T_6090 | _T_5836; // @[Mux.scala 27:72]
  wire [21:0] _T_5837 = _T_4446 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6092 = _T_6091 | _T_5837; // @[Mux.scala 27:72]
  wire [21:0] _T_5838 = _T_4448 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6093 = _T_6092 | _T_5838; // @[Mux.scala 27:72]
  wire [21:0] _T_5839 = _T_4450 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6094 = _T_6093 | _T_5839; // @[Mux.scala 27:72]
  wire [21:0] _T_5840 = _T_4452 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6095 = _T_6094 | _T_5840; // @[Mux.scala 27:72]
  wire [21:0] _T_5841 = _T_4454 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6096 = _T_6095 | _T_5841; // @[Mux.scala 27:72]
  wire [21:0] _T_5842 = _T_4456 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6097 = _T_6096 | _T_5842; // @[Mux.scala 27:72]
  wire [21:0] _T_5843 = _T_4458 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6098 = _T_6097 | _T_5843; // @[Mux.scala 27:72]
  wire [21:0] _T_5844 = _T_4460 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6099 = _T_6098 | _T_5844; // @[Mux.scala 27:72]
  wire [21:0] _T_5845 = _T_4462 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6100 = _T_6099 | _T_5845; // @[Mux.scala 27:72]
  wire [21:0] _T_5846 = _T_4464 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6101 = _T_6100 | _T_5846; // @[Mux.scala 27:72]
  wire [21:0] _T_5847 = _T_4466 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6102 = _T_6101 | _T_5847; // @[Mux.scala 27:72]
  wire [21:0] _T_5848 = _T_4468 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6103 = _T_6102 | _T_5848; // @[Mux.scala 27:72]
  wire [21:0] _T_5849 = _T_4470 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6104 = _T_6103 | _T_5849; // @[Mux.scala 27:72]
  wire [21:0] _T_5850 = _T_4472 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6105 = _T_6104 | _T_5850; // @[Mux.scala 27:72]
  wire [21:0] _T_5851 = _T_4474 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6106 = _T_6105 | _T_5851; // @[Mux.scala 27:72]
  wire [21:0] _T_5852 = _T_4476 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6107 = _T_6106 | _T_5852; // @[Mux.scala 27:72]
  wire [21:0] _T_5853 = _T_4478 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6108 = _T_6107 | _T_5853; // @[Mux.scala 27:72]
  wire [21:0] _T_5854 = _T_4480 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6109 = _T_6108 | _T_5854; // @[Mux.scala 27:72]
  wire [21:0] _T_5855 = _T_4482 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6110 = _T_6109 | _T_5855; // @[Mux.scala 27:72]
  wire [21:0] _T_5856 = _T_4484 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6111 = _T_6110 | _T_5856; // @[Mux.scala 27:72]
  wire [21:0] _T_5857 = _T_4486 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6112 = _T_6111 | _T_5857; // @[Mux.scala 27:72]
  wire [21:0] _T_5858 = _T_4488 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6113 = _T_6112 | _T_5858; // @[Mux.scala 27:72]
  wire [21:0] _T_5859 = _T_4490 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6114 = _T_6113 | _T_5859; // @[Mux.scala 27:72]
  wire [21:0] _T_5860 = _T_4492 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6115 = _T_6114 | _T_5860; // @[Mux.scala 27:72]
  wire [21:0] _T_5861 = _T_4494 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6116 = _T_6115 | _T_5861; // @[Mux.scala 27:72]
  wire [21:0] _T_5862 = _T_4496 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6117 = _T_6116 | _T_5862; // @[Mux.scala 27:72]
  wire [21:0] _T_5863 = _T_4498 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6118 = _T_6117 | _T_5863; // @[Mux.scala 27:72]
  wire [21:0] _T_5864 = _T_4500 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6119 = _T_6118 | _T_5864; // @[Mux.scala 27:72]
  wire [21:0] _T_5865 = _T_4502 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6120 = _T_6119 | _T_5865; // @[Mux.scala 27:72]
  wire [21:0] _T_5866 = _T_4504 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6121 = _T_6120 | _T_5866; // @[Mux.scala 27:72]
  wire [21:0] _T_5867 = _T_4506 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6122 = _T_6121 | _T_5867; // @[Mux.scala 27:72]
  wire [21:0] _T_5868 = _T_4508 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6123 = _T_6122 | _T_5868; // @[Mux.scala 27:72]
  wire [21:0] _T_5869 = _T_4510 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6124 = _T_6123 | _T_5869; // @[Mux.scala 27:72]
  wire [21:0] _T_5870 = _T_4512 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6125 = _T_6124 | _T_5870; // @[Mux.scala 27:72]
  wire [21:0] _T_5871 = _T_4514 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6126 = _T_6125 | _T_5871; // @[Mux.scala 27:72]
  wire [21:0] _T_5872 = _T_4516 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6127 = _T_6126 | _T_5872; // @[Mux.scala 27:72]
  wire [21:0] _T_5873 = _T_4518 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6128 = _T_6127 | _T_5873; // @[Mux.scala 27:72]
  wire [21:0] _T_5874 = _T_4520 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6129 = _T_6128 | _T_5874; // @[Mux.scala 27:72]
  wire [21:0] _T_5875 = _T_4522 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6130 = _T_6129 | _T_5875; // @[Mux.scala 27:72]
  wire [21:0] _T_5876 = _T_4524 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6131 = _T_6130 | _T_5876; // @[Mux.scala 27:72]
  wire [21:0] _T_5877 = _T_4526 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6132 = _T_6131 | _T_5877; // @[Mux.scala 27:72]
  wire [21:0] _T_5878 = _T_4528 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6133 = _T_6132 | _T_5878; // @[Mux.scala 27:72]
  wire [21:0] _T_5879 = _T_4530 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6134 = _T_6133 | _T_5879; // @[Mux.scala 27:72]
  wire [21:0] _T_5880 = _T_4532 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6135 = _T_6134 | _T_5880; // @[Mux.scala 27:72]
  wire [21:0] _T_5881 = _T_4534 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6136 = _T_6135 | _T_5881; // @[Mux.scala 27:72]
  wire [21:0] _T_5882 = _T_4536 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6137 = _T_6136 | _T_5882; // @[Mux.scala 27:72]
  wire [21:0] _T_5883 = _T_4538 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6138 = _T_6137 | _T_5883; // @[Mux.scala 27:72]
  wire [21:0] _T_5884 = _T_4540 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6139 = _T_6138 | _T_5884; // @[Mux.scala 27:72]
  wire [21:0] _T_5885 = _T_4542 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6140 = _T_6139 | _T_5885; // @[Mux.scala 27:72]
  wire [21:0] _T_5886 = _T_4544 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6141 = _T_6140 | _T_5886; // @[Mux.scala 27:72]
  wire [21:0] _T_5887 = _T_4546 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6142 = _T_6141 | _T_5887; // @[Mux.scala 27:72]
  wire [21:0] _T_5888 = _T_4548 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6143 = _T_6142 | _T_5888; // @[Mux.scala 27:72]
  wire [21:0] _T_5889 = _T_4550 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6144 = _T_6143 | _T_5889; // @[Mux.scala 27:72]
  wire [21:0] _T_5890 = _T_4552 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6145 = _T_6144 | _T_5890; // @[Mux.scala 27:72]
  wire [21:0] _T_5891 = _T_4554 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6146 = _T_6145 | _T_5891; // @[Mux.scala 27:72]
  wire [21:0] _T_5892 = _T_4556 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6147 = _T_6146 | _T_5892; // @[Mux.scala 27:72]
  wire [21:0] _T_5893 = _T_4558 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6148 = _T_6147 | _T_5893; // @[Mux.scala 27:72]
  wire [21:0] _T_5894 = _T_4560 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6149 = _T_6148 | _T_5894; // @[Mux.scala 27:72]
  wire [21:0] _T_5895 = _T_4562 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6150 = _T_6149 | _T_5895; // @[Mux.scala 27:72]
  wire [21:0] _T_5896 = _T_4564 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6151 = _T_6150 | _T_5896; // @[Mux.scala 27:72]
  wire [21:0] _T_5897 = _T_4566 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6152 = _T_6151 | _T_5897; // @[Mux.scala 27:72]
  wire [21:0] _T_5898 = _T_4568 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6153 = _T_6152 | _T_5898; // @[Mux.scala 27:72]
  wire [21:0] _T_5899 = _T_4570 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6154 = _T_6153 | _T_5899; // @[Mux.scala 27:72]
  wire [21:0] _T_5900 = _T_4572 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6155 = _T_6154 | _T_5900; // @[Mux.scala 27:72]
  wire [21:0] _T_5901 = _T_4574 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6156 = _T_6155 | _T_5901; // @[Mux.scala 27:72]
  wire [21:0] _T_5902 = _T_4576 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6157 = _T_6156 | _T_5902; // @[Mux.scala 27:72]
  wire [21:0] _T_5903 = _T_4578 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6158 = _T_6157 | _T_5903; // @[Mux.scala 27:72]
  wire [21:0] _T_5904 = _T_4580 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6159 = _T_6158 | _T_5904; // @[Mux.scala 27:72]
  wire [21:0] _T_5905 = _T_4582 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6160 = _T_6159 | _T_5905; // @[Mux.scala 27:72]
  wire [21:0] _T_5906 = _T_4584 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6161 = _T_6160 | _T_5906; // @[Mux.scala 27:72]
  wire [21:0] _T_5907 = _T_4586 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6162 = _T_6161 | _T_5907; // @[Mux.scala 27:72]
  wire [21:0] _T_5908 = _T_4588 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6163 = _T_6162 | _T_5908; // @[Mux.scala 27:72]
  wire [21:0] _T_5909 = _T_4590 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6164 = _T_6163 | _T_5909; // @[Mux.scala 27:72]
  wire [21:0] _T_5910 = _T_4592 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6165 = _T_6164 | _T_5910; // @[Mux.scala 27:72]
  wire [21:0] _T_5911 = _T_4594 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6166 = _T_6165 | _T_5911; // @[Mux.scala 27:72]
  wire [21:0] _T_5912 = _T_4596 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6167 = _T_6166 | _T_5912; // @[Mux.scala 27:72]
  wire [21:0] _T_5913 = _T_4598 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6168 = _T_6167 | _T_5913; // @[Mux.scala 27:72]
  wire [21:0] _T_5914 = _T_4600 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6169 = _T_6168 | _T_5914; // @[Mux.scala 27:72]
  wire [21:0] _T_5915 = _T_4602 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6170 = _T_6169 | _T_5915; // @[Mux.scala 27:72]
  wire [21:0] _T_5916 = _T_4604 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6171 = _T_6170 | _T_5916; // @[Mux.scala 27:72]
  wire [21:0] _T_5917 = _T_4606 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6172 = _T_6171 | _T_5917; // @[Mux.scala 27:72]
  wire [21:0] _T_5918 = _T_4608 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6173 = _T_6172 | _T_5918; // @[Mux.scala 27:72]
  wire [21:0] _T_5919 = _T_4610 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6174 = _T_6173 | _T_5919; // @[Mux.scala 27:72]
  wire [21:0] _T_5920 = _T_4612 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6175 = _T_6174 | _T_5920; // @[Mux.scala 27:72]
  wire [21:0] _T_5921 = _T_4614 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6176 = _T_6175 | _T_5921; // @[Mux.scala 27:72]
  wire [21:0] _T_5922 = _T_4616 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6177 = _T_6176 | _T_5922; // @[Mux.scala 27:72]
  wire [21:0] _T_5923 = _T_4618 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6178 = _T_6177 | _T_5923; // @[Mux.scala 27:72]
  wire [21:0] _T_5924 = _T_4620 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6179 = _T_6178 | _T_5924; // @[Mux.scala 27:72]
  wire [21:0] _T_5925 = _T_4622 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6180 = _T_6179 | _T_5925; // @[Mux.scala 27:72]
  wire [21:0] _T_5926 = _T_4624 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6181 = _T_6180 | _T_5926; // @[Mux.scala 27:72]
  wire [21:0] _T_5927 = _T_4626 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6182 = _T_6181 | _T_5927; // @[Mux.scala 27:72]
  wire [21:0] _T_5928 = _T_4628 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6183 = _T_6182 | _T_5928; // @[Mux.scala 27:72]
  wire [21:0] _T_5929 = _T_4630 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6184 = _T_6183 | _T_5929; // @[Mux.scala 27:72]
  wire [21:0] _T_5930 = _T_4632 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6185 = _T_6184 | _T_5930; // @[Mux.scala 27:72]
  wire [21:0] _T_5931 = _T_4634 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6186 = _T_6185 | _T_5931; // @[Mux.scala 27:72]
  wire [21:0] _T_5932 = _T_4636 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6187 = _T_6186 | _T_5932; // @[Mux.scala 27:72]
  wire [21:0] _T_5933 = _T_4638 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6188 = _T_6187 | _T_5933; // @[Mux.scala 27:72]
  wire [21:0] _T_5934 = _T_4640 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6189 = _T_6188 | _T_5934; // @[Mux.scala 27:72]
  wire [21:0] _T_5935 = _T_4642 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6190 = _T_6189 | _T_5935; // @[Mux.scala 27:72]
  wire [21:0] _T_5936 = _T_4644 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6191 = _T_6190 | _T_5936; // @[Mux.scala 27:72]
  wire [21:0] _T_5937 = _T_4646 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6192 = _T_6191 | _T_5937; // @[Mux.scala 27:72]
  wire [21:0] _T_5938 = _T_4648 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6193 = _T_6192 | _T_5938; // @[Mux.scala 27:72]
  wire [21:0] _T_5939 = _T_4650 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6194 = _T_6193 | _T_5939; // @[Mux.scala 27:72]
  wire [21:0] _T_5940 = _T_4652 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6195 = _T_6194 | _T_5940; // @[Mux.scala 27:72]
  wire [21:0] _T_5941 = _T_4654 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6196 = _T_6195 | _T_5941; // @[Mux.scala 27:72]
  wire [21:0] _T_5942 = _T_4656 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6197 = _T_6196 | _T_5942; // @[Mux.scala 27:72]
  wire [21:0] _T_5943 = _T_4658 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6198 = _T_6197 | _T_5943; // @[Mux.scala 27:72]
  wire [21:0] _T_5944 = _T_4660 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6199 = _T_6198 | _T_5944; // @[Mux.scala 27:72]
  wire [21:0] _T_5945 = _T_4662 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6200 = _T_6199 | _T_5945; // @[Mux.scala 27:72]
  wire [21:0] _T_5946 = _T_4664 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6201 = _T_6200 | _T_5946; // @[Mux.scala 27:72]
  wire [21:0] _T_5947 = _T_4666 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6201 | _T_5947; // @[Mux.scala 27:72]
  wire  _T_72 = btb_bank0_rd_data_way1_p1_f[21:17] == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 145:106]
  wire  _T_73 = btb_bank0_rd_data_way1_p1_f[0] & _T_72; // @[el2_ifu_bp_ctl.scala 145:61]
  wire  _T_76 = _T_73 & _T_48; // @[el2_ifu_bp_ctl.scala 145:129]
  wire  _T_77 = _T_76 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 146:56]
  wire  tag_match_way1_p1_f = _T_77 & _T; // @[el2_ifu_bp_ctl.scala 146:77]
  wire  _T_108 = btb_bank0_rd_data_way1_p1_f[3] ^ btb_bank0_rd_data_way1_p1_f[4]; // @[el2_ifu_bp_ctl.scala 159:100]
  wire  _T_109 = tag_match_way1_p1_f & _T_108; // @[el2_ifu_bp_ctl.scala 159:62]
  wire  _T_113 = ~_T_108; // @[el2_ifu_bp_ctl.scala 160:64]
  wire  _T_114 = tag_match_way1_p1_f & _T_113; // @[el2_ifu_bp_ctl.scala 160:62]
  wire [1:0] tag_match_way1_expanded_p1_f = {_T_109,_T_114}; // @[Cat.scala 29:58]
  wire [21:0] _T_134 = tag_match_way1_expanded_p1_f[1] ? btb_bank0_rd_data_way1_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_p1_f = _T_133 | _T_134; // @[Mux.scala 27:72]
  wire [21:0] _T_146 = io_ifc_fetch_addr_f[0] ? btb_bank0e_rd_data_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_145 | _T_146; // @[Mux.scala 27:72]
  wire  _T_241 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 236:59]
  wire [21:0] _T_119 = tag_match_way0_expanded_f[0] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_120 = tag_match_way1_expanded_f[0] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_f = _T_119 | _T_120; // @[Mux.scala 27:72]
  wire [21:0] _T_139 = _T_143 ? btb_bank0e_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_140 = io_ifc_fetch_addr_f[0] ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_139 | _T_140; // @[Mux.scala 27:72]
  wire  _T_244 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 237:59]
  wire [1:0] bht_force_taken_f = {_T_241,_T_244}; // @[Cat.scala 29:58]
  wire [9:0] _T_566 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[el2_ifu_bp_ctl.scala 284:18]
  wire [7:0] bht_rd_addr_f = _T_566[9:2] ^ fghr; // @[el2_lib.scala 188:35]
  wire  _T_20797 = bht_rd_addr_f == 8'h0; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_21564 = _T_20797 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_20800 = bht_rd_addr_f == 8'h1; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_21565 = _T_20800 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21820 = _T_21564 | _T_21565; // @[Mux.scala 27:72]
  wire  _T_20803 = bht_rd_addr_f == 8'h2; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_21566 = _T_20803 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21821 = _T_21820 | _T_21566; // @[Mux.scala 27:72]
  wire  _T_20806 = bht_rd_addr_f == 8'h3; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_21567 = _T_20806 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21822 = _T_21821 | _T_21567; // @[Mux.scala 27:72]
  wire  _T_20809 = bht_rd_addr_f == 8'h4; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_21568 = _T_20809 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21823 = _T_21822 | _T_21568; // @[Mux.scala 27:72]
  wire  _T_20812 = bht_rd_addr_f == 8'h5; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_21569 = _T_20812 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21824 = _T_21823 | _T_21569; // @[Mux.scala 27:72]
  wire  _T_20815 = bht_rd_addr_f == 8'h6; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_21570 = _T_20815 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21825 = _T_21824 | _T_21570; // @[Mux.scala 27:72]
  wire  _T_20818 = bht_rd_addr_f == 8'h7; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_21571 = _T_20818 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21826 = _T_21825 | _T_21571; // @[Mux.scala 27:72]
  wire  _T_20821 = bht_rd_addr_f == 8'h8; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_21572 = _T_20821 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21827 = _T_21826 | _T_21572; // @[Mux.scala 27:72]
  wire  _T_20824 = bht_rd_addr_f == 8'h9; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_21573 = _T_20824 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21828 = _T_21827 | _T_21573; // @[Mux.scala 27:72]
  wire  _T_20827 = bht_rd_addr_f == 8'ha; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_21574 = _T_20827 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21829 = _T_21828 | _T_21574; // @[Mux.scala 27:72]
  wire  _T_20830 = bht_rd_addr_f == 8'hb; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_21575 = _T_20830 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21830 = _T_21829 | _T_21575; // @[Mux.scala 27:72]
  wire  _T_20833 = bht_rd_addr_f == 8'hc; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_21576 = _T_20833 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21831 = _T_21830 | _T_21576; // @[Mux.scala 27:72]
  wire  _T_20836 = bht_rd_addr_f == 8'hd; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_21577 = _T_20836 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21832 = _T_21831 | _T_21577; // @[Mux.scala 27:72]
  wire  _T_20839 = bht_rd_addr_f == 8'he; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_21578 = _T_20839 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21833 = _T_21832 | _T_21578; // @[Mux.scala 27:72]
  wire  _T_20842 = bht_rd_addr_f == 8'hf; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_21579 = _T_20842 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21834 = _T_21833 | _T_21579; // @[Mux.scala 27:72]
  wire  _T_20845 = bht_rd_addr_f == 8'h10; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_21580 = _T_20845 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21835 = _T_21834 | _T_21580; // @[Mux.scala 27:72]
  wire  _T_20848 = bht_rd_addr_f == 8'h11; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_21581 = _T_20848 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21836 = _T_21835 | _T_21581; // @[Mux.scala 27:72]
  wire  _T_20851 = bht_rd_addr_f == 8'h12; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_21582 = _T_20851 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21837 = _T_21836 | _T_21582; // @[Mux.scala 27:72]
  wire  _T_20854 = bht_rd_addr_f == 8'h13; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_21583 = _T_20854 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21838 = _T_21837 | _T_21583; // @[Mux.scala 27:72]
  wire  _T_20857 = bht_rd_addr_f == 8'h14; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_21584 = _T_20857 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21839 = _T_21838 | _T_21584; // @[Mux.scala 27:72]
  wire  _T_20860 = bht_rd_addr_f == 8'h15; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_21585 = _T_20860 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21840 = _T_21839 | _T_21585; // @[Mux.scala 27:72]
  wire  _T_20863 = bht_rd_addr_f == 8'h16; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_21586 = _T_20863 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21841 = _T_21840 | _T_21586; // @[Mux.scala 27:72]
  wire  _T_20866 = bht_rd_addr_f == 8'h17; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_21587 = _T_20866 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21842 = _T_21841 | _T_21587; // @[Mux.scala 27:72]
  wire  _T_20869 = bht_rd_addr_f == 8'h18; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_21588 = _T_20869 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21843 = _T_21842 | _T_21588; // @[Mux.scala 27:72]
  wire  _T_20872 = bht_rd_addr_f == 8'h19; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_21589 = _T_20872 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21844 = _T_21843 | _T_21589; // @[Mux.scala 27:72]
  wire  _T_20875 = bht_rd_addr_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_21590 = _T_20875 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21845 = _T_21844 | _T_21590; // @[Mux.scala 27:72]
  wire  _T_20878 = bht_rd_addr_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_21591 = _T_20878 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21846 = _T_21845 | _T_21591; // @[Mux.scala 27:72]
  wire  _T_20881 = bht_rd_addr_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_21592 = _T_20881 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21847 = _T_21846 | _T_21592; // @[Mux.scala 27:72]
  wire  _T_20884 = bht_rd_addr_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_21593 = _T_20884 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21848 = _T_21847 | _T_21593; // @[Mux.scala 27:72]
  wire  _T_20887 = bht_rd_addr_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_21594 = _T_20887 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21849 = _T_21848 | _T_21594; // @[Mux.scala 27:72]
  wire  _T_20890 = bht_rd_addr_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_21595 = _T_20890 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21850 = _T_21849 | _T_21595; // @[Mux.scala 27:72]
  wire  _T_20893 = bht_rd_addr_f == 8'h20; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_21596 = _T_20893 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21851 = _T_21850 | _T_21596; // @[Mux.scala 27:72]
  wire  _T_20896 = bht_rd_addr_f == 8'h21; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_21597 = _T_20896 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21852 = _T_21851 | _T_21597; // @[Mux.scala 27:72]
  wire  _T_20899 = bht_rd_addr_f == 8'h22; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_21598 = _T_20899 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21853 = _T_21852 | _T_21598; // @[Mux.scala 27:72]
  wire  _T_20902 = bht_rd_addr_f == 8'h23; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_21599 = _T_20902 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21854 = _T_21853 | _T_21599; // @[Mux.scala 27:72]
  wire  _T_20905 = bht_rd_addr_f == 8'h24; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_21600 = _T_20905 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21855 = _T_21854 | _T_21600; // @[Mux.scala 27:72]
  wire  _T_20908 = bht_rd_addr_f == 8'h25; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_21601 = _T_20908 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21856 = _T_21855 | _T_21601; // @[Mux.scala 27:72]
  wire  _T_20911 = bht_rd_addr_f == 8'h26; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_21602 = _T_20911 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21857 = _T_21856 | _T_21602; // @[Mux.scala 27:72]
  wire  _T_20914 = bht_rd_addr_f == 8'h27; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_21603 = _T_20914 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21858 = _T_21857 | _T_21603; // @[Mux.scala 27:72]
  wire  _T_20917 = bht_rd_addr_f == 8'h28; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_21604 = _T_20917 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21859 = _T_21858 | _T_21604; // @[Mux.scala 27:72]
  wire  _T_20920 = bht_rd_addr_f == 8'h29; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_21605 = _T_20920 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21860 = _T_21859 | _T_21605; // @[Mux.scala 27:72]
  wire  _T_20923 = bht_rd_addr_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_21606 = _T_20923 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21861 = _T_21860 | _T_21606; // @[Mux.scala 27:72]
  wire  _T_20926 = bht_rd_addr_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_21607 = _T_20926 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21862 = _T_21861 | _T_21607; // @[Mux.scala 27:72]
  wire  _T_20929 = bht_rd_addr_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_21608 = _T_20929 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21863 = _T_21862 | _T_21608; // @[Mux.scala 27:72]
  wire  _T_20932 = bht_rd_addr_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_21609 = _T_20932 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21864 = _T_21863 | _T_21609; // @[Mux.scala 27:72]
  wire  _T_20935 = bht_rd_addr_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_21610 = _T_20935 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21865 = _T_21864 | _T_21610; // @[Mux.scala 27:72]
  wire  _T_20938 = bht_rd_addr_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_21611 = _T_20938 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21866 = _T_21865 | _T_21611; // @[Mux.scala 27:72]
  wire  _T_20941 = bht_rd_addr_f == 8'h30; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_21612 = _T_20941 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21867 = _T_21866 | _T_21612; // @[Mux.scala 27:72]
  wire  _T_20944 = bht_rd_addr_f == 8'h31; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_21613 = _T_20944 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21868 = _T_21867 | _T_21613; // @[Mux.scala 27:72]
  wire  _T_20947 = bht_rd_addr_f == 8'h32; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_21614 = _T_20947 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21869 = _T_21868 | _T_21614; // @[Mux.scala 27:72]
  wire  _T_20950 = bht_rd_addr_f == 8'h33; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_21615 = _T_20950 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21870 = _T_21869 | _T_21615; // @[Mux.scala 27:72]
  wire  _T_20953 = bht_rd_addr_f == 8'h34; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_21616 = _T_20953 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21871 = _T_21870 | _T_21616; // @[Mux.scala 27:72]
  wire  _T_20956 = bht_rd_addr_f == 8'h35; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_21617 = _T_20956 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21872 = _T_21871 | _T_21617; // @[Mux.scala 27:72]
  wire  _T_20959 = bht_rd_addr_f == 8'h36; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_21618 = _T_20959 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21873 = _T_21872 | _T_21618; // @[Mux.scala 27:72]
  wire  _T_20962 = bht_rd_addr_f == 8'h37; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_21619 = _T_20962 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21874 = _T_21873 | _T_21619; // @[Mux.scala 27:72]
  wire  _T_20965 = bht_rd_addr_f == 8'h38; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_21620 = _T_20965 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21875 = _T_21874 | _T_21620; // @[Mux.scala 27:72]
  wire  _T_20968 = bht_rd_addr_f == 8'h39; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_21621 = _T_20968 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21876 = _T_21875 | _T_21621; // @[Mux.scala 27:72]
  wire  _T_20971 = bht_rd_addr_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_21622 = _T_20971 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21877 = _T_21876 | _T_21622; // @[Mux.scala 27:72]
  wire  _T_20974 = bht_rd_addr_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_21623 = _T_20974 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21878 = _T_21877 | _T_21623; // @[Mux.scala 27:72]
  wire  _T_20977 = bht_rd_addr_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_21624 = _T_20977 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21879 = _T_21878 | _T_21624; // @[Mux.scala 27:72]
  wire  _T_20980 = bht_rd_addr_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_21625 = _T_20980 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21880 = _T_21879 | _T_21625; // @[Mux.scala 27:72]
  wire  _T_20983 = bht_rd_addr_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_21626 = _T_20983 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21881 = _T_21880 | _T_21626; // @[Mux.scala 27:72]
  wire  _T_20986 = bht_rd_addr_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_21627 = _T_20986 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21882 = _T_21881 | _T_21627; // @[Mux.scala 27:72]
  wire  _T_20989 = bht_rd_addr_f == 8'h40; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_21628 = _T_20989 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21883 = _T_21882 | _T_21628; // @[Mux.scala 27:72]
  wire  _T_20992 = bht_rd_addr_f == 8'h41; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_21629 = _T_20992 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21884 = _T_21883 | _T_21629; // @[Mux.scala 27:72]
  wire  _T_20995 = bht_rd_addr_f == 8'h42; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_21630 = _T_20995 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21885 = _T_21884 | _T_21630; // @[Mux.scala 27:72]
  wire  _T_20998 = bht_rd_addr_f == 8'h43; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_21631 = _T_20998 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21886 = _T_21885 | _T_21631; // @[Mux.scala 27:72]
  wire  _T_21001 = bht_rd_addr_f == 8'h44; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_21632 = _T_21001 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21887 = _T_21886 | _T_21632; // @[Mux.scala 27:72]
  wire  _T_21004 = bht_rd_addr_f == 8'h45; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_21633 = _T_21004 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21888 = _T_21887 | _T_21633; // @[Mux.scala 27:72]
  wire  _T_21007 = bht_rd_addr_f == 8'h46; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_21634 = _T_21007 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21889 = _T_21888 | _T_21634; // @[Mux.scala 27:72]
  wire  _T_21010 = bht_rd_addr_f == 8'h47; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_21635 = _T_21010 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21890 = _T_21889 | _T_21635; // @[Mux.scala 27:72]
  wire  _T_21013 = bht_rd_addr_f == 8'h48; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_21636 = _T_21013 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21891 = _T_21890 | _T_21636; // @[Mux.scala 27:72]
  wire  _T_21016 = bht_rd_addr_f == 8'h49; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_21637 = _T_21016 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21892 = _T_21891 | _T_21637; // @[Mux.scala 27:72]
  wire  _T_21019 = bht_rd_addr_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_21638 = _T_21019 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21893 = _T_21892 | _T_21638; // @[Mux.scala 27:72]
  wire  _T_21022 = bht_rd_addr_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_21639 = _T_21022 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21894 = _T_21893 | _T_21639; // @[Mux.scala 27:72]
  wire  _T_21025 = bht_rd_addr_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_21640 = _T_21025 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21895 = _T_21894 | _T_21640; // @[Mux.scala 27:72]
  wire  _T_21028 = bht_rd_addr_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_21641 = _T_21028 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21896 = _T_21895 | _T_21641; // @[Mux.scala 27:72]
  wire  _T_21031 = bht_rd_addr_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_21642 = _T_21031 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21897 = _T_21896 | _T_21642; // @[Mux.scala 27:72]
  wire  _T_21034 = bht_rd_addr_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_21643 = _T_21034 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21898 = _T_21897 | _T_21643; // @[Mux.scala 27:72]
  wire  _T_21037 = bht_rd_addr_f == 8'h50; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_21644 = _T_21037 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21899 = _T_21898 | _T_21644; // @[Mux.scala 27:72]
  wire  _T_21040 = bht_rd_addr_f == 8'h51; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_21645 = _T_21040 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21900 = _T_21899 | _T_21645; // @[Mux.scala 27:72]
  wire  _T_21043 = bht_rd_addr_f == 8'h52; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_21646 = _T_21043 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21901 = _T_21900 | _T_21646; // @[Mux.scala 27:72]
  wire  _T_21046 = bht_rd_addr_f == 8'h53; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_21647 = _T_21046 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21902 = _T_21901 | _T_21647; // @[Mux.scala 27:72]
  wire  _T_21049 = bht_rd_addr_f == 8'h54; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_21648 = _T_21049 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21903 = _T_21902 | _T_21648; // @[Mux.scala 27:72]
  wire  _T_21052 = bht_rd_addr_f == 8'h55; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_21649 = _T_21052 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21904 = _T_21903 | _T_21649; // @[Mux.scala 27:72]
  wire  _T_21055 = bht_rd_addr_f == 8'h56; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_21650 = _T_21055 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21905 = _T_21904 | _T_21650; // @[Mux.scala 27:72]
  wire  _T_21058 = bht_rd_addr_f == 8'h57; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_21651 = _T_21058 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21906 = _T_21905 | _T_21651; // @[Mux.scala 27:72]
  wire  _T_21061 = bht_rd_addr_f == 8'h58; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_21652 = _T_21061 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21907 = _T_21906 | _T_21652; // @[Mux.scala 27:72]
  wire  _T_21064 = bht_rd_addr_f == 8'h59; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_21653 = _T_21064 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21908 = _T_21907 | _T_21653; // @[Mux.scala 27:72]
  wire  _T_21067 = bht_rd_addr_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_21654 = _T_21067 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21909 = _T_21908 | _T_21654; // @[Mux.scala 27:72]
  wire  _T_21070 = bht_rd_addr_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_21655 = _T_21070 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21910 = _T_21909 | _T_21655; // @[Mux.scala 27:72]
  wire  _T_21073 = bht_rd_addr_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_21656 = _T_21073 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21911 = _T_21910 | _T_21656; // @[Mux.scala 27:72]
  wire  _T_21076 = bht_rd_addr_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_21657 = _T_21076 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21912 = _T_21911 | _T_21657; // @[Mux.scala 27:72]
  wire  _T_21079 = bht_rd_addr_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_21658 = _T_21079 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21913 = _T_21912 | _T_21658; // @[Mux.scala 27:72]
  wire  _T_21082 = bht_rd_addr_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_21659 = _T_21082 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21914 = _T_21913 | _T_21659; // @[Mux.scala 27:72]
  wire  _T_21085 = bht_rd_addr_f == 8'h60; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_21660 = _T_21085 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21915 = _T_21914 | _T_21660; // @[Mux.scala 27:72]
  wire  _T_21088 = bht_rd_addr_f == 8'h61; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_21661 = _T_21088 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21916 = _T_21915 | _T_21661; // @[Mux.scala 27:72]
  wire  _T_21091 = bht_rd_addr_f == 8'h62; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_21662 = _T_21091 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21917 = _T_21916 | _T_21662; // @[Mux.scala 27:72]
  wire  _T_21094 = bht_rd_addr_f == 8'h63; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_21663 = _T_21094 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21918 = _T_21917 | _T_21663; // @[Mux.scala 27:72]
  wire  _T_21097 = bht_rd_addr_f == 8'h64; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_21664 = _T_21097 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21919 = _T_21918 | _T_21664; // @[Mux.scala 27:72]
  wire  _T_21100 = bht_rd_addr_f == 8'h65; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_21665 = _T_21100 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21920 = _T_21919 | _T_21665; // @[Mux.scala 27:72]
  wire  _T_21103 = bht_rd_addr_f == 8'h66; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_21666 = _T_21103 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21921 = _T_21920 | _T_21666; // @[Mux.scala 27:72]
  wire  _T_21106 = bht_rd_addr_f == 8'h67; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_21667 = _T_21106 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21922 = _T_21921 | _T_21667; // @[Mux.scala 27:72]
  wire  _T_21109 = bht_rd_addr_f == 8'h68; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_21668 = _T_21109 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21923 = _T_21922 | _T_21668; // @[Mux.scala 27:72]
  wire  _T_21112 = bht_rd_addr_f == 8'h69; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_21669 = _T_21112 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21924 = _T_21923 | _T_21669; // @[Mux.scala 27:72]
  wire  _T_21115 = bht_rd_addr_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_21670 = _T_21115 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21925 = _T_21924 | _T_21670; // @[Mux.scala 27:72]
  wire  _T_21118 = bht_rd_addr_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_21671 = _T_21118 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21926 = _T_21925 | _T_21671; // @[Mux.scala 27:72]
  wire  _T_21121 = bht_rd_addr_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_21672 = _T_21121 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21927 = _T_21926 | _T_21672; // @[Mux.scala 27:72]
  wire  _T_21124 = bht_rd_addr_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_21673 = _T_21124 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21928 = _T_21927 | _T_21673; // @[Mux.scala 27:72]
  wire  _T_21127 = bht_rd_addr_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_21674 = _T_21127 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21929 = _T_21928 | _T_21674; // @[Mux.scala 27:72]
  wire  _T_21130 = bht_rd_addr_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_21675 = _T_21130 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21930 = _T_21929 | _T_21675; // @[Mux.scala 27:72]
  wire  _T_21133 = bht_rd_addr_f == 8'h70; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_21676 = _T_21133 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21931 = _T_21930 | _T_21676; // @[Mux.scala 27:72]
  wire  _T_21136 = bht_rd_addr_f == 8'h71; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_21677 = _T_21136 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21932 = _T_21931 | _T_21677; // @[Mux.scala 27:72]
  wire  _T_21139 = bht_rd_addr_f == 8'h72; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_21678 = _T_21139 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21933 = _T_21932 | _T_21678; // @[Mux.scala 27:72]
  wire  _T_21142 = bht_rd_addr_f == 8'h73; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_21679 = _T_21142 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21934 = _T_21933 | _T_21679; // @[Mux.scala 27:72]
  wire  _T_21145 = bht_rd_addr_f == 8'h74; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_21680 = _T_21145 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21935 = _T_21934 | _T_21680; // @[Mux.scala 27:72]
  wire  _T_21148 = bht_rd_addr_f == 8'h75; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_21681 = _T_21148 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21936 = _T_21935 | _T_21681; // @[Mux.scala 27:72]
  wire  _T_21151 = bht_rd_addr_f == 8'h76; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_21682 = _T_21151 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21937 = _T_21936 | _T_21682; // @[Mux.scala 27:72]
  wire  _T_21154 = bht_rd_addr_f == 8'h77; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_21683 = _T_21154 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21938 = _T_21937 | _T_21683; // @[Mux.scala 27:72]
  wire  _T_21157 = bht_rd_addr_f == 8'h78; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_21684 = _T_21157 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21939 = _T_21938 | _T_21684; // @[Mux.scala 27:72]
  wire  _T_21160 = bht_rd_addr_f == 8'h79; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_21685 = _T_21160 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21940 = _T_21939 | _T_21685; // @[Mux.scala 27:72]
  wire  _T_21163 = bht_rd_addr_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_21686 = _T_21163 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21941 = _T_21940 | _T_21686; // @[Mux.scala 27:72]
  wire  _T_21166 = bht_rd_addr_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_21687 = _T_21166 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21942 = _T_21941 | _T_21687; // @[Mux.scala 27:72]
  wire  _T_21169 = bht_rd_addr_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_21688 = _T_21169 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21943 = _T_21942 | _T_21688; // @[Mux.scala 27:72]
  wire  _T_21172 = bht_rd_addr_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_21689 = _T_21172 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21944 = _T_21943 | _T_21689; // @[Mux.scala 27:72]
  wire  _T_21175 = bht_rd_addr_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_21690 = _T_21175 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21945 = _T_21944 | _T_21690; // @[Mux.scala 27:72]
  wire  _T_21178 = bht_rd_addr_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_21691 = _T_21178 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21946 = _T_21945 | _T_21691; // @[Mux.scala 27:72]
  wire  _T_21181 = bht_rd_addr_f == 8'h80; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_21692 = _T_21181 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21947 = _T_21946 | _T_21692; // @[Mux.scala 27:72]
  wire  _T_21184 = bht_rd_addr_f == 8'h81; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_21693 = _T_21184 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21948 = _T_21947 | _T_21693; // @[Mux.scala 27:72]
  wire  _T_21187 = bht_rd_addr_f == 8'h82; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_21694 = _T_21187 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21949 = _T_21948 | _T_21694; // @[Mux.scala 27:72]
  wire  _T_21190 = bht_rd_addr_f == 8'h83; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_21695 = _T_21190 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21950 = _T_21949 | _T_21695; // @[Mux.scala 27:72]
  wire  _T_21193 = bht_rd_addr_f == 8'h84; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_21696 = _T_21193 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21951 = _T_21950 | _T_21696; // @[Mux.scala 27:72]
  wire  _T_21196 = bht_rd_addr_f == 8'h85; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_21697 = _T_21196 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21952 = _T_21951 | _T_21697; // @[Mux.scala 27:72]
  wire  _T_21199 = bht_rd_addr_f == 8'h86; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_21698 = _T_21199 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21953 = _T_21952 | _T_21698; // @[Mux.scala 27:72]
  wire  _T_21202 = bht_rd_addr_f == 8'h87; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_21699 = _T_21202 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21954 = _T_21953 | _T_21699; // @[Mux.scala 27:72]
  wire  _T_21205 = bht_rd_addr_f == 8'h88; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_21700 = _T_21205 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21955 = _T_21954 | _T_21700; // @[Mux.scala 27:72]
  wire  _T_21208 = bht_rd_addr_f == 8'h89; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_21701 = _T_21208 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21956 = _T_21955 | _T_21701; // @[Mux.scala 27:72]
  wire  _T_21211 = bht_rd_addr_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_21702 = _T_21211 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21957 = _T_21956 | _T_21702; // @[Mux.scala 27:72]
  wire  _T_21214 = bht_rd_addr_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_21703 = _T_21214 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21958 = _T_21957 | _T_21703; // @[Mux.scala 27:72]
  wire  _T_21217 = bht_rd_addr_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_21704 = _T_21217 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21959 = _T_21958 | _T_21704; // @[Mux.scala 27:72]
  wire  _T_21220 = bht_rd_addr_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_21705 = _T_21220 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21960 = _T_21959 | _T_21705; // @[Mux.scala 27:72]
  wire  _T_21223 = bht_rd_addr_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_21706 = _T_21223 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21961 = _T_21960 | _T_21706; // @[Mux.scala 27:72]
  wire  _T_21226 = bht_rd_addr_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_21707 = _T_21226 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21962 = _T_21961 | _T_21707; // @[Mux.scala 27:72]
  wire  _T_21229 = bht_rd_addr_f == 8'h90; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_21708 = _T_21229 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21963 = _T_21962 | _T_21708; // @[Mux.scala 27:72]
  wire  _T_21232 = bht_rd_addr_f == 8'h91; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_21709 = _T_21232 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21964 = _T_21963 | _T_21709; // @[Mux.scala 27:72]
  wire  _T_21235 = bht_rd_addr_f == 8'h92; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_21710 = _T_21235 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21965 = _T_21964 | _T_21710; // @[Mux.scala 27:72]
  wire  _T_21238 = bht_rd_addr_f == 8'h93; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_21711 = _T_21238 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21966 = _T_21965 | _T_21711; // @[Mux.scala 27:72]
  wire  _T_21241 = bht_rd_addr_f == 8'h94; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_21712 = _T_21241 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21967 = _T_21966 | _T_21712; // @[Mux.scala 27:72]
  wire  _T_21244 = bht_rd_addr_f == 8'h95; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_21713 = _T_21244 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21968 = _T_21967 | _T_21713; // @[Mux.scala 27:72]
  wire  _T_21247 = bht_rd_addr_f == 8'h96; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_21714 = _T_21247 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21969 = _T_21968 | _T_21714; // @[Mux.scala 27:72]
  wire  _T_21250 = bht_rd_addr_f == 8'h97; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_21715 = _T_21250 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21970 = _T_21969 | _T_21715; // @[Mux.scala 27:72]
  wire  _T_21253 = bht_rd_addr_f == 8'h98; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_21716 = _T_21253 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21971 = _T_21970 | _T_21716; // @[Mux.scala 27:72]
  wire  _T_21256 = bht_rd_addr_f == 8'h99; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_21717 = _T_21256 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21972 = _T_21971 | _T_21717; // @[Mux.scala 27:72]
  wire  _T_21259 = bht_rd_addr_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_21718 = _T_21259 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21973 = _T_21972 | _T_21718; // @[Mux.scala 27:72]
  wire  _T_21262 = bht_rd_addr_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_21719 = _T_21262 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21974 = _T_21973 | _T_21719; // @[Mux.scala 27:72]
  wire  _T_21265 = bht_rd_addr_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_21720 = _T_21265 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21975 = _T_21974 | _T_21720; // @[Mux.scala 27:72]
  wire  _T_21268 = bht_rd_addr_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_21721 = _T_21268 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21976 = _T_21975 | _T_21721; // @[Mux.scala 27:72]
  wire  _T_21271 = bht_rd_addr_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_21722 = _T_21271 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21977 = _T_21976 | _T_21722; // @[Mux.scala 27:72]
  wire  _T_21274 = bht_rd_addr_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_21723 = _T_21274 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21978 = _T_21977 | _T_21723; // @[Mux.scala 27:72]
  wire  _T_21277 = bht_rd_addr_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_21724 = _T_21277 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21979 = _T_21978 | _T_21724; // @[Mux.scala 27:72]
  wire  _T_21280 = bht_rd_addr_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_21725 = _T_21280 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21980 = _T_21979 | _T_21725; // @[Mux.scala 27:72]
  wire  _T_21283 = bht_rd_addr_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_21726 = _T_21283 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21981 = _T_21980 | _T_21726; // @[Mux.scala 27:72]
  wire  _T_21286 = bht_rd_addr_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_21727 = _T_21286 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21982 = _T_21981 | _T_21727; // @[Mux.scala 27:72]
  wire  _T_21289 = bht_rd_addr_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_21728 = _T_21289 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21983 = _T_21982 | _T_21728; // @[Mux.scala 27:72]
  wire  _T_21292 = bht_rd_addr_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_21729 = _T_21292 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21984 = _T_21983 | _T_21729; // @[Mux.scala 27:72]
  wire  _T_21295 = bht_rd_addr_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_21730 = _T_21295 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21985 = _T_21984 | _T_21730; // @[Mux.scala 27:72]
  wire  _T_21298 = bht_rd_addr_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_21731 = _T_21298 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21986 = _T_21985 | _T_21731; // @[Mux.scala 27:72]
  wire  _T_21301 = bht_rd_addr_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_21732 = _T_21301 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21987 = _T_21986 | _T_21732; // @[Mux.scala 27:72]
  wire  _T_21304 = bht_rd_addr_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_21733 = _T_21304 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21988 = _T_21987 | _T_21733; // @[Mux.scala 27:72]
  wire  _T_21307 = bht_rd_addr_f == 8'haa; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_21734 = _T_21307 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21989 = _T_21988 | _T_21734; // @[Mux.scala 27:72]
  wire  _T_21310 = bht_rd_addr_f == 8'hab; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_21735 = _T_21310 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21990 = _T_21989 | _T_21735; // @[Mux.scala 27:72]
  wire  _T_21313 = bht_rd_addr_f == 8'hac; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_21736 = _T_21313 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21991 = _T_21990 | _T_21736; // @[Mux.scala 27:72]
  wire  _T_21316 = bht_rd_addr_f == 8'had; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_21737 = _T_21316 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21992 = _T_21991 | _T_21737; // @[Mux.scala 27:72]
  wire  _T_21319 = bht_rd_addr_f == 8'hae; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_21738 = _T_21319 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21993 = _T_21992 | _T_21738; // @[Mux.scala 27:72]
  wire  _T_21322 = bht_rd_addr_f == 8'haf; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_21739 = _T_21322 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21994 = _T_21993 | _T_21739; // @[Mux.scala 27:72]
  wire  _T_21325 = bht_rd_addr_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_21740 = _T_21325 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21995 = _T_21994 | _T_21740; // @[Mux.scala 27:72]
  wire  _T_21328 = bht_rd_addr_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_21741 = _T_21328 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21996 = _T_21995 | _T_21741; // @[Mux.scala 27:72]
  wire  _T_21331 = bht_rd_addr_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_21742 = _T_21331 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21997 = _T_21996 | _T_21742; // @[Mux.scala 27:72]
  wire  _T_21334 = bht_rd_addr_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_21743 = _T_21334 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21998 = _T_21997 | _T_21743; // @[Mux.scala 27:72]
  wire  _T_21337 = bht_rd_addr_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_21744 = _T_21337 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21999 = _T_21998 | _T_21744; // @[Mux.scala 27:72]
  wire  _T_21340 = bht_rd_addr_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_21745 = _T_21340 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22000 = _T_21999 | _T_21745; // @[Mux.scala 27:72]
  wire  _T_21343 = bht_rd_addr_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_21746 = _T_21343 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22001 = _T_22000 | _T_21746; // @[Mux.scala 27:72]
  wire  _T_21346 = bht_rd_addr_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_21747 = _T_21346 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22002 = _T_22001 | _T_21747; // @[Mux.scala 27:72]
  wire  _T_21349 = bht_rd_addr_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_21748 = _T_21349 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22003 = _T_22002 | _T_21748; // @[Mux.scala 27:72]
  wire  _T_21352 = bht_rd_addr_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_21749 = _T_21352 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22004 = _T_22003 | _T_21749; // @[Mux.scala 27:72]
  wire  _T_21355 = bht_rd_addr_f == 8'hba; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_21750 = _T_21355 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22005 = _T_22004 | _T_21750; // @[Mux.scala 27:72]
  wire  _T_21358 = bht_rd_addr_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_21751 = _T_21358 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22006 = _T_22005 | _T_21751; // @[Mux.scala 27:72]
  wire  _T_21361 = bht_rd_addr_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_21752 = _T_21361 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22007 = _T_22006 | _T_21752; // @[Mux.scala 27:72]
  wire  _T_21364 = bht_rd_addr_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_21753 = _T_21364 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22008 = _T_22007 | _T_21753; // @[Mux.scala 27:72]
  wire  _T_21367 = bht_rd_addr_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_21754 = _T_21367 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22009 = _T_22008 | _T_21754; // @[Mux.scala 27:72]
  wire  _T_21370 = bht_rd_addr_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_21755 = _T_21370 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22010 = _T_22009 | _T_21755; // @[Mux.scala 27:72]
  wire  _T_21373 = bht_rd_addr_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_21756 = _T_21373 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22011 = _T_22010 | _T_21756; // @[Mux.scala 27:72]
  wire  _T_21376 = bht_rd_addr_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_21757 = _T_21376 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22012 = _T_22011 | _T_21757; // @[Mux.scala 27:72]
  wire  _T_21379 = bht_rd_addr_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_21758 = _T_21379 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22013 = _T_22012 | _T_21758; // @[Mux.scala 27:72]
  wire  _T_21382 = bht_rd_addr_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_21759 = _T_21382 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22014 = _T_22013 | _T_21759; // @[Mux.scala 27:72]
  wire  _T_21385 = bht_rd_addr_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_21760 = _T_21385 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22015 = _T_22014 | _T_21760; // @[Mux.scala 27:72]
  wire  _T_21388 = bht_rd_addr_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_21761 = _T_21388 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22016 = _T_22015 | _T_21761; // @[Mux.scala 27:72]
  wire  _T_21391 = bht_rd_addr_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_21762 = _T_21391 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22017 = _T_22016 | _T_21762; // @[Mux.scala 27:72]
  wire  _T_21394 = bht_rd_addr_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_21763 = _T_21394 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22018 = _T_22017 | _T_21763; // @[Mux.scala 27:72]
  wire  _T_21397 = bht_rd_addr_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_21764 = _T_21397 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22019 = _T_22018 | _T_21764; // @[Mux.scala 27:72]
  wire  _T_21400 = bht_rd_addr_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_21765 = _T_21400 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22020 = _T_22019 | _T_21765; // @[Mux.scala 27:72]
  wire  _T_21403 = bht_rd_addr_f == 8'hca; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_21766 = _T_21403 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22021 = _T_22020 | _T_21766; // @[Mux.scala 27:72]
  wire  _T_21406 = bht_rd_addr_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_21767 = _T_21406 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22022 = _T_22021 | _T_21767; // @[Mux.scala 27:72]
  wire  _T_21409 = bht_rd_addr_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_21768 = _T_21409 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22023 = _T_22022 | _T_21768; // @[Mux.scala 27:72]
  wire  _T_21412 = bht_rd_addr_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_21769 = _T_21412 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22024 = _T_22023 | _T_21769; // @[Mux.scala 27:72]
  wire  _T_21415 = bht_rd_addr_f == 8'hce; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_21770 = _T_21415 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22025 = _T_22024 | _T_21770; // @[Mux.scala 27:72]
  wire  _T_21418 = bht_rd_addr_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_21771 = _T_21418 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22026 = _T_22025 | _T_21771; // @[Mux.scala 27:72]
  wire  _T_21421 = bht_rd_addr_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_21772 = _T_21421 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22027 = _T_22026 | _T_21772; // @[Mux.scala 27:72]
  wire  _T_21424 = bht_rd_addr_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_21773 = _T_21424 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22028 = _T_22027 | _T_21773; // @[Mux.scala 27:72]
  wire  _T_21427 = bht_rd_addr_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_21774 = _T_21427 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22029 = _T_22028 | _T_21774; // @[Mux.scala 27:72]
  wire  _T_21430 = bht_rd_addr_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_21775 = _T_21430 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22030 = _T_22029 | _T_21775; // @[Mux.scala 27:72]
  wire  _T_21433 = bht_rd_addr_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_21776 = _T_21433 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22031 = _T_22030 | _T_21776; // @[Mux.scala 27:72]
  wire  _T_21436 = bht_rd_addr_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_21777 = _T_21436 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22032 = _T_22031 | _T_21777; // @[Mux.scala 27:72]
  wire  _T_21439 = bht_rd_addr_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_21778 = _T_21439 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22033 = _T_22032 | _T_21778; // @[Mux.scala 27:72]
  wire  _T_21442 = bht_rd_addr_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_21779 = _T_21442 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22034 = _T_22033 | _T_21779; // @[Mux.scala 27:72]
  wire  _T_21445 = bht_rd_addr_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_21780 = _T_21445 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22035 = _T_22034 | _T_21780; // @[Mux.scala 27:72]
  wire  _T_21448 = bht_rd_addr_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_21781 = _T_21448 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22036 = _T_22035 | _T_21781; // @[Mux.scala 27:72]
  wire  _T_21451 = bht_rd_addr_f == 8'hda; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_21782 = _T_21451 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22037 = _T_22036 | _T_21782; // @[Mux.scala 27:72]
  wire  _T_21454 = bht_rd_addr_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_21783 = _T_21454 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22038 = _T_22037 | _T_21783; // @[Mux.scala 27:72]
  wire  _T_21457 = bht_rd_addr_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_21784 = _T_21457 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22039 = _T_22038 | _T_21784; // @[Mux.scala 27:72]
  wire  _T_21460 = bht_rd_addr_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_21785 = _T_21460 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22040 = _T_22039 | _T_21785; // @[Mux.scala 27:72]
  wire  _T_21463 = bht_rd_addr_f == 8'hde; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_21786 = _T_21463 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22041 = _T_22040 | _T_21786; // @[Mux.scala 27:72]
  wire  _T_21466 = bht_rd_addr_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_21787 = _T_21466 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22042 = _T_22041 | _T_21787; // @[Mux.scala 27:72]
  wire  _T_21469 = bht_rd_addr_f == 8'he0; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_21788 = _T_21469 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22043 = _T_22042 | _T_21788; // @[Mux.scala 27:72]
  wire  _T_21472 = bht_rd_addr_f == 8'he1; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_21789 = _T_21472 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22044 = _T_22043 | _T_21789; // @[Mux.scala 27:72]
  wire  _T_21475 = bht_rd_addr_f == 8'he2; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_21790 = _T_21475 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22045 = _T_22044 | _T_21790; // @[Mux.scala 27:72]
  wire  _T_21478 = bht_rd_addr_f == 8'he3; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_21791 = _T_21478 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22046 = _T_22045 | _T_21791; // @[Mux.scala 27:72]
  wire  _T_21481 = bht_rd_addr_f == 8'he4; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_21792 = _T_21481 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22047 = _T_22046 | _T_21792; // @[Mux.scala 27:72]
  wire  _T_21484 = bht_rd_addr_f == 8'he5; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_21793 = _T_21484 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22048 = _T_22047 | _T_21793; // @[Mux.scala 27:72]
  wire  _T_21487 = bht_rd_addr_f == 8'he6; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_21794 = _T_21487 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22049 = _T_22048 | _T_21794; // @[Mux.scala 27:72]
  wire  _T_21490 = bht_rd_addr_f == 8'he7; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_21795 = _T_21490 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22050 = _T_22049 | _T_21795; // @[Mux.scala 27:72]
  wire  _T_21493 = bht_rd_addr_f == 8'he8; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_21796 = _T_21493 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22051 = _T_22050 | _T_21796; // @[Mux.scala 27:72]
  wire  _T_21496 = bht_rd_addr_f == 8'he9; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_21797 = _T_21496 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22052 = _T_22051 | _T_21797; // @[Mux.scala 27:72]
  wire  _T_21499 = bht_rd_addr_f == 8'hea; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_21798 = _T_21499 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22053 = _T_22052 | _T_21798; // @[Mux.scala 27:72]
  wire  _T_21502 = bht_rd_addr_f == 8'heb; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_21799 = _T_21502 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22054 = _T_22053 | _T_21799; // @[Mux.scala 27:72]
  wire  _T_21505 = bht_rd_addr_f == 8'hec; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_21800 = _T_21505 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22055 = _T_22054 | _T_21800; // @[Mux.scala 27:72]
  wire  _T_21508 = bht_rd_addr_f == 8'hed; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_21801 = _T_21508 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22056 = _T_22055 | _T_21801; // @[Mux.scala 27:72]
  wire  _T_21511 = bht_rd_addr_f == 8'hee; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_21802 = _T_21511 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22057 = _T_22056 | _T_21802; // @[Mux.scala 27:72]
  wire  _T_21514 = bht_rd_addr_f == 8'hef; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_21803 = _T_21514 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22058 = _T_22057 | _T_21803; // @[Mux.scala 27:72]
  wire  _T_21517 = bht_rd_addr_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_21804 = _T_21517 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22059 = _T_22058 | _T_21804; // @[Mux.scala 27:72]
  wire  _T_21520 = bht_rd_addr_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_21805 = _T_21520 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22060 = _T_22059 | _T_21805; // @[Mux.scala 27:72]
  wire  _T_21523 = bht_rd_addr_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_21806 = _T_21523 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22061 = _T_22060 | _T_21806; // @[Mux.scala 27:72]
  wire  _T_21526 = bht_rd_addr_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_21807 = _T_21526 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22062 = _T_22061 | _T_21807; // @[Mux.scala 27:72]
  wire  _T_21529 = bht_rd_addr_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_21808 = _T_21529 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22063 = _T_22062 | _T_21808; // @[Mux.scala 27:72]
  wire  _T_21532 = bht_rd_addr_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_21809 = _T_21532 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22064 = _T_22063 | _T_21809; // @[Mux.scala 27:72]
  wire  _T_21535 = bht_rd_addr_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_21810 = _T_21535 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22065 = _T_22064 | _T_21810; // @[Mux.scala 27:72]
  wire  _T_21538 = bht_rd_addr_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_21811 = _T_21538 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22066 = _T_22065 | _T_21811; // @[Mux.scala 27:72]
  wire  _T_21541 = bht_rd_addr_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_21812 = _T_21541 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22067 = _T_22066 | _T_21812; // @[Mux.scala 27:72]
  wire  _T_21544 = bht_rd_addr_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_21813 = _T_21544 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22068 = _T_22067 | _T_21813; // @[Mux.scala 27:72]
  wire  _T_21547 = bht_rd_addr_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_21814 = _T_21547 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22069 = _T_22068 | _T_21814; // @[Mux.scala 27:72]
  wire  _T_21550 = bht_rd_addr_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_21815 = _T_21550 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22070 = _T_22069 | _T_21815; // @[Mux.scala 27:72]
  wire  _T_21553 = bht_rd_addr_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_21816 = _T_21553 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22071 = _T_22070 | _T_21816; // @[Mux.scala 27:72]
  wire  _T_21556 = bht_rd_addr_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_21817 = _T_21556 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22072 = _T_22071 | _T_21817; // @[Mux.scala 27:72]
  wire  _T_21559 = bht_rd_addr_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_21818 = _T_21559 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22073 = _T_22072 | _T_21818; // @[Mux.scala 27:72]
  wire  _T_21562 = bht_rd_addr_f == 8'hff; // @[el2_ifu_bp_ctl.scala 388:106]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_21819 = _T_21562 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_22073 | _T_21819; // @[Mux.scala 27:72]
  wire [1:0] _T_258 = _T_143 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_569 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_569[9:2] ^ fghr; // @[el2_lib.scala 188:35]
  wire  _T_22077 = bht_rd_addr_hashed_p1_f == 8'h0; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22844 = _T_22077 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22080 = bht_rd_addr_hashed_p1_f == 8'h1; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22845 = _T_22080 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23100 = _T_22844 | _T_22845; // @[Mux.scala 27:72]
  wire  _T_22083 = bht_rd_addr_hashed_p1_f == 8'h2; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22846 = _T_22083 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23101 = _T_23100 | _T_22846; // @[Mux.scala 27:72]
  wire  _T_22086 = bht_rd_addr_hashed_p1_f == 8'h3; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22847 = _T_22086 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23102 = _T_23101 | _T_22847; // @[Mux.scala 27:72]
  wire  _T_22089 = bht_rd_addr_hashed_p1_f == 8'h4; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22848 = _T_22089 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23103 = _T_23102 | _T_22848; // @[Mux.scala 27:72]
  wire  _T_22092 = bht_rd_addr_hashed_p1_f == 8'h5; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22849 = _T_22092 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23104 = _T_23103 | _T_22849; // @[Mux.scala 27:72]
  wire  _T_22095 = bht_rd_addr_hashed_p1_f == 8'h6; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22850 = _T_22095 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23105 = _T_23104 | _T_22850; // @[Mux.scala 27:72]
  wire  _T_22098 = bht_rd_addr_hashed_p1_f == 8'h7; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22851 = _T_22098 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23106 = _T_23105 | _T_22851; // @[Mux.scala 27:72]
  wire  _T_22101 = bht_rd_addr_hashed_p1_f == 8'h8; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22852 = _T_22101 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23107 = _T_23106 | _T_22852; // @[Mux.scala 27:72]
  wire  _T_22104 = bht_rd_addr_hashed_p1_f == 8'h9; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22853 = _T_22104 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23108 = _T_23107 | _T_22853; // @[Mux.scala 27:72]
  wire  _T_22107 = bht_rd_addr_hashed_p1_f == 8'ha; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22854 = _T_22107 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23109 = _T_23108 | _T_22854; // @[Mux.scala 27:72]
  wire  _T_22110 = bht_rd_addr_hashed_p1_f == 8'hb; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22855 = _T_22110 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23110 = _T_23109 | _T_22855; // @[Mux.scala 27:72]
  wire  _T_22113 = bht_rd_addr_hashed_p1_f == 8'hc; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22856 = _T_22113 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23111 = _T_23110 | _T_22856; // @[Mux.scala 27:72]
  wire  _T_22116 = bht_rd_addr_hashed_p1_f == 8'hd; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22857 = _T_22116 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23112 = _T_23111 | _T_22857; // @[Mux.scala 27:72]
  wire  _T_22119 = bht_rd_addr_hashed_p1_f == 8'he; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22858 = _T_22119 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23113 = _T_23112 | _T_22858; // @[Mux.scala 27:72]
  wire  _T_22122 = bht_rd_addr_hashed_p1_f == 8'hf; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22859 = _T_22122 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23114 = _T_23113 | _T_22859; // @[Mux.scala 27:72]
  wire  _T_22125 = bht_rd_addr_hashed_p1_f == 8'h10; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22860 = _T_22125 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23115 = _T_23114 | _T_22860; // @[Mux.scala 27:72]
  wire  _T_22128 = bht_rd_addr_hashed_p1_f == 8'h11; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22861 = _T_22128 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23116 = _T_23115 | _T_22861; // @[Mux.scala 27:72]
  wire  _T_22131 = bht_rd_addr_hashed_p1_f == 8'h12; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22862 = _T_22131 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23117 = _T_23116 | _T_22862; // @[Mux.scala 27:72]
  wire  _T_22134 = bht_rd_addr_hashed_p1_f == 8'h13; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22863 = _T_22134 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23118 = _T_23117 | _T_22863; // @[Mux.scala 27:72]
  wire  _T_22137 = bht_rd_addr_hashed_p1_f == 8'h14; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22864 = _T_22137 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23119 = _T_23118 | _T_22864; // @[Mux.scala 27:72]
  wire  _T_22140 = bht_rd_addr_hashed_p1_f == 8'h15; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22865 = _T_22140 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23120 = _T_23119 | _T_22865; // @[Mux.scala 27:72]
  wire  _T_22143 = bht_rd_addr_hashed_p1_f == 8'h16; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22866 = _T_22143 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23121 = _T_23120 | _T_22866; // @[Mux.scala 27:72]
  wire  _T_22146 = bht_rd_addr_hashed_p1_f == 8'h17; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22867 = _T_22146 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23122 = _T_23121 | _T_22867; // @[Mux.scala 27:72]
  wire  _T_22149 = bht_rd_addr_hashed_p1_f == 8'h18; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22868 = _T_22149 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23123 = _T_23122 | _T_22868; // @[Mux.scala 27:72]
  wire  _T_22152 = bht_rd_addr_hashed_p1_f == 8'h19; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22869 = _T_22152 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23124 = _T_23123 | _T_22869; // @[Mux.scala 27:72]
  wire  _T_22155 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22870 = _T_22155 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23125 = _T_23124 | _T_22870; // @[Mux.scala 27:72]
  wire  _T_22158 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22871 = _T_22158 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23126 = _T_23125 | _T_22871; // @[Mux.scala 27:72]
  wire  _T_22161 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22872 = _T_22161 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23127 = _T_23126 | _T_22872; // @[Mux.scala 27:72]
  wire  _T_22164 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22873 = _T_22164 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23128 = _T_23127 | _T_22873; // @[Mux.scala 27:72]
  wire  _T_22167 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22874 = _T_22167 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23129 = _T_23128 | _T_22874; // @[Mux.scala 27:72]
  wire  _T_22170 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22875 = _T_22170 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23130 = _T_23129 | _T_22875; // @[Mux.scala 27:72]
  wire  _T_22173 = bht_rd_addr_hashed_p1_f == 8'h20; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22876 = _T_22173 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23131 = _T_23130 | _T_22876; // @[Mux.scala 27:72]
  wire  _T_22176 = bht_rd_addr_hashed_p1_f == 8'h21; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22877 = _T_22176 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23132 = _T_23131 | _T_22877; // @[Mux.scala 27:72]
  wire  _T_22179 = bht_rd_addr_hashed_p1_f == 8'h22; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22878 = _T_22179 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23133 = _T_23132 | _T_22878; // @[Mux.scala 27:72]
  wire  _T_22182 = bht_rd_addr_hashed_p1_f == 8'h23; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22879 = _T_22182 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23134 = _T_23133 | _T_22879; // @[Mux.scala 27:72]
  wire  _T_22185 = bht_rd_addr_hashed_p1_f == 8'h24; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22880 = _T_22185 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23135 = _T_23134 | _T_22880; // @[Mux.scala 27:72]
  wire  _T_22188 = bht_rd_addr_hashed_p1_f == 8'h25; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22881 = _T_22188 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23136 = _T_23135 | _T_22881; // @[Mux.scala 27:72]
  wire  _T_22191 = bht_rd_addr_hashed_p1_f == 8'h26; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22882 = _T_22191 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23137 = _T_23136 | _T_22882; // @[Mux.scala 27:72]
  wire  _T_22194 = bht_rd_addr_hashed_p1_f == 8'h27; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22883 = _T_22194 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23138 = _T_23137 | _T_22883; // @[Mux.scala 27:72]
  wire  _T_22197 = bht_rd_addr_hashed_p1_f == 8'h28; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22884 = _T_22197 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23139 = _T_23138 | _T_22884; // @[Mux.scala 27:72]
  wire  _T_22200 = bht_rd_addr_hashed_p1_f == 8'h29; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22885 = _T_22200 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23140 = _T_23139 | _T_22885; // @[Mux.scala 27:72]
  wire  _T_22203 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22886 = _T_22203 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23141 = _T_23140 | _T_22886; // @[Mux.scala 27:72]
  wire  _T_22206 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22887 = _T_22206 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23142 = _T_23141 | _T_22887; // @[Mux.scala 27:72]
  wire  _T_22209 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22888 = _T_22209 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23143 = _T_23142 | _T_22888; // @[Mux.scala 27:72]
  wire  _T_22212 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22889 = _T_22212 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23144 = _T_23143 | _T_22889; // @[Mux.scala 27:72]
  wire  _T_22215 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22890 = _T_22215 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23145 = _T_23144 | _T_22890; // @[Mux.scala 27:72]
  wire  _T_22218 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22891 = _T_22218 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23146 = _T_23145 | _T_22891; // @[Mux.scala 27:72]
  wire  _T_22221 = bht_rd_addr_hashed_p1_f == 8'h30; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22892 = _T_22221 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23147 = _T_23146 | _T_22892; // @[Mux.scala 27:72]
  wire  _T_22224 = bht_rd_addr_hashed_p1_f == 8'h31; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22893 = _T_22224 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23148 = _T_23147 | _T_22893; // @[Mux.scala 27:72]
  wire  _T_22227 = bht_rd_addr_hashed_p1_f == 8'h32; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22894 = _T_22227 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23149 = _T_23148 | _T_22894; // @[Mux.scala 27:72]
  wire  _T_22230 = bht_rd_addr_hashed_p1_f == 8'h33; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22895 = _T_22230 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23150 = _T_23149 | _T_22895; // @[Mux.scala 27:72]
  wire  _T_22233 = bht_rd_addr_hashed_p1_f == 8'h34; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22896 = _T_22233 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23151 = _T_23150 | _T_22896; // @[Mux.scala 27:72]
  wire  _T_22236 = bht_rd_addr_hashed_p1_f == 8'h35; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22897 = _T_22236 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23152 = _T_23151 | _T_22897; // @[Mux.scala 27:72]
  wire  _T_22239 = bht_rd_addr_hashed_p1_f == 8'h36; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22898 = _T_22239 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23153 = _T_23152 | _T_22898; // @[Mux.scala 27:72]
  wire  _T_22242 = bht_rd_addr_hashed_p1_f == 8'h37; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22899 = _T_22242 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23154 = _T_23153 | _T_22899; // @[Mux.scala 27:72]
  wire  _T_22245 = bht_rd_addr_hashed_p1_f == 8'h38; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22900 = _T_22245 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23155 = _T_23154 | _T_22900; // @[Mux.scala 27:72]
  wire  _T_22248 = bht_rd_addr_hashed_p1_f == 8'h39; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22901 = _T_22248 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23156 = _T_23155 | _T_22901; // @[Mux.scala 27:72]
  wire  _T_22251 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22902 = _T_22251 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23157 = _T_23156 | _T_22902; // @[Mux.scala 27:72]
  wire  _T_22254 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22903 = _T_22254 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23158 = _T_23157 | _T_22903; // @[Mux.scala 27:72]
  wire  _T_22257 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22904 = _T_22257 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23159 = _T_23158 | _T_22904; // @[Mux.scala 27:72]
  wire  _T_22260 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22905 = _T_22260 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23160 = _T_23159 | _T_22905; // @[Mux.scala 27:72]
  wire  _T_22263 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22906 = _T_22263 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23161 = _T_23160 | _T_22906; // @[Mux.scala 27:72]
  wire  _T_22266 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22907 = _T_22266 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23162 = _T_23161 | _T_22907; // @[Mux.scala 27:72]
  wire  _T_22269 = bht_rd_addr_hashed_p1_f == 8'h40; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22908 = _T_22269 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23163 = _T_23162 | _T_22908; // @[Mux.scala 27:72]
  wire  _T_22272 = bht_rd_addr_hashed_p1_f == 8'h41; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22909 = _T_22272 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23164 = _T_23163 | _T_22909; // @[Mux.scala 27:72]
  wire  _T_22275 = bht_rd_addr_hashed_p1_f == 8'h42; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22910 = _T_22275 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23165 = _T_23164 | _T_22910; // @[Mux.scala 27:72]
  wire  _T_22278 = bht_rd_addr_hashed_p1_f == 8'h43; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22911 = _T_22278 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23166 = _T_23165 | _T_22911; // @[Mux.scala 27:72]
  wire  _T_22281 = bht_rd_addr_hashed_p1_f == 8'h44; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22912 = _T_22281 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23167 = _T_23166 | _T_22912; // @[Mux.scala 27:72]
  wire  _T_22284 = bht_rd_addr_hashed_p1_f == 8'h45; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22913 = _T_22284 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23168 = _T_23167 | _T_22913; // @[Mux.scala 27:72]
  wire  _T_22287 = bht_rd_addr_hashed_p1_f == 8'h46; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22914 = _T_22287 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23169 = _T_23168 | _T_22914; // @[Mux.scala 27:72]
  wire  _T_22290 = bht_rd_addr_hashed_p1_f == 8'h47; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22915 = _T_22290 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23170 = _T_23169 | _T_22915; // @[Mux.scala 27:72]
  wire  _T_22293 = bht_rd_addr_hashed_p1_f == 8'h48; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22916 = _T_22293 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23171 = _T_23170 | _T_22916; // @[Mux.scala 27:72]
  wire  _T_22296 = bht_rd_addr_hashed_p1_f == 8'h49; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22917 = _T_22296 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23172 = _T_23171 | _T_22917; // @[Mux.scala 27:72]
  wire  _T_22299 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22918 = _T_22299 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23173 = _T_23172 | _T_22918; // @[Mux.scala 27:72]
  wire  _T_22302 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22919 = _T_22302 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23174 = _T_23173 | _T_22919; // @[Mux.scala 27:72]
  wire  _T_22305 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22920 = _T_22305 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23175 = _T_23174 | _T_22920; // @[Mux.scala 27:72]
  wire  _T_22308 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22921 = _T_22308 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23176 = _T_23175 | _T_22921; // @[Mux.scala 27:72]
  wire  _T_22311 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22922 = _T_22311 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23177 = _T_23176 | _T_22922; // @[Mux.scala 27:72]
  wire  _T_22314 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22923 = _T_22314 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23178 = _T_23177 | _T_22923; // @[Mux.scala 27:72]
  wire  _T_22317 = bht_rd_addr_hashed_p1_f == 8'h50; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22924 = _T_22317 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23179 = _T_23178 | _T_22924; // @[Mux.scala 27:72]
  wire  _T_22320 = bht_rd_addr_hashed_p1_f == 8'h51; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22925 = _T_22320 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23180 = _T_23179 | _T_22925; // @[Mux.scala 27:72]
  wire  _T_22323 = bht_rd_addr_hashed_p1_f == 8'h52; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22926 = _T_22323 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23181 = _T_23180 | _T_22926; // @[Mux.scala 27:72]
  wire  _T_22326 = bht_rd_addr_hashed_p1_f == 8'h53; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22927 = _T_22326 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23182 = _T_23181 | _T_22927; // @[Mux.scala 27:72]
  wire  _T_22329 = bht_rd_addr_hashed_p1_f == 8'h54; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22928 = _T_22329 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23183 = _T_23182 | _T_22928; // @[Mux.scala 27:72]
  wire  _T_22332 = bht_rd_addr_hashed_p1_f == 8'h55; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22929 = _T_22332 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23184 = _T_23183 | _T_22929; // @[Mux.scala 27:72]
  wire  _T_22335 = bht_rd_addr_hashed_p1_f == 8'h56; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22930 = _T_22335 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23185 = _T_23184 | _T_22930; // @[Mux.scala 27:72]
  wire  _T_22338 = bht_rd_addr_hashed_p1_f == 8'h57; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22931 = _T_22338 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23186 = _T_23185 | _T_22931; // @[Mux.scala 27:72]
  wire  _T_22341 = bht_rd_addr_hashed_p1_f == 8'h58; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22932 = _T_22341 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23187 = _T_23186 | _T_22932; // @[Mux.scala 27:72]
  wire  _T_22344 = bht_rd_addr_hashed_p1_f == 8'h59; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22933 = _T_22344 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23188 = _T_23187 | _T_22933; // @[Mux.scala 27:72]
  wire  _T_22347 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22934 = _T_22347 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23189 = _T_23188 | _T_22934; // @[Mux.scala 27:72]
  wire  _T_22350 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22935 = _T_22350 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23190 = _T_23189 | _T_22935; // @[Mux.scala 27:72]
  wire  _T_22353 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22936 = _T_22353 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23191 = _T_23190 | _T_22936; // @[Mux.scala 27:72]
  wire  _T_22356 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22937 = _T_22356 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23192 = _T_23191 | _T_22937; // @[Mux.scala 27:72]
  wire  _T_22359 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22938 = _T_22359 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23193 = _T_23192 | _T_22938; // @[Mux.scala 27:72]
  wire  _T_22362 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22939 = _T_22362 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23194 = _T_23193 | _T_22939; // @[Mux.scala 27:72]
  wire  _T_22365 = bht_rd_addr_hashed_p1_f == 8'h60; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22940 = _T_22365 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23195 = _T_23194 | _T_22940; // @[Mux.scala 27:72]
  wire  _T_22368 = bht_rd_addr_hashed_p1_f == 8'h61; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22941 = _T_22368 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23196 = _T_23195 | _T_22941; // @[Mux.scala 27:72]
  wire  _T_22371 = bht_rd_addr_hashed_p1_f == 8'h62; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22942 = _T_22371 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23197 = _T_23196 | _T_22942; // @[Mux.scala 27:72]
  wire  _T_22374 = bht_rd_addr_hashed_p1_f == 8'h63; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22943 = _T_22374 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23198 = _T_23197 | _T_22943; // @[Mux.scala 27:72]
  wire  _T_22377 = bht_rd_addr_hashed_p1_f == 8'h64; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22944 = _T_22377 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23199 = _T_23198 | _T_22944; // @[Mux.scala 27:72]
  wire  _T_22380 = bht_rd_addr_hashed_p1_f == 8'h65; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22945 = _T_22380 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23200 = _T_23199 | _T_22945; // @[Mux.scala 27:72]
  wire  _T_22383 = bht_rd_addr_hashed_p1_f == 8'h66; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22946 = _T_22383 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23201 = _T_23200 | _T_22946; // @[Mux.scala 27:72]
  wire  _T_22386 = bht_rd_addr_hashed_p1_f == 8'h67; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22947 = _T_22386 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23202 = _T_23201 | _T_22947; // @[Mux.scala 27:72]
  wire  _T_22389 = bht_rd_addr_hashed_p1_f == 8'h68; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22948 = _T_22389 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23203 = _T_23202 | _T_22948; // @[Mux.scala 27:72]
  wire  _T_22392 = bht_rd_addr_hashed_p1_f == 8'h69; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22949 = _T_22392 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23204 = _T_23203 | _T_22949; // @[Mux.scala 27:72]
  wire  _T_22395 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22950 = _T_22395 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23205 = _T_23204 | _T_22950; // @[Mux.scala 27:72]
  wire  _T_22398 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22951 = _T_22398 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23206 = _T_23205 | _T_22951; // @[Mux.scala 27:72]
  wire  _T_22401 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22952 = _T_22401 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23207 = _T_23206 | _T_22952; // @[Mux.scala 27:72]
  wire  _T_22404 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22953 = _T_22404 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23208 = _T_23207 | _T_22953; // @[Mux.scala 27:72]
  wire  _T_22407 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22954 = _T_22407 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23209 = _T_23208 | _T_22954; // @[Mux.scala 27:72]
  wire  _T_22410 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22955 = _T_22410 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23210 = _T_23209 | _T_22955; // @[Mux.scala 27:72]
  wire  _T_22413 = bht_rd_addr_hashed_p1_f == 8'h70; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22956 = _T_22413 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23211 = _T_23210 | _T_22956; // @[Mux.scala 27:72]
  wire  _T_22416 = bht_rd_addr_hashed_p1_f == 8'h71; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22957 = _T_22416 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23212 = _T_23211 | _T_22957; // @[Mux.scala 27:72]
  wire  _T_22419 = bht_rd_addr_hashed_p1_f == 8'h72; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22958 = _T_22419 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23213 = _T_23212 | _T_22958; // @[Mux.scala 27:72]
  wire  _T_22422 = bht_rd_addr_hashed_p1_f == 8'h73; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22959 = _T_22422 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23214 = _T_23213 | _T_22959; // @[Mux.scala 27:72]
  wire  _T_22425 = bht_rd_addr_hashed_p1_f == 8'h74; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22960 = _T_22425 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23215 = _T_23214 | _T_22960; // @[Mux.scala 27:72]
  wire  _T_22428 = bht_rd_addr_hashed_p1_f == 8'h75; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22961 = _T_22428 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23216 = _T_23215 | _T_22961; // @[Mux.scala 27:72]
  wire  _T_22431 = bht_rd_addr_hashed_p1_f == 8'h76; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22962 = _T_22431 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23217 = _T_23216 | _T_22962; // @[Mux.scala 27:72]
  wire  _T_22434 = bht_rd_addr_hashed_p1_f == 8'h77; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22963 = _T_22434 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23218 = _T_23217 | _T_22963; // @[Mux.scala 27:72]
  wire  _T_22437 = bht_rd_addr_hashed_p1_f == 8'h78; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22964 = _T_22437 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23219 = _T_23218 | _T_22964; // @[Mux.scala 27:72]
  wire  _T_22440 = bht_rd_addr_hashed_p1_f == 8'h79; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22965 = _T_22440 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23220 = _T_23219 | _T_22965; // @[Mux.scala 27:72]
  wire  _T_22443 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22966 = _T_22443 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23221 = _T_23220 | _T_22966; // @[Mux.scala 27:72]
  wire  _T_22446 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22967 = _T_22446 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23222 = _T_23221 | _T_22967; // @[Mux.scala 27:72]
  wire  _T_22449 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22968 = _T_22449 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23223 = _T_23222 | _T_22968; // @[Mux.scala 27:72]
  wire  _T_22452 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22969 = _T_22452 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23224 = _T_23223 | _T_22969; // @[Mux.scala 27:72]
  wire  _T_22455 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22970 = _T_22455 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23225 = _T_23224 | _T_22970; // @[Mux.scala 27:72]
  wire  _T_22458 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22971 = _T_22458 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23226 = _T_23225 | _T_22971; // @[Mux.scala 27:72]
  wire  _T_22461 = bht_rd_addr_hashed_p1_f == 8'h80; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22972 = _T_22461 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23227 = _T_23226 | _T_22972; // @[Mux.scala 27:72]
  wire  _T_22464 = bht_rd_addr_hashed_p1_f == 8'h81; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22973 = _T_22464 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23228 = _T_23227 | _T_22973; // @[Mux.scala 27:72]
  wire  _T_22467 = bht_rd_addr_hashed_p1_f == 8'h82; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22974 = _T_22467 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23229 = _T_23228 | _T_22974; // @[Mux.scala 27:72]
  wire  _T_22470 = bht_rd_addr_hashed_p1_f == 8'h83; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22975 = _T_22470 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23230 = _T_23229 | _T_22975; // @[Mux.scala 27:72]
  wire  _T_22473 = bht_rd_addr_hashed_p1_f == 8'h84; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22976 = _T_22473 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23231 = _T_23230 | _T_22976; // @[Mux.scala 27:72]
  wire  _T_22476 = bht_rd_addr_hashed_p1_f == 8'h85; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22977 = _T_22476 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23232 = _T_23231 | _T_22977; // @[Mux.scala 27:72]
  wire  _T_22479 = bht_rd_addr_hashed_p1_f == 8'h86; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22978 = _T_22479 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23233 = _T_23232 | _T_22978; // @[Mux.scala 27:72]
  wire  _T_22482 = bht_rd_addr_hashed_p1_f == 8'h87; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22979 = _T_22482 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23234 = _T_23233 | _T_22979; // @[Mux.scala 27:72]
  wire  _T_22485 = bht_rd_addr_hashed_p1_f == 8'h88; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22980 = _T_22485 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23235 = _T_23234 | _T_22980; // @[Mux.scala 27:72]
  wire  _T_22488 = bht_rd_addr_hashed_p1_f == 8'h89; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22981 = _T_22488 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23236 = _T_23235 | _T_22981; // @[Mux.scala 27:72]
  wire  _T_22491 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22982 = _T_22491 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23237 = _T_23236 | _T_22982; // @[Mux.scala 27:72]
  wire  _T_22494 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22983 = _T_22494 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23238 = _T_23237 | _T_22983; // @[Mux.scala 27:72]
  wire  _T_22497 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22984 = _T_22497 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23239 = _T_23238 | _T_22984; // @[Mux.scala 27:72]
  wire  _T_22500 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22985 = _T_22500 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23240 = _T_23239 | _T_22985; // @[Mux.scala 27:72]
  wire  _T_22503 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22986 = _T_22503 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23241 = _T_23240 | _T_22986; // @[Mux.scala 27:72]
  wire  _T_22506 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22987 = _T_22506 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23242 = _T_23241 | _T_22987; // @[Mux.scala 27:72]
  wire  _T_22509 = bht_rd_addr_hashed_p1_f == 8'h90; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22988 = _T_22509 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23243 = _T_23242 | _T_22988; // @[Mux.scala 27:72]
  wire  _T_22512 = bht_rd_addr_hashed_p1_f == 8'h91; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22989 = _T_22512 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23244 = _T_23243 | _T_22989; // @[Mux.scala 27:72]
  wire  _T_22515 = bht_rd_addr_hashed_p1_f == 8'h92; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22990 = _T_22515 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23245 = _T_23244 | _T_22990; // @[Mux.scala 27:72]
  wire  _T_22518 = bht_rd_addr_hashed_p1_f == 8'h93; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22991 = _T_22518 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23246 = _T_23245 | _T_22991; // @[Mux.scala 27:72]
  wire  _T_22521 = bht_rd_addr_hashed_p1_f == 8'h94; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22992 = _T_22521 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23247 = _T_23246 | _T_22992; // @[Mux.scala 27:72]
  wire  _T_22524 = bht_rd_addr_hashed_p1_f == 8'h95; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22993 = _T_22524 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23248 = _T_23247 | _T_22993; // @[Mux.scala 27:72]
  wire  _T_22527 = bht_rd_addr_hashed_p1_f == 8'h96; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22994 = _T_22527 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23249 = _T_23248 | _T_22994; // @[Mux.scala 27:72]
  wire  _T_22530 = bht_rd_addr_hashed_p1_f == 8'h97; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22995 = _T_22530 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23250 = _T_23249 | _T_22995; // @[Mux.scala 27:72]
  wire  _T_22533 = bht_rd_addr_hashed_p1_f == 8'h98; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22996 = _T_22533 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23251 = _T_23250 | _T_22996; // @[Mux.scala 27:72]
  wire  _T_22536 = bht_rd_addr_hashed_p1_f == 8'h99; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22997 = _T_22536 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23252 = _T_23251 | _T_22997; // @[Mux.scala 27:72]
  wire  _T_22539 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22998 = _T_22539 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23253 = _T_23252 | _T_22998; // @[Mux.scala 27:72]
  wire  _T_22542 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_22999 = _T_22542 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23254 = _T_23253 | _T_22999; // @[Mux.scala 27:72]
  wire  _T_22545 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23000 = _T_22545 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23255 = _T_23254 | _T_23000; // @[Mux.scala 27:72]
  wire  _T_22548 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23001 = _T_22548 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23256 = _T_23255 | _T_23001; // @[Mux.scala 27:72]
  wire  _T_22551 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23002 = _T_22551 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23257 = _T_23256 | _T_23002; // @[Mux.scala 27:72]
  wire  _T_22554 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23003 = _T_22554 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23258 = _T_23257 | _T_23003; // @[Mux.scala 27:72]
  wire  _T_22557 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23004 = _T_22557 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23259 = _T_23258 | _T_23004; // @[Mux.scala 27:72]
  wire  _T_22560 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23005 = _T_22560 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23260 = _T_23259 | _T_23005; // @[Mux.scala 27:72]
  wire  _T_22563 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23006 = _T_22563 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23261 = _T_23260 | _T_23006; // @[Mux.scala 27:72]
  wire  _T_22566 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23007 = _T_22566 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23262 = _T_23261 | _T_23007; // @[Mux.scala 27:72]
  wire  _T_22569 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23008 = _T_22569 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23263 = _T_23262 | _T_23008; // @[Mux.scala 27:72]
  wire  _T_22572 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23009 = _T_22572 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23264 = _T_23263 | _T_23009; // @[Mux.scala 27:72]
  wire  _T_22575 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23010 = _T_22575 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23265 = _T_23264 | _T_23010; // @[Mux.scala 27:72]
  wire  _T_22578 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23011 = _T_22578 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23266 = _T_23265 | _T_23011; // @[Mux.scala 27:72]
  wire  _T_22581 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23012 = _T_22581 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23267 = _T_23266 | _T_23012; // @[Mux.scala 27:72]
  wire  _T_22584 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23013 = _T_22584 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23268 = _T_23267 | _T_23013; // @[Mux.scala 27:72]
  wire  _T_22587 = bht_rd_addr_hashed_p1_f == 8'haa; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23014 = _T_22587 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23269 = _T_23268 | _T_23014; // @[Mux.scala 27:72]
  wire  _T_22590 = bht_rd_addr_hashed_p1_f == 8'hab; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23015 = _T_22590 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23270 = _T_23269 | _T_23015; // @[Mux.scala 27:72]
  wire  _T_22593 = bht_rd_addr_hashed_p1_f == 8'hac; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23016 = _T_22593 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23271 = _T_23270 | _T_23016; // @[Mux.scala 27:72]
  wire  _T_22596 = bht_rd_addr_hashed_p1_f == 8'had; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23017 = _T_22596 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23272 = _T_23271 | _T_23017; // @[Mux.scala 27:72]
  wire  _T_22599 = bht_rd_addr_hashed_p1_f == 8'hae; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23018 = _T_22599 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23273 = _T_23272 | _T_23018; // @[Mux.scala 27:72]
  wire  _T_22602 = bht_rd_addr_hashed_p1_f == 8'haf; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23019 = _T_22602 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23274 = _T_23273 | _T_23019; // @[Mux.scala 27:72]
  wire  _T_22605 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23020 = _T_22605 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23275 = _T_23274 | _T_23020; // @[Mux.scala 27:72]
  wire  _T_22608 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23021 = _T_22608 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23276 = _T_23275 | _T_23021; // @[Mux.scala 27:72]
  wire  _T_22611 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23022 = _T_22611 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23277 = _T_23276 | _T_23022; // @[Mux.scala 27:72]
  wire  _T_22614 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23023 = _T_22614 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23278 = _T_23277 | _T_23023; // @[Mux.scala 27:72]
  wire  _T_22617 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23024 = _T_22617 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23279 = _T_23278 | _T_23024; // @[Mux.scala 27:72]
  wire  _T_22620 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23025 = _T_22620 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23280 = _T_23279 | _T_23025; // @[Mux.scala 27:72]
  wire  _T_22623 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23026 = _T_22623 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23281 = _T_23280 | _T_23026; // @[Mux.scala 27:72]
  wire  _T_22626 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23027 = _T_22626 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23282 = _T_23281 | _T_23027; // @[Mux.scala 27:72]
  wire  _T_22629 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23028 = _T_22629 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23283 = _T_23282 | _T_23028; // @[Mux.scala 27:72]
  wire  _T_22632 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23029 = _T_22632 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23284 = _T_23283 | _T_23029; // @[Mux.scala 27:72]
  wire  _T_22635 = bht_rd_addr_hashed_p1_f == 8'hba; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23030 = _T_22635 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23285 = _T_23284 | _T_23030; // @[Mux.scala 27:72]
  wire  _T_22638 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23031 = _T_22638 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23286 = _T_23285 | _T_23031; // @[Mux.scala 27:72]
  wire  _T_22641 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23032 = _T_22641 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23287 = _T_23286 | _T_23032; // @[Mux.scala 27:72]
  wire  _T_22644 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23033 = _T_22644 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23288 = _T_23287 | _T_23033; // @[Mux.scala 27:72]
  wire  _T_22647 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23034 = _T_22647 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23289 = _T_23288 | _T_23034; // @[Mux.scala 27:72]
  wire  _T_22650 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23035 = _T_22650 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23290 = _T_23289 | _T_23035; // @[Mux.scala 27:72]
  wire  _T_22653 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23036 = _T_22653 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23291 = _T_23290 | _T_23036; // @[Mux.scala 27:72]
  wire  _T_22656 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23037 = _T_22656 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23292 = _T_23291 | _T_23037; // @[Mux.scala 27:72]
  wire  _T_22659 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23038 = _T_22659 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23293 = _T_23292 | _T_23038; // @[Mux.scala 27:72]
  wire  _T_22662 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23039 = _T_22662 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23294 = _T_23293 | _T_23039; // @[Mux.scala 27:72]
  wire  _T_22665 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23040 = _T_22665 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23295 = _T_23294 | _T_23040; // @[Mux.scala 27:72]
  wire  _T_22668 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23041 = _T_22668 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23296 = _T_23295 | _T_23041; // @[Mux.scala 27:72]
  wire  _T_22671 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23042 = _T_22671 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23297 = _T_23296 | _T_23042; // @[Mux.scala 27:72]
  wire  _T_22674 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23043 = _T_22674 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23298 = _T_23297 | _T_23043; // @[Mux.scala 27:72]
  wire  _T_22677 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23044 = _T_22677 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23299 = _T_23298 | _T_23044; // @[Mux.scala 27:72]
  wire  _T_22680 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23045 = _T_22680 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23300 = _T_23299 | _T_23045; // @[Mux.scala 27:72]
  wire  _T_22683 = bht_rd_addr_hashed_p1_f == 8'hca; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23046 = _T_22683 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23301 = _T_23300 | _T_23046; // @[Mux.scala 27:72]
  wire  _T_22686 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23047 = _T_22686 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23302 = _T_23301 | _T_23047; // @[Mux.scala 27:72]
  wire  _T_22689 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23048 = _T_22689 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23303 = _T_23302 | _T_23048; // @[Mux.scala 27:72]
  wire  _T_22692 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23049 = _T_22692 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23304 = _T_23303 | _T_23049; // @[Mux.scala 27:72]
  wire  _T_22695 = bht_rd_addr_hashed_p1_f == 8'hce; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23050 = _T_22695 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23305 = _T_23304 | _T_23050; // @[Mux.scala 27:72]
  wire  _T_22698 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23051 = _T_22698 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23306 = _T_23305 | _T_23051; // @[Mux.scala 27:72]
  wire  _T_22701 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23052 = _T_22701 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23307 = _T_23306 | _T_23052; // @[Mux.scala 27:72]
  wire  _T_22704 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23053 = _T_22704 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23308 = _T_23307 | _T_23053; // @[Mux.scala 27:72]
  wire  _T_22707 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23054 = _T_22707 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23309 = _T_23308 | _T_23054; // @[Mux.scala 27:72]
  wire  _T_22710 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23055 = _T_22710 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23310 = _T_23309 | _T_23055; // @[Mux.scala 27:72]
  wire  _T_22713 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23056 = _T_22713 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23311 = _T_23310 | _T_23056; // @[Mux.scala 27:72]
  wire  _T_22716 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23057 = _T_22716 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23312 = _T_23311 | _T_23057; // @[Mux.scala 27:72]
  wire  _T_22719 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23058 = _T_22719 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23313 = _T_23312 | _T_23058; // @[Mux.scala 27:72]
  wire  _T_22722 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23059 = _T_22722 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23314 = _T_23313 | _T_23059; // @[Mux.scala 27:72]
  wire  _T_22725 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23060 = _T_22725 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23315 = _T_23314 | _T_23060; // @[Mux.scala 27:72]
  wire  _T_22728 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23061 = _T_22728 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23316 = _T_23315 | _T_23061; // @[Mux.scala 27:72]
  wire  _T_22731 = bht_rd_addr_hashed_p1_f == 8'hda; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23062 = _T_22731 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23317 = _T_23316 | _T_23062; // @[Mux.scala 27:72]
  wire  _T_22734 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23063 = _T_22734 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23318 = _T_23317 | _T_23063; // @[Mux.scala 27:72]
  wire  _T_22737 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23064 = _T_22737 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23319 = _T_23318 | _T_23064; // @[Mux.scala 27:72]
  wire  _T_22740 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23065 = _T_22740 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23320 = _T_23319 | _T_23065; // @[Mux.scala 27:72]
  wire  _T_22743 = bht_rd_addr_hashed_p1_f == 8'hde; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23066 = _T_22743 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23321 = _T_23320 | _T_23066; // @[Mux.scala 27:72]
  wire  _T_22746 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23067 = _T_22746 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23322 = _T_23321 | _T_23067; // @[Mux.scala 27:72]
  wire  _T_22749 = bht_rd_addr_hashed_p1_f == 8'he0; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23068 = _T_22749 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23323 = _T_23322 | _T_23068; // @[Mux.scala 27:72]
  wire  _T_22752 = bht_rd_addr_hashed_p1_f == 8'he1; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23069 = _T_22752 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23324 = _T_23323 | _T_23069; // @[Mux.scala 27:72]
  wire  _T_22755 = bht_rd_addr_hashed_p1_f == 8'he2; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23070 = _T_22755 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23325 = _T_23324 | _T_23070; // @[Mux.scala 27:72]
  wire  _T_22758 = bht_rd_addr_hashed_p1_f == 8'he3; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23071 = _T_22758 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23326 = _T_23325 | _T_23071; // @[Mux.scala 27:72]
  wire  _T_22761 = bht_rd_addr_hashed_p1_f == 8'he4; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23072 = _T_22761 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23327 = _T_23326 | _T_23072; // @[Mux.scala 27:72]
  wire  _T_22764 = bht_rd_addr_hashed_p1_f == 8'he5; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23073 = _T_22764 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23328 = _T_23327 | _T_23073; // @[Mux.scala 27:72]
  wire  _T_22767 = bht_rd_addr_hashed_p1_f == 8'he6; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23074 = _T_22767 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23329 = _T_23328 | _T_23074; // @[Mux.scala 27:72]
  wire  _T_22770 = bht_rd_addr_hashed_p1_f == 8'he7; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23075 = _T_22770 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23330 = _T_23329 | _T_23075; // @[Mux.scala 27:72]
  wire  _T_22773 = bht_rd_addr_hashed_p1_f == 8'he8; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23076 = _T_22773 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23331 = _T_23330 | _T_23076; // @[Mux.scala 27:72]
  wire  _T_22776 = bht_rd_addr_hashed_p1_f == 8'he9; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23077 = _T_22776 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23332 = _T_23331 | _T_23077; // @[Mux.scala 27:72]
  wire  _T_22779 = bht_rd_addr_hashed_p1_f == 8'hea; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23078 = _T_22779 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23333 = _T_23332 | _T_23078; // @[Mux.scala 27:72]
  wire  _T_22782 = bht_rd_addr_hashed_p1_f == 8'heb; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23079 = _T_22782 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23334 = _T_23333 | _T_23079; // @[Mux.scala 27:72]
  wire  _T_22785 = bht_rd_addr_hashed_p1_f == 8'hec; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23080 = _T_22785 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23335 = _T_23334 | _T_23080; // @[Mux.scala 27:72]
  wire  _T_22788 = bht_rd_addr_hashed_p1_f == 8'hed; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23081 = _T_22788 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23336 = _T_23335 | _T_23081; // @[Mux.scala 27:72]
  wire  _T_22791 = bht_rd_addr_hashed_p1_f == 8'hee; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23082 = _T_22791 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23337 = _T_23336 | _T_23082; // @[Mux.scala 27:72]
  wire  _T_22794 = bht_rd_addr_hashed_p1_f == 8'hef; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23083 = _T_22794 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23338 = _T_23337 | _T_23083; // @[Mux.scala 27:72]
  wire  _T_22797 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23084 = _T_22797 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23339 = _T_23338 | _T_23084; // @[Mux.scala 27:72]
  wire  _T_22800 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23085 = _T_22800 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23340 = _T_23339 | _T_23085; // @[Mux.scala 27:72]
  wire  _T_22803 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23086 = _T_22803 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23341 = _T_23340 | _T_23086; // @[Mux.scala 27:72]
  wire  _T_22806 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23087 = _T_22806 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23342 = _T_23341 | _T_23087; // @[Mux.scala 27:72]
  wire  _T_22809 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23088 = _T_22809 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23343 = _T_23342 | _T_23088; // @[Mux.scala 27:72]
  wire  _T_22812 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23089 = _T_22812 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23344 = _T_23343 | _T_23089; // @[Mux.scala 27:72]
  wire  _T_22815 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23090 = _T_22815 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23345 = _T_23344 | _T_23090; // @[Mux.scala 27:72]
  wire  _T_22818 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23091 = _T_22818 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23346 = _T_23345 | _T_23091; // @[Mux.scala 27:72]
  wire  _T_22821 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23092 = _T_22821 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23347 = _T_23346 | _T_23092; // @[Mux.scala 27:72]
  wire  _T_22824 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23093 = _T_22824 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23348 = _T_23347 | _T_23093; // @[Mux.scala 27:72]
  wire  _T_22827 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23094 = _T_22827 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23349 = _T_23348 | _T_23094; // @[Mux.scala 27:72]
  wire  _T_22830 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23095 = _T_22830 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23350 = _T_23349 | _T_23095; // @[Mux.scala 27:72]
  wire  _T_22833 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23096 = _T_22833 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23351 = _T_23350 | _T_23096; // @[Mux.scala 27:72]
  wire  _T_22836 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23097 = _T_22836 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23352 = _T_23351 | _T_23097; // @[Mux.scala 27:72]
  wire  _T_22839 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23098 = _T_22839 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23353 = _T_23352 | _T_23098; // @[Mux.scala 27:72]
  wire  _T_22842 = bht_rd_addr_hashed_p1_f == 8'hff; // @[el2_ifu_bp_ctl.scala 389:112]
  wire [1:0] _T_23099 = _T_22842 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_23353 | _T_23099; // @[Mux.scala 27:72]
  wire [1:0] _T_259 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_258 | _T_259; // @[Mux.scala 27:72]
  wire  _T_263 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 251:42]
  wire [1:0] wayhit_f = tag_match_way0_expanded_f | tag_match_way1_expanded_f; // @[el2_ifu_bp_ctl.scala 162:44]
  wire [1:0] _T_158 = _T_143 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = tag_match_way0_expanded_p1_f | tag_match_way1_expanded_p1_f; // @[el2_ifu_bp_ctl.scala 164:50]
  wire [1:0] _T_157 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_159 = io_ifc_fetch_addr_f[0] ? _T_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_160 = _T_158 | _T_159; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[el2_ifu_bp_ctl.scala 220:64]
  wire  _T_217 = ~eoc_near; // @[el2_ifu_bp_ctl.scala 222:15]
  wire  _T_219 = |io_ifc_fetch_addr_f[1:0]; // @[el2_ifu_bp_ctl.scala 222:57]
  wire  _T_220 = ~_T_219; // @[el2_ifu_bp_ctl.scala 222:28]
  wire  eoc_mask = _T_217 | _T_220; // @[el2_ifu_bp_ctl.scala 222:25]
  wire [1:0] _T_162 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] bht_valid_f = _T_160 & _T_162; // @[el2_ifu_bp_ctl.scala 191:71]
  wire  _T_265 = _T_263 & bht_valid_f[1]; // @[el2_ifu_bp_ctl.scala 251:69]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_20284 = _T_20797 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_20285 = _T_20800 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20540 = _T_20284 | _T_20285; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_20286 = _T_20803 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20541 = _T_20540 | _T_20286; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_20287 = _T_20806 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20542 = _T_20541 | _T_20287; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_20288 = _T_20809 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20543 = _T_20542 | _T_20288; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_20289 = _T_20812 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20544 = _T_20543 | _T_20289; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_20290 = _T_20815 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20545 = _T_20544 | _T_20290; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_20291 = _T_20818 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20546 = _T_20545 | _T_20291; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_20292 = _T_20821 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20547 = _T_20546 | _T_20292; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_20293 = _T_20824 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20548 = _T_20547 | _T_20293; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_20294 = _T_20827 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20549 = _T_20548 | _T_20294; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_20295 = _T_20830 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20550 = _T_20549 | _T_20295; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_20296 = _T_20833 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20551 = _T_20550 | _T_20296; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_20297 = _T_20836 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20552 = _T_20551 | _T_20297; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_20298 = _T_20839 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20553 = _T_20552 | _T_20298; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_20299 = _T_20842 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20554 = _T_20553 | _T_20299; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_20300 = _T_20845 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20555 = _T_20554 | _T_20300; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_20301 = _T_20848 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20556 = _T_20555 | _T_20301; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_20302 = _T_20851 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20557 = _T_20556 | _T_20302; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_20303 = _T_20854 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20558 = _T_20557 | _T_20303; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_20304 = _T_20857 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20559 = _T_20558 | _T_20304; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_20305 = _T_20860 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20560 = _T_20559 | _T_20305; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_20306 = _T_20863 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20561 = _T_20560 | _T_20306; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_20307 = _T_20866 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20562 = _T_20561 | _T_20307; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_20308 = _T_20869 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20563 = _T_20562 | _T_20308; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_20309 = _T_20872 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20564 = _T_20563 | _T_20309; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_20310 = _T_20875 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20565 = _T_20564 | _T_20310; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_20311 = _T_20878 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20566 = _T_20565 | _T_20311; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_20312 = _T_20881 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20567 = _T_20566 | _T_20312; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_20313 = _T_20884 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20568 = _T_20567 | _T_20313; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_20314 = _T_20887 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20569 = _T_20568 | _T_20314; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_20315 = _T_20890 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20570 = _T_20569 | _T_20315; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_20316 = _T_20893 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20571 = _T_20570 | _T_20316; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_20317 = _T_20896 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20572 = _T_20571 | _T_20317; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_20318 = _T_20899 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20573 = _T_20572 | _T_20318; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_20319 = _T_20902 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20574 = _T_20573 | _T_20319; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_20320 = _T_20905 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20575 = _T_20574 | _T_20320; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_20321 = _T_20908 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20576 = _T_20575 | _T_20321; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_20322 = _T_20911 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20577 = _T_20576 | _T_20322; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_20323 = _T_20914 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20578 = _T_20577 | _T_20323; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_20324 = _T_20917 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20579 = _T_20578 | _T_20324; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_20325 = _T_20920 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20580 = _T_20579 | _T_20325; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_20326 = _T_20923 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20581 = _T_20580 | _T_20326; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_20327 = _T_20926 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20582 = _T_20581 | _T_20327; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_20328 = _T_20929 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20583 = _T_20582 | _T_20328; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_20329 = _T_20932 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20584 = _T_20583 | _T_20329; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_20330 = _T_20935 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20585 = _T_20584 | _T_20330; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_20331 = _T_20938 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20586 = _T_20585 | _T_20331; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_20332 = _T_20941 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20587 = _T_20586 | _T_20332; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_20333 = _T_20944 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20588 = _T_20587 | _T_20333; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_20334 = _T_20947 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20589 = _T_20588 | _T_20334; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_20335 = _T_20950 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20590 = _T_20589 | _T_20335; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_20336 = _T_20953 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20591 = _T_20590 | _T_20336; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_20337 = _T_20956 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20592 = _T_20591 | _T_20337; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_20338 = _T_20959 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20593 = _T_20592 | _T_20338; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_20339 = _T_20962 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20594 = _T_20593 | _T_20339; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_20340 = _T_20965 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20595 = _T_20594 | _T_20340; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_20341 = _T_20968 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20596 = _T_20595 | _T_20341; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_20342 = _T_20971 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20597 = _T_20596 | _T_20342; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_20343 = _T_20974 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20598 = _T_20597 | _T_20343; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_20344 = _T_20977 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20599 = _T_20598 | _T_20344; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_20345 = _T_20980 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20600 = _T_20599 | _T_20345; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_20346 = _T_20983 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20601 = _T_20600 | _T_20346; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_20347 = _T_20986 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20602 = _T_20601 | _T_20347; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_20348 = _T_20989 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20603 = _T_20602 | _T_20348; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_20349 = _T_20992 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20604 = _T_20603 | _T_20349; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_20350 = _T_20995 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20605 = _T_20604 | _T_20350; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_20351 = _T_20998 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20606 = _T_20605 | _T_20351; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_20352 = _T_21001 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20607 = _T_20606 | _T_20352; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_20353 = _T_21004 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20608 = _T_20607 | _T_20353; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_20354 = _T_21007 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20609 = _T_20608 | _T_20354; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_20355 = _T_21010 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20610 = _T_20609 | _T_20355; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_20356 = _T_21013 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20611 = _T_20610 | _T_20356; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_20357 = _T_21016 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20612 = _T_20611 | _T_20357; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_20358 = _T_21019 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20613 = _T_20612 | _T_20358; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_20359 = _T_21022 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20614 = _T_20613 | _T_20359; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_20360 = _T_21025 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20615 = _T_20614 | _T_20360; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_20361 = _T_21028 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20616 = _T_20615 | _T_20361; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_20362 = _T_21031 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20617 = _T_20616 | _T_20362; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_20363 = _T_21034 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20618 = _T_20617 | _T_20363; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_20364 = _T_21037 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20619 = _T_20618 | _T_20364; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_20365 = _T_21040 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20620 = _T_20619 | _T_20365; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_20366 = _T_21043 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20621 = _T_20620 | _T_20366; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_20367 = _T_21046 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20622 = _T_20621 | _T_20367; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_20368 = _T_21049 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20623 = _T_20622 | _T_20368; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_20369 = _T_21052 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20624 = _T_20623 | _T_20369; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_20370 = _T_21055 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20625 = _T_20624 | _T_20370; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_20371 = _T_21058 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20626 = _T_20625 | _T_20371; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_20372 = _T_21061 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20627 = _T_20626 | _T_20372; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_20373 = _T_21064 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20628 = _T_20627 | _T_20373; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_20374 = _T_21067 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20629 = _T_20628 | _T_20374; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_20375 = _T_21070 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20630 = _T_20629 | _T_20375; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_20376 = _T_21073 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20631 = _T_20630 | _T_20376; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_20377 = _T_21076 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20632 = _T_20631 | _T_20377; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_20378 = _T_21079 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20633 = _T_20632 | _T_20378; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_20379 = _T_21082 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20634 = _T_20633 | _T_20379; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_20380 = _T_21085 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20635 = _T_20634 | _T_20380; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_20381 = _T_21088 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20636 = _T_20635 | _T_20381; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_20382 = _T_21091 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20637 = _T_20636 | _T_20382; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_20383 = _T_21094 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20638 = _T_20637 | _T_20383; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_20384 = _T_21097 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20639 = _T_20638 | _T_20384; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_20385 = _T_21100 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20640 = _T_20639 | _T_20385; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_20386 = _T_21103 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20641 = _T_20640 | _T_20386; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_20387 = _T_21106 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20642 = _T_20641 | _T_20387; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_20388 = _T_21109 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20643 = _T_20642 | _T_20388; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_20389 = _T_21112 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20644 = _T_20643 | _T_20389; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_20390 = _T_21115 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20645 = _T_20644 | _T_20390; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_20391 = _T_21118 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20646 = _T_20645 | _T_20391; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_20392 = _T_21121 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20647 = _T_20646 | _T_20392; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_20393 = _T_21124 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20648 = _T_20647 | _T_20393; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_20394 = _T_21127 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20649 = _T_20648 | _T_20394; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_20395 = _T_21130 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20650 = _T_20649 | _T_20395; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_20396 = _T_21133 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20651 = _T_20650 | _T_20396; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_20397 = _T_21136 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20652 = _T_20651 | _T_20397; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_20398 = _T_21139 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20653 = _T_20652 | _T_20398; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_20399 = _T_21142 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20654 = _T_20653 | _T_20399; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_20400 = _T_21145 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20655 = _T_20654 | _T_20400; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_20401 = _T_21148 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20656 = _T_20655 | _T_20401; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_20402 = _T_21151 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20657 = _T_20656 | _T_20402; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_20403 = _T_21154 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20658 = _T_20657 | _T_20403; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_20404 = _T_21157 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20659 = _T_20658 | _T_20404; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_20405 = _T_21160 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20660 = _T_20659 | _T_20405; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_20406 = _T_21163 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20661 = _T_20660 | _T_20406; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_20407 = _T_21166 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20662 = _T_20661 | _T_20407; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_20408 = _T_21169 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20663 = _T_20662 | _T_20408; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_20409 = _T_21172 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20664 = _T_20663 | _T_20409; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_20410 = _T_21175 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20665 = _T_20664 | _T_20410; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_20411 = _T_21178 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20666 = _T_20665 | _T_20411; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_20412 = _T_21181 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20667 = _T_20666 | _T_20412; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_20413 = _T_21184 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20668 = _T_20667 | _T_20413; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_20414 = _T_21187 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20669 = _T_20668 | _T_20414; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_20415 = _T_21190 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20670 = _T_20669 | _T_20415; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_20416 = _T_21193 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20671 = _T_20670 | _T_20416; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_20417 = _T_21196 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20672 = _T_20671 | _T_20417; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_20418 = _T_21199 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20673 = _T_20672 | _T_20418; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_20419 = _T_21202 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20674 = _T_20673 | _T_20419; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_20420 = _T_21205 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20675 = _T_20674 | _T_20420; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_20421 = _T_21208 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20676 = _T_20675 | _T_20421; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_20422 = _T_21211 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20677 = _T_20676 | _T_20422; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_20423 = _T_21214 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20678 = _T_20677 | _T_20423; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_20424 = _T_21217 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20679 = _T_20678 | _T_20424; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_20425 = _T_21220 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20680 = _T_20679 | _T_20425; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_20426 = _T_21223 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20681 = _T_20680 | _T_20426; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_20427 = _T_21226 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20682 = _T_20681 | _T_20427; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_20428 = _T_21229 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20683 = _T_20682 | _T_20428; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_20429 = _T_21232 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20684 = _T_20683 | _T_20429; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_20430 = _T_21235 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20685 = _T_20684 | _T_20430; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_20431 = _T_21238 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20686 = _T_20685 | _T_20431; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_20432 = _T_21241 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20687 = _T_20686 | _T_20432; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_20433 = _T_21244 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20688 = _T_20687 | _T_20433; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_20434 = _T_21247 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20689 = _T_20688 | _T_20434; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_20435 = _T_21250 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20690 = _T_20689 | _T_20435; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_20436 = _T_21253 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20691 = _T_20690 | _T_20436; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_20437 = _T_21256 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20692 = _T_20691 | _T_20437; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_20438 = _T_21259 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20693 = _T_20692 | _T_20438; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_20439 = _T_21262 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20694 = _T_20693 | _T_20439; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_20440 = _T_21265 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20695 = _T_20694 | _T_20440; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_20441 = _T_21268 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20696 = _T_20695 | _T_20441; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_20442 = _T_21271 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20697 = _T_20696 | _T_20442; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_20443 = _T_21274 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20698 = _T_20697 | _T_20443; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_20444 = _T_21277 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20699 = _T_20698 | _T_20444; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_20445 = _T_21280 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20700 = _T_20699 | _T_20445; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_20446 = _T_21283 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20701 = _T_20700 | _T_20446; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_20447 = _T_21286 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20702 = _T_20701 | _T_20447; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_20448 = _T_21289 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20703 = _T_20702 | _T_20448; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_20449 = _T_21292 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20704 = _T_20703 | _T_20449; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_20450 = _T_21295 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20705 = _T_20704 | _T_20450; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_20451 = _T_21298 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20706 = _T_20705 | _T_20451; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_20452 = _T_21301 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20707 = _T_20706 | _T_20452; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_20453 = _T_21304 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20708 = _T_20707 | _T_20453; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_20454 = _T_21307 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20709 = _T_20708 | _T_20454; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_20455 = _T_21310 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20710 = _T_20709 | _T_20455; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_20456 = _T_21313 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20711 = _T_20710 | _T_20456; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_20457 = _T_21316 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20712 = _T_20711 | _T_20457; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_20458 = _T_21319 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20713 = _T_20712 | _T_20458; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_20459 = _T_21322 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20714 = _T_20713 | _T_20459; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_20460 = _T_21325 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20715 = _T_20714 | _T_20460; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_20461 = _T_21328 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20716 = _T_20715 | _T_20461; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_20462 = _T_21331 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20717 = _T_20716 | _T_20462; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_20463 = _T_21334 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20718 = _T_20717 | _T_20463; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_20464 = _T_21337 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20719 = _T_20718 | _T_20464; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_20465 = _T_21340 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20720 = _T_20719 | _T_20465; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_20466 = _T_21343 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20721 = _T_20720 | _T_20466; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_20467 = _T_21346 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20722 = _T_20721 | _T_20467; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_20468 = _T_21349 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20723 = _T_20722 | _T_20468; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_20469 = _T_21352 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20724 = _T_20723 | _T_20469; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_20470 = _T_21355 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20725 = _T_20724 | _T_20470; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_20471 = _T_21358 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20726 = _T_20725 | _T_20471; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_20472 = _T_21361 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20727 = _T_20726 | _T_20472; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_20473 = _T_21364 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20728 = _T_20727 | _T_20473; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_20474 = _T_21367 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20729 = _T_20728 | _T_20474; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_20475 = _T_21370 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20730 = _T_20729 | _T_20475; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_20476 = _T_21373 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20731 = _T_20730 | _T_20476; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_20477 = _T_21376 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20732 = _T_20731 | _T_20477; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_20478 = _T_21379 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20733 = _T_20732 | _T_20478; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_20479 = _T_21382 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20734 = _T_20733 | _T_20479; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_20480 = _T_21385 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20735 = _T_20734 | _T_20480; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_20481 = _T_21388 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20736 = _T_20735 | _T_20481; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_20482 = _T_21391 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20737 = _T_20736 | _T_20482; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_20483 = _T_21394 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20738 = _T_20737 | _T_20483; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_20484 = _T_21397 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20739 = _T_20738 | _T_20484; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_20485 = _T_21400 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20740 = _T_20739 | _T_20485; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_20486 = _T_21403 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20741 = _T_20740 | _T_20486; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_20487 = _T_21406 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20742 = _T_20741 | _T_20487; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_20488 = _T_21409 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20743 = _T_20742 | _T_20488; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_20489 = _T_21412 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20744 = _T_20743 | _T_20489; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_20490 = _T_21415 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20745 = _T_20744 | _T_20490; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_20491 = _T_21418 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20746 = _T_20745 | _T_20491; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_20492 = _T_21421 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20747 = _T_20746 | _T_20492; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_20493 = _T_21424 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20748 = _T_20747 | _T_20493; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_20494 = _T_21427 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20749 = _T_20748 | _T_20494; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_20495 = _T_21430 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20750 = _T_20749 | _T_20495; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_20496 = _T_21433 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20751 = _T_20750 | _T_20496; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_20497 = _T_21436 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20752 = _T_20751 | _T_20497; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_20498 = _T_21439 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20753 = _T_20752 | _T_20498; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_20499 = _T_21442 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20754 = _T_20753 | _T_20499; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_20500 = _T_21445 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20755 = _T_20754 | _T_20500; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_20501 = _T_21448 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20756 = _T_20755 | _T_20501; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_20502 = _T_21451 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20757 = _T_20756 | _T_20502; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_20503 = _T_21454 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20758 = _T_20757 | _T_20503; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_20504 = _T_21457 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20759 = _T_20758 | _T_20504; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_20505 = _T_21460 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20760 = _T_20759 | _T_20505; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_20506 = _T_21463 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20761 = _T_20760 | _T_20506; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_20507 = _T_21466 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20762 = _T_20761 | _T_20507; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_20508 = _T_21469 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20763 = _T_20762 | _T_20508; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_20509 = _T_21472 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20764 = _T_20763 | _T_20509; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_20510 = _T_21475 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20765 = _T_20764 | _T_20510; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_20511 = _T_21478 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20766 = _T_20765 | _T_20511; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_20512 = _T_21481 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20767 = _T_20766 | _T_20512; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_20513 = _T_21484 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20768 = _T_20767 | _T_20513; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_20514 = _T_21487 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20769 = _T_20768 | _T_20514; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_20515 = _T_21490 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20770 = _T_20769 | _T_20515; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_20516 = _T_21493 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20771 = _T_20770 | _T_20516; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_20517 = _T_21496 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20772 = _T_20771 | _T_20517; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_20518 = _T_21499 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20773 = _T_20772 | _T_20518; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_20519 = _T_21502 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20774 = _T_20773 | _T_20519; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_20520 = _T_21505 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20775 = _T_20774 | _T_20520; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_20521 = _T_21508 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20776 = _T_20775 | _T_20521; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_20522 = _T_21511 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20777 = _T_20776 | _T_20522; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_20523 = _T_21514 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20778 = _T_20777 | _T_20523; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_20524 = _T_21517 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20779 = _T_20778 | _T_20524; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_20525 = _T_21520 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20780 = _T_20779 | _T_20525; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_20526 = _T_21523 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20781 = _T_20780 | _T_20526; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_20527 = _T_21526 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20782 = _T_20781 | _T_20527; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_20528 = _T_21529 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20783 = _T_20782 | _T_20528; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_20529 = _T_21532 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20784 = _T_20783 | _T_20529; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_20530 = _T_21535 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20785 = _T_20784 | _T_20530; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_20531 = _T_21538 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20786 = _T_20785 | _T_20531; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_20532 = _T_21541 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20787 = _T_20786 | _T_20532; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_20533 = _T_21544 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20788 = _T_20787 | _T_20533; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_20534 = _T_21547 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20789 = _T_20788 | _T_20534; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_20535 = _T_21550 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20790 = _T_20789 | _T_20535; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_20536 = _T_21553 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20791 = _T_20790 | _T_20536; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_20537 = _T_21556 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20792 = _T_20791 | _T_20537; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_20538 = _T_21559 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_20793 = _T_20792 | _T_20538; // @[Mux.scala 27:72]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_20539 = _T_21562 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_20793 | _T_20539; // @[Mux.scala 27:72]
  wire [1:0] _T_250 = _T_143 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_251 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_250 | _T_251; // @[Mux.scala 27:72]
  wire  _T_268 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 252:45]
  wire  _T_270 = _T_268 & bht_valid_f[0]; // @[el2_ifu_bp_ctl.scala 252:72]
  wire [1:0] bht_dir_f = {_T_265,_T_270}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[el2_ifu_bp_ctl.scala 108:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_143}; // @[Cat.scala 29:58]
  wire  _T_32 = io_exu_mp_btag == fetch_rd_tag_f; // @[el2_ifu_bp_ctl.scala 124:46]
  wire  _T_33 = _T_32 & exu_mp_valid; // @[el2_ifu_bp_ctl.scala 124:66]
  wire  _T_34 = _T_33 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 124:81]
  wire  _T_35 = io_exu_mp_index == btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 124:117]
  wire  fetch_mp_collision_f = _T_34 & _T_35; // @[el2_ifu_bp_ctl.scala 124:102]
  wire  _T_36 = io_exu_mp_btag == fetch_rd_tag_p1_f; // @[el2_ifu_bp_ctl.scala 125:49]
  wire  _T_37 = _T_36 & exu_mp_valid; // @[el2_ifu_bp_ctl.scala 125:72]
  wire  _T_38 = _T_37 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 125:87]
  wire  _T_39 = io_exu_mp_index == btb_rd_addr_p1_f; // @[el2_ifu_bp_ctl.scala 125:123]
  wire  fetch_mp_collision_p1_f = _T_38 & _T_39; // @[el2_ifu_bp_ctl.scala 125:108]
  reg  exu_mp_way_f; // @[el2_ifu_bp_ctl.scala 129:29]
  reg  exu_flush_final_d1; // @[el2_ifu_bp_ctl.scala 130:35]
  wire [255:0] mp_wrindex_dec = 256'h0 << io_exu_mp_index; // @[el2_ifu_bp_ctl.scala 183:38]
  wire [255:0] fetch_wrindex_dec = 256'h0 << btb_rd_addr_f; // @[el2_ifu_bp_ctl.scala 185:41]
  wire [255:0] fetch_wrindex_p1_dec = 256'h0 << btb_rd_addr_p1_f; // @[el2_ifu_bp_ctl.scala 187:44]
  wire [255:0] _T_149 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] mp_wrlru_b0 = mp_wrindex_dec & _T_149; // @[el2_ifu_bp_ctl.scala 189:36]
  wire  _T_165 = bht_valid_f[0] | bht_valid_f[1]; // @[el2_ifu_bp_ctl.scala 193:42]
  wire  _T_166 = _T_165 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 193:58]
  wire  lru_update_valid_f = _T_166 & _T; // @[el2_ifu_bp_ctl.scala 193:79]
  wire [255:0] _T_169 = lru_update_valid_f ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] fetch_wrlru_b0 = fetch_wrindex_dec & _T_169; // @[el2_ifu_bp_ctl.scala 195:42]
  wire [255:0] fetch_wrlru_p1_b0 = fetch_wrindex_p1_dec & _T_169; // @[el2_ifu_bp_ctl.scala 196:48]
  wire  _T_172 = mp_wrlru_b0 == 256'h0; // @[el2_ifu_bp_ctl.scala 198:25]
  wire  _T_173 = fetch_wrlru_b0 == 256'h0; // @[el2_ifu_bp_ctl.scala 198:40]
  wire  btb_lru_b0_hold = _T_172 & _T_173; // @[el2_ifu_bp_ctl.scala 198:38]
  wire  _T_175 = ~io_exu_mp_pkt_way; // @[el2_ifu_bp_ctl.scala 202:33]
  wire [255:0] _T_178 = _T_175 ? mp_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_179 = tag_match_way0_f ? fetch_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_180 = tag_match_way0_p1_f ? fetch_wrlru_p1_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_181 = _T_178 | _T_179; // @[Mux.scala 27:72]
  wire [255:0] _T_182 = _T_181 | _T_180; // @[Mux.scala 27:72]
  reg [255:0] btb_lru_b0_f; // @[Reg.scala 27:20]
  wire [255:0] _GEN_1036 = {{255'd0}, btb_lru_b0_hold}; // @[el2_ifu_bp_ctl.scala 204:100]
  wire [255:0] _T_184 = _GEN_1036 & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 204:100]
  wire [255:0] btb_lru_b0_ns = _T_182 | _T_184; // @[el2_ifu_bp_ctl.scala 204:82]
  wire [255:0] _T_186 = fetch_wrindex_dec & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 206:78]
  wire  _T_187 = |_T_186; // @[el2_ifu_bp_ctl.scala 206:94]
  wire  btb_lru_rd_f = fetch_mp_collision_f ? exu_mp_way_f : _T_187; // @[el2_ifu_bp_ctl.scala 206:25]
  wire [255:0] _T_189 = fetch_wrindex_p1_dec & btb_lru_b0_f; // @[el2_ifu_bp_ctl.scala 208:87]
  wire  _T_190 = |_T_189; // @[el2_ifu_bp_ctl.scala 208:103]
  wire  btb_lru_rd_p1_f = fetch_mp_collision_p1_f ? exu_mp_way_f : _T_190; // @[el2_ifu_bp_ctl.scala 208:28]
  wire [1:0] _T_193 = {btb_lru_rd_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_196 = {btb_lru_rd_p1_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_197 = _T_143 ? _T_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_198 = io_ifc_fetch_addr_f[0] ? _T_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_197 | _T_198; // @[Mux.scala 27:72]
  wire [1:0] _T_207 = {tag_match_way1_expanded_p1_f[0],tag_match_way1_expanded_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_208 = _T_143 ? tag_match_way1_expanded_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_209 = io_ifc_fetch_addr_f[0] ? _T_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_208 | _T_209; // @[Mux.scala 27:72]
  wire  _T_211 = bht_valid_f == 2'h0; // @[el2_ifu_bp_ctl.scala 216:47]
  wire [1:0] _GEN_1037 = {{1'd0}, _T_211}; // @[el2_ifu_bp_ctl.scala 216:58]
  wire [1:0] _T_212 = _GEN_1037 & btb_vlru_rd_f; // @[el2_ifu_bp_ctl.scala 216:58]
  wire  _T_213 = io_ifc_fetch_req_f | exu_mp_valid; // @[el2_ifu_bp_ctl.scala 218:75]
  wire [15:0] _T_228 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_229 = btb_sel_f[0] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_230 = _T_228 | _T_229; // @[Mux.scala 27:72]
  wire [16:0] btb_sel_data_f = {{1'd0}, _T_230}; // @[el2_ifu_bp_ctl.scala 231:18]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[el2_ifu_bp_ctl.scala 226:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[el2_ifu_bp_ctl.scala 227:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[el2_ifu_bp_ctl.scala 228:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[el2_ifu_bp_ctl.scala 229:36]
  wire [1:0] _T_278 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_278; // @[el2_ifu_bp_ctl.scala 257:34]
  wire [1:0] _T_232 = bht_valid_f & hist1_raw; // @[el2_ifu_bp_ctl.scala 234:39]
  wire  _T_233 = |_T_232; // @[el2_ifu_bp_ctl.scala 234:52]
  wire  _T_234 = _T_233 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 234:56]
  wire  _T_235 = ~leak_one_f_d1; // @[el2_ifu_bp_ctl.scala 234:79]
  wire  _T_236 = _T_234 & _T_235; // @[el2_ifu_bp_ctl.scala 234:77]
  wire  _T_237 = ~io_dec_tlu_bpred_disable; // @[el2_ifu_bp_ctl.scala 234:96]
  wire  _T_273 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[el2_ifu_bp_ctl.scala 254:51]
  wire  _T_274 = ~io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 254:69]
  wire  _T_284 = bht_valid_f[1] & btb_vbank1_rd_data_f[4]; // @[el2_ifu_bp_ctl.scala 261:34]
  wire  _T_287 = bht_valid_f[0] & btb_vbank0_rd_data_f[4]; // @[el2_ifu_bp_ctl.scala 262:34]
  wire  _T_290 = ~btb_vbank1_rd_data_f[2]; // @[el2_ifu_bp_ctl.scala 264:37]
  wire  _T_291 = bht_valid_f[1] & _T_290; // @[el2_ifu_bp_ctl.scala 264:35]
  wire  _T_293 = _T_291 & btb_vbank1_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 264:65]
  wire  _T_296 = ~btb_vbank0_rd_data_f[2]; // @[el2_ifu_bp_ctl.scala 265:37]
  wire  _T_297 = bht_valid_f[0] & _T_296; // @[el2_ifu_bp_ctl.scala 265:35]
  wire  _T_299 = _T_297 & btb_vbank0_rd_data_f[1]; // @[el2_ifu_bp_ctl.scala 265:65]
  wire [1:0] num_valids = bht_valid_f[1] + bht_valid_f[0]; // @[el2_ifu_bp_ctl.scala 268:35]
  wire [1:0] _T_302 = btb_sel_f & bht_dir_f; // @[el2_ifu_bp_ctl.scala 270:28]
  wire  final_h = &_T_302; // @[el2_ifu_bp_ctl.scala 270:41]
  wire  _T_303 = num_valids == 2'h2; // @[el2_ifu_bp_ctl.scala 274:41]
  wire [7:0] _T_307 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_308 = num_valids == 2'h1; // @[el2_ifu_bp_ctl.scala 275:41]
  wire [7:0] _T_311 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_312 = num_valids == 2'h0; // @[el2_ifu_bp_ctl.scala 276:41]
  wire [7:0] _T_315 = _T_303 ? _T_307 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_316 = _T_308 ? _T_311 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_317 = _T_312 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_318 = _T_315 | _T_316; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_318 | _T_317; // @[Mux.scala 27:72]
  wire  _T_321 = ~exu_flush_final_d1; // @[el2_ifu_bp_ctl.scala 281:27]
  wire  _T_322 = _T_321 & io_ifc_fetch_req_f; // @[el2_ifu_bp_ctl.scala 281:47]
  wire  _T_323 = _T_322 & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 281:68]
  wire  _T_325 = _T_323 & _T_235; // @[el2_ifu_bp_ctl.scala 281:82]
  wire  _T_328 = io_ifc_fetch_req_f & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 282:70]
  wire  _T_330 = _T_328 & _T_235; // @[el2_ifu_bp_ctl.scala 282:84]
  wire  _T_331 = ~_T_330; // @[el2_ifu_bp_ctl.scala 282:49]
  wire  _T_332 = _T_321 & _T_331; // @[el2_ifu_bp_ctl.scala 282:47]
  wire [7:0] _T_334 = exu_flush_final_d1 ? io_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_335 = _T_325 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_336 = _T_332 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_337 = _T_334 | _T_335; // @[Mux.scala 27:72]
  wire [7:0] fghr_ns = _T_337 | _T_336; // @[Mux.scala 27:72]
  wire [1:0] _T_341 = io_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_342 = ~_T_341; // @[el2_ifu_bp_ctl.scala 293:36]
  wire  _T_346 = ~fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 296:36]
  wire  _T_347 = bht_dir_f[0] & _T_346; // @[el2_ifu_bp_ctl.scala 296:34]
  wire  _T_351 = _T_14 & fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 296:72]
  wire  _T_352 = _T_347 | _T_351; // @[el2_ifu_bp_ctl.scala 296:55]
  wire  _T_355 = bht_dir_f[0] & fetch_start_f[0]; // @[el2_ifu_bp_ctl.scala 297:19]
  wire  _T_360 = _T_14 & _T_346; // @[el2_ifu_bp_ctl.scala 297:56]
  wire  _T_361 = _T_355 | _T_360; // @[el2_ifu_bp_ctl.scala 297:39]
  wire [1:0] bloc_f = {_T_352,_T_361}; // @[Cat.scala 29:58]
  wire  _T_365 = _T_14 & io_ifc_fetch_addr_f[0]; // @[el2_ifu_bp_ctl.scala 299:35]
  wire  _T_366 = ~btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 299:62]
  wire  use_fa_plus = _T_365 & _T_366; // @[el2_ifu_bp_ctl.scala 299:60]
  wire  _T_369 = fetch_start_f[0] & btb_sel_f[0]; // @[el2_ifu_bp_ctl.scala 301:44]
  wire  btb_fg_crossing_f = _T_369 & btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 301:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[el2_ifu_bp_ctl.scala 302:43]
  wire  _T_372 = io_ifc_fetch_req_f & _T_274; // @[el2_ifu_bp_ctl.scala 304:87]
  wire  _T_373 = _T_372 & io_ic_hit_f; // @[el2_ifu_bp_ctl.scala 304:112]
  reg [30:0] ifc_fetch_adder_prior; // @[Reg.scala 27:20]
  wire  _T_377 = ~btb_fg_crossing_f; // @[el2_ifu_bp_ctl.scala 309:32]
  wire  _T_378 = ~use_fa_plus; // @[el2_ifu_bp_ctl.scala 309:53]
  wire  _T_379 = _T_377 & _T_378; // @[el2_ifu_bp_ctl.scala 309:51]
  wire [29:0] _T_382 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_383 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 31'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_384 = _T_379 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [30:0] _GEN_1038 = {{1'd0}, _T_382}; // @[Mux.scala 27:72]
  wire [30:0] _T_385 = _GEN_1038 | _T_383; // @[Mux.scala 27:72]
  wire [30:0] _GEN_1039 = {{1'd0}, _T_384}; // @[Mux.scala 27:72]
  wire [30:0] adder_pc_in_f = _T_385 | _GEN_1039; // @[Mux.scala 27:72]
  wire [31:0] _T_389 = {adder_pc_in_f[29:0],bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_390 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_393 = _T_389[12:1] + _T_390[12:1]; // @[el2_lib.scala 198:31]
  wire [18:0] _T_396 = _T_389[31:13] + 19'h1; // @[el2_lib.scala 199:27]
  wire [18:0] _T_399 = _T_389[31:13] - 19'h1; // @[el2_lib.scala 200:27]
  wire  _T_402 = ~_T_393[12]; // @[el2_lib.scala 202:27]
  wire  _T_403 = _T_390[12] ^ _T_402; // @[el2_lib.scala 202:25]
  wire  _T_406 = ~_T_390[12]; // @[el2_lib.scala 203:8]
  wire  _T_408 = _T_406 & _T_393[12]; // @[el2_lib.scala 203:14]
  wire  _T_412 = _T_390[12] & _T_402; // @[el2_lib.scala 204:13]
  wire [18:0] _T_414 = _T_403 ? _T_389[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_415 = _T_408 ? _T_396 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_416 = _T_412 ? _T_399 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_417 = _T_414 | _T_415; // @[Mux.scala 27:72]
  wire [18:0] _T_418 = _T_417 | _T_416; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_418,_T_393[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_422 = ~btb_rd_call_f; // @[el2_ifu_bp_ctl.scala 316:49]
  wire  _T_423 = btb_rd_ret_f & _T_422; // @[el2_ifu_bp_ctl.scala 316:47]
  reg [31:0] rets_out_0; // @[Reg.scala 27:20]
  wire  _T_425 = _T_423 & rets_out_0[0]; // @[el2_ifu_bp_ctl.scala 316:64]
  wire [12:0] _T_436 = {11'h0,_T_366,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_439 = _T_389[12:1] + _T_436[12:1]; // @[el2_lib.scala 198:31]
  wire  _T_448 = ~_T_439[12]; // @[el2_lib.scala 202:27]
  wire  _T_449 = _T_436[12] ^ _T_448; // @[el2_lib.scala 202:25]
  wire  _T_452 = ~_T_436[12]; // @[el2_lib.scala 203:8]
  wire  _T_454 = _T_452 & _T_439[12]; // @[el2_lib.scala 203:14]
  wire  _T_458 = _T_436[12] & _T_448; // @[el2_lib.scala 204:13]
  wire [18:0] _T_460 = _T_449 ? _T_389[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_461 = _T_454 ? _T_396 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_462 = _T_458 ? _T_399 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_463 = _T_460 | _T_461; // @[Mux.scala 27:72]
  wire [18:0] _T_464 = _T_463 | _T_462; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_464,_T_439[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_468 = ~btb_rd_ret_f; // @[el2_ifu_bp_ctl.scala 322:33]
  wire  _T_469 = btb_rd_call_f & _T_468; // @[el2_ifu_bp_ctl.scala 322:31]
  wire  rs_push = _T_469 & io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 322:47]
  wire  rs_pop = _T_423 & io_ifu_bp_hit_taken_f; // @[el2_ifu_bp_ctl.scala 323:46]
  wire  _T_472 = ~rs_push; // @[el2_ifu_bp_ctl.scala 324:17]
  wire  _T_473 = ~rs_pop; // @[el2_ifu_bp_ctl.scala 324:28]
  wire  rs_hold = _T_472 & _T_473; // @[el2_ifu_bp_ctl.scala 324:26]
  wire  rsenable_0 = ~rs_hold; // @[el2_ifu_bp_ctl.scala 326:60]
  wire  rsenable_1 = rs_push | rs_pop; // @[el2_ifu_bp_ctl.scala 326:119]
  wire [31:0] _T_476 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_478 = rs_push ? _T_476 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[Reg.scala 27:20]
  wire [31:0] _T_479 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_0 = _T_478 | _T_479; // @[Mux.scala 27:72]
  wire [31:0] _T_483 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[Reg.scala 27:20]
  wire [31:0] _T_484 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_1 = _T_483 | _T_484; // @[Mux.scala 27:72]
  wire [31:0] _T_488 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[Reg.scala 27:20]
  wire [31:0] _T_489 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_2 = _T_488 | _T_489; // @[Mux.scala 27:72]
  wire [31:0] _T_493 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[Reg.scala 27:20]
  wire [31:0] _T_494 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_3 = _T_493 | _T_494; // @[Mux.scala 27:72]
  wire [31:0] _T_498 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[Reg.scala 27:20]
  wire [31:0] _T_499 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_4 = _T_498 | _T_499; // @[Mux.scala 27:72]
  wire [31:0] _T_503 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[Reg.scala 27:20]
  wire [31:0] _T_504 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_5 = _T_503 | _T_504; // @[Mux.scala 27:72]
  wire [31:0] _T_508 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[Reg.scala 27:20]
  wire [31:0] _T_509 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_6 = _T_508 | _T_509; // @[Mux.scala 27:72]
  wire  _T_527 = ~dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 337:35]
  wire  btb_valid = exu_mp_valid & _T_527; // @[el2_ifu_bp_ctl.scala 337:32]
  wire  _T_528 = io_exu_mp_pkt_pcall | io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 340:89]
  wire  _T_529 = io_exu_mp_pkt_pret | io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 340:113]
  wire [21:0] btb_wr_data = {io_exu_mp_btag,io_exu_mp_pkt_toffset,io_exu_mp_pkt_pc4,io_exu_mp_pkt_boffset,_T_528,_T_529,btb_valid}; // @[Cat.scala 29:58]
  wire  exu_mp_valid_write = exu_mp_valid & io_exu_mp_pkt_ataken; // @[el2_ifu_bp_ctl.scala 341:41]
  wire  _T_536 = _T_175 & exu_mp_valid_write; // @[el2_ifu_bp_ctl.scala 343:39]
  wire  _T_538 = _T_536 & _T_527; // @[el2_ifu_bp_ctl.scala 343:60]
  wire  _T_539 = ~io_dec_tlu_br0_r_pkt_way; // @[el2_ifu_bp_ctl.scala 343:87]
  wire  _T_540 = _T_539 & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 343:104]
  wire  btb_wr_en_way0 = _T_538 | _T_540; // @[el2_ifu_bp_ctl.scala 343:83]
  wire  _T_541 = io_exu_mp_pkt_way & exu_mp_valid_write; // @[el2_ifu_bp_ctl.scala 344:36]
  wire  _T_543 = _T_541 & _T_527; // @[el2_ifu_bp_ctl.scala 344:57]
  wire  _T_544 = io_dec_tlu_br0_r_pkt_way & dec_tlu_error_wb; // @[el2_ifu_bp_ctl.scala 344:98]
  wire  btb_wr_en_way1 = _T_543 | _T_544; // @[el2_ifu_bp_ctl.scala 344:80]
  wire [7:0] btb_wr_addr = dec_tlu_error_wb ? {{1'd0}, btb_error_addr_wb} : io_exu_mp_index; // @[el2_ifu_bp_ctl.scala 346:24]
  wire  middle_of_bank = io_exu_mp_pkt_pc4 ^ io_exu_mp_pkt_boffset; // @[el2_ifu_bp_ctl.scala 347:35]
  wire  _T_546 = ~io_exu_mp_pkt_pcall; // @[el2_ifu_bp_ctl.scala 348:43]
  wire  _T_547 = exu_mp_valid & _T_546; // @[el2_ifu_bp_ctl.scala 348:41]
  wire  _T_548 = ~io_exu_mp_pkt_pret; // @[el2_ifu_bp_ctl.scala 348:58]
  wire  _T_549 = _T_547 & _T_548; // @[el2_ifu_bp_ctl.scala 348:56]
  wire  _T_550 = ~io_exu_mp_pkt_pja; // @[el2_ifu_bp_ctl.scala 348:72]
  wire  _T_551 = _T_549 & _T_550; // @[el2_ifu_bp_ctl.scala 348:70]
  wire [1:0] _T_553 = _T_551 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_554 = ~middle_of_bank; // @[el2_ifu_bp_ctl.scala 348:106]
  wire [1:0] _T_555 = {middle_of_bank,_T_554}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_553 & _T_555; // @[el2_ifu_bp_ctl.scala 348:84]
  wire [1:0] _T_557 = io_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_558 = ~io_dec_tlu_br0_r_pkt_middle; // @[el2_ifu_bp_ctl.scala 349:75]
  wire [1:0] _T_559 = {io_dec_tlu_br0_r_pkt_middle,_T_558}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_557 & _T_559; // @[el2_ifu_bp_ctl.scala 349:46]
  wire [9:0] _T_560 = {io_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr0 = _T_560[9:2] ^ io_exu_mp_eghr; // @[el2_lib.scala 188:35]
  wire [9:0] _T_563 = {io_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_wr_addr2 = _T_563[9:2] ^ io_exu_i0_br_fghr_r; // @[el2_lib.scala 188:35]
  wire  _T_572 = btb_wr_addr == 8'h0; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_573 = _T_572 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_575 = btb_wr_addr == 8'h1; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_576 = _T_575 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_578 = btb_wr_addr == 8'h2; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_579 = _T_578 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_581 = btb_wr_addr == 8'h3; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_582 = _T_581 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_584 = btb_wr_addr == 8'h4; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_585 = _T_584 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_587 = btb_wr_addr == 8'h5; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_588 = _T_587 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_590 = btb_wr_addr == 8'h6; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_591 = _T_590 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_593 = btb_wr_addr == 8'h7; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_594 = _T_593 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_596 = btb_wr_addr == 8'h8; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_597 = _T_596 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_599 = btb_wr_addr == 8'h9; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_600 = _T_599 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_602 = btb_wr_addr == 8'ha; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_603 = _T_602 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_605 = btb_wr_addr == 8'hb; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_606 = _T_605 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_608 = btb_wr_addr == 8'hc; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_609 = _T_608 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_611 = btb_wr_addr == 8'hd; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_612 = _T_611 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_614 = btb_wr_addr == 8'he; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_615 = _T_614 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_617 = btb_wr_addr == 8'hf; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_618 = _T_617 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_620 = btb_wr_addr == 8'h10; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_621 = _T_620 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_623 = btb_wr_addr == 8'h11; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_624 = _T_623 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_626 = btb_wr_addr == 8'h12; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_627 = _T_626 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_629 = btb_wr_addr == 8'h13; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_630 = _T_629 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_632 = btb_wr_addr == 8'h14; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_633 = _T_632 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_635 = btb_wr_addr == 8'h15; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_636 = _T_635 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_638 = btb_wr_addr == 8'h16; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_639 = _T_638 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_641 = btb_wr_addr == 8'h17; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_642 = _T_641 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_644 = btb_wr_addr == 8'h18; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_645 = _T_644 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_647 = btb_wr_addr == 8'h19; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_648 = _T_647 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_650 = btb_wr_addr == 8'h1a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_651 = _T_650 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_653 = btb_wr_addr == 8'h1b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_654 = _T_653 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_656 = btb_wr_addr == 8'h1c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_657 = _T_656 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_659 = btb_wr_addr == 8'h1d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_660 = _T_659 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_662 = btb_wr_addr == 8'h1e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_663 = _T_662 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_665 = btb_wr_addr == 8'h1f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_666 = _T_665 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_668 = btb_wr_addr == 8'h20; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_669 = _T_668 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_671 = btb_wr_addr == 8'h21; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_672 = _T_671 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_674 = btb_wr_addr == 8'h22; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_675 = _T_674 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_677 = btb_wr_addr == 8'h23; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_678 = _T_677 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_680 = btb_wr_addr == 8'h24; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_681 = _T_680 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_683 = btb_wr_addr == 8'h25; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_684 = _T_683 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_686 = btb_wr_addr == 8'h26; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_687 = _T_686 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_689 = btb_wr_addr == 8'h27; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_690 = _T_689 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_692 = btb_wr_addr == 8'h28; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_693 = _T_692 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_695 = btb_wr_addr == 8'h29; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_696 = _T_695 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_698 = btb_wr_addr == 8'h2a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_699 = _T_698 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_701 = btb_wr_addr == 8'h2b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_702 = _T_701 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_704 = btb_wr_addr == 8'h2c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_705 = _T_704 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_707 = btb_wr_addr == 8'h2d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_708 = _T_707 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_710 = btb_wr_addr == 8'h2e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_711 = _T_710 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_713 = btb_wr_addr == 8'h2f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_714 = _T_713 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_716 = btb_wr_addr == 8'h30; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_717 = _T_716 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_719 = btb_wr_addr == 8'h31; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_720 = _T_719 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_722 = btb_wr_addr == 8'h32; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_723 = _T_722 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_725 = btb_wr_addr == 8'h33; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_726 = _T_725 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_728 = btb_wr_addr == 8'h34; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_729 = _T_728 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_731 = btb_wr_addr == 8'h35; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_732 = _T_731 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_734 = btb_wr_addr == 8'h36; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_735 = _T_734 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_737 = btb_wr_addr == 8'h37; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_738 = _T_737 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_740 = btb_wr_addr == 8'h38; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_741 = _T_740 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_743 = btb_wr_addr == 8'h39; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_744 = _T_743 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_746 = btb_wr_addr == 8'h3a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_747 = _T_746 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_749 = btb_wr_addr == 8'h3b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_750 = _T_749 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_752 = btb_wr_addr == 8'h3c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_753 = _T_752 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_755 = btb_wr_addr == 8'h3d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_756 = _T_755 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_758 = btb_wr_addr == 8'h3e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_759 = _T_758 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_761 = btb_wr_addr == 8'h3f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_762 = _T_761 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_764 = btb_wr_addr == 8'h40; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_765 = _T_764 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_767 = btb_wr_addr == 8'h41; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_768 = _T_767 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_770 = btb_wr_addr == 8'h42; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_771 = _T_770 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_773 = btb_wr_addr == 8'h43; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_774 = _T_773 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_776 = btb_wr_addr == 8'h44; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_777 = _T_776 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_779 = btb_wr_addr == 8'h45; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_780 = _T_779 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_782 = btb_wr_addr == 8'h46; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_783 = _T_782 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_785 = btb_wr_addr == 8'h47; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_786 = _T_785 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_788 = btb_wr_addr == 8'h48; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_789 = _T_788 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_791 = btb_wr_addr == 8'h49; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_792 = _T_791 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_794 = btb_wr_addr == 8'h4a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_795 = _T_794 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_797 = btb_wr_addr == 8'h4b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_798 = _T_797 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_800 = btb_wr_addr == 8'h4c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_801 = _T_800 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_803 = btb_wr_addr == 8'h4d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_804 = _T_803 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_806 = btb_wr_addr == 8'h4e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_807 = _T_806 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_809 = btb_wr_addr == 8'h4f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_810 = _T_809 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_812 = btb_wr_addr == 8'h50; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_813 = _T_812 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_815 = btb_wr_addr == 8'h51; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_816 = _T_815 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_818 = btb_wr_addr == 8'h52; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_819 = _T_818 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_821 = btb_wr_addr == 8'h53; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_822 = _T_821 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_824 = btb_wr_addr == 8'h54; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_825 = _T_824 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_827 = btb_wr_addr == 8'h55; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_828 = _T_827 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_830 = btb_wr_addr == 8'h56; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_831 = _T_830 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_833 = btb_wr_addr == 8'h57; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_834 = _T_833 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_836 = btb_wr_addr == 8'h58; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_837 = _T_836 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_839 = btb_wr_addr == 8'h59; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_840 = _T_839 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_842 = btb_wr_addr == 8'h5a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_843 = _T_842 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_845 = btb_wr_addr == 8'h5b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_846 = _T_845 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_848 = btb_wr_addr == 8'h5c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_849 = _T_848 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_851 = btb_wr_addr == 8'h5d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_852 = _T_851 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_854 = btb_wr_addr == 8'h5e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_855 = _T_854 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_857 = btb_wr_addr == 8'h5f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_858 = _T_857 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_860 = btb_wr_addr == 8'h60; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_861 = _T_860 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_863 = btb_wr_addr == 8'h61; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_864 = _T_863 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_866 = btb_wr_addr == 8'h62; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_867 = _T_866 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_869 = btb_wr_addr == 8'h63; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_870 = _T_869 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_872 = btb_wr_addr == 8'h64; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_873 = _T_872 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_875 = btb_wr_addr == 8'h65; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_876 = _T_875 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_878 = btb_wr_addr == 8'h66; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_879 = _T_878 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_881 = btb_wr_addr == 8'h67; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_882 = _T_881 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_884 = btb_wr_addr == 8'h68; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_885 = _T_884 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_887 = btb_wr_addr == 8'h69; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_888 = _T_887 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_890 = btb_wr_addr == 8'h6a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_891 = _T_890 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_893 = btb_wr_addr == 8'h6b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_894 = _T_893 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_896 = btb_wr_addr == 8'h6c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_897 = _T_896 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_899 = btb_wr_addr == 8'h6d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_900 = _T_899 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_902 = btb_wr_addr == 8'h6e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_903 = _T_902 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_905 = btb_wr_addr == 8'h6f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_906 = _T_905 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_908 = btb_wr_addr == 8'h70; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_909 = _T_908 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_911 = btb_wr_addr == 8'h71; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_912 = _T_911 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_914 = btb_wr_addr == 8'h72; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_915 = _T_914 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_917 = btb_wr_addr == 8'h73; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_918 = _T_917 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_920 = btb_wr_addr == 8'h74; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_921 = _T_920 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_923 = btb_wr_addr == 8'h75; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_924 = _T_923 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_926 = btb_wr_addr == 8'h76; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_927 = _T_926 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_929 = btb_wr_addr == 8'h77; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_930 = _T_929 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_932 = btb_wr_addr == 8'h78; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_933 = _T_932 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_935 = btb_wr_addr == 8'h79; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_936 = _T_935 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_938 = btb_wr_addr == 8'h7a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_939 = _T_938 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_941 = btb_wr_addr == 8'h7b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_942 = _T_941 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_944 = btb_wr_addr == 8'h7c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_945 = _T_944 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_947 = btb_wr_addr == 8'h7d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_948 = _T_947 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_950 = btb_wr_addr == 8'h7e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_951 = _T_950 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_953 = btb_wr_addr == 8'h7f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_954 = _T_953 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_956 = btb_wr_addr == 8'h80; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_957 = _T_956 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_959 = btb_wr_addr == 8'h81; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_960 = _T_959 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_962 = btb_wr_addr == 8'h82; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_963 = _T_962 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_965 = btb_wr_addr == 8'h83; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_966 = _T_965 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_968 = btb_wr_addr == 8'h84; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_969 = _T_968 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_971 = btb_wr_addr == 8'h85; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_972 = _T_971 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_974 = btb_wr_addr == 8'h86; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_975 = _T_974 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_977 = btb_wr_addr == 8'h87; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_978 = _T_977 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_980 = btb_wr_addr == 8'h88; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_981 = _T_980 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_983 = btb_wr_addr == 8'h89; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_984 = _T_983 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_986 = btb_wr_addr == 8'h8a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_987 = _T_986 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_989 = btb_wr_addr == 8'h8b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_990 = _T_989 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_992 = btb_wr_addr == 8'h8c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_993 = _T_992 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_995 = btb_wr_addr == 8'h8d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_996 = _T_995 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_998 = btb_wr_addr == 8'h8e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_999 = _T_998 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1001 = btb_wr_addr == 8'h8f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1002 = _T_1001 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1004 = btb_wr_addr == 8'h90; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1005 = _T_1004 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1007 = btb_wr_addr == 8'h91; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1008 = _T_1007 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1010 = btb_wr_addr == 8'h92; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1011 = _T_1010 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1013 = btb_wr_addr == 8'h93; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1014 = _T_1013 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1016 = btb_wr_addr == 8'h94; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1017 = _T_1016 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1019 = btb_wr_addr == 8'h95; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1020 = _T_1019 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1022 = btb_wr_addr == 8'h96; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1023 = _T_1022 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1025 = btb_wr_addr == 8'h97; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1026 = _T_1025 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1028 = btb_wr_addr == 8'h98; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1029 = _T_1028 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1031 = btb_wr_addr == 8'h99; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1032 = _T_1031 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1034 = btb_wr_addr == 8'h9a; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1035 = _T_1034 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1037 = btb_wr_addr == 8'h9b; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1038 = _T_1037 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1040 = btb_wr_addr == 8'h9c; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1041 = _T_1040 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1043 = btb_wr_addr == 8'h9d; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1044 = _T_1043 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1046 = btb_wr_addr == 8'h9e; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1047 = _T_1046 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1049 = btb_wr_addr == 8'h9f; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1050 = _T_1049 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1052 = btb_wr_addr == 8'ha0; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1053 = _T_1052 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1055 = btb_wr_addr == 8'ha1; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1056 = _T_1055 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1058 = btb_wr_addr == 8'ha2; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1059 = _T_1058 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1061 = btb_wr_addr == 8'ha3; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1062 = _T_1061 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1064 = btb_wr_addr == 8'ha4; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1065 = _T_1064 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1067 = btb_wr_addr == 8'ha5; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1068 = _T_1067 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1070 = btb_wr_addr == 8'ha6; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1071 = _T_1070 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1073 = btb_wr_addr == 8'ha7; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1074 = _T_1073 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1076 = btb_wr_addr == 8'ha8; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1077 = _T_1076 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1079 = btb_wr_addr == 8'ha9; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1080 = _T_1079 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1082 = btb_wr_addr == 8'haa; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1083 = _T_1082 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1085 = btb_wr_addr == 8'hab; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1086 = _T_1085 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1088 = btb_wr_addr == 8'hac; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1089 = _T_1088 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1091 = btb_wr_addr == 8'had; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1092 = _T_1091 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1094 = btb_wr_addr == 8'hae; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1095 = _T_1094 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1097 = btb_wr_addr == 8'haf; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1098 = _T_1097 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1100 = btb_wr_addr == 8'hb0; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1101 = _T_1100 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1103 = btb_wr_addr == 8'hb1; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1104 = _T_1103 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1106 = btb_wr_addr == 8'hb2; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1107 = _T_1106 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1109 = btb_wr_addr == 8'hb3; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1110 = _T_1109 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1112 = btb_wr_addr == 8'hb4; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1113 = _T_1112 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1115 = btb_wr_addr == 8'hb5; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1116 = _T_1115 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1118 = btb_wr_addr == 8'hb6; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1119 = _T_1118 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1121 = btb_wr_addr == 8'hb7; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1122 = _T_1121 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1124 = btb_wr_addr == 8'hb8; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1125 = _T_1124 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1127 = btb_wr_addr == 8'hb9; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1128 = _T_1127 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1130 = btb_wr_addr == 8'hba; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1131 = _T_1130 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1133 = btb_wr_addr == 8'hbb; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1134 = _T_1133 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1136 = btb_wr_addr == 8'hbc; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1137 = _T_1136 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1139 = btb_wr_addr == 8'hbd; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1140 = _T_1139 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1142 = btb_wr_addr == 8'hbe; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1143 = _T_1142 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1145 = btb_wr_addr == 8'hbf; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1146 = _T_1145 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1148 = btb_wr_addr == 8'hc0; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1149 = _T_1148 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1151 = btb_wr_addr == 8'hc1; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1152 = _T_1151 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1154 = btb_wr_addr == 8'hc2; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1155 = _T_1154 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1157 = btb_wr_addr == 8'hc3; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1158 = _T_1157 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1160 = btb_wr_addr == 8'hc4; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1161 = _T_1160 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1163 = btb_wr_addr == 8'hc5; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1164 = _T_1163 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1166 = btb_wr_addr == 8'hc6; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1167 = _T_1166 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1169 = btb_wr_addr == 8'hc7; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1170 = _T_1169 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1172 = btb_wr_addr == 8'hc8; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1173 = _T_1172 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1175 = btb_wr_addr == 8'hc9; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1176 = _T_1175 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1178 = btb_wr_addr == 8'hca; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1179 = _T_1178 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1181 = btb_wr_addr == 8'hcb; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1182 = _T_1181 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1184 = btb_wr_addr == 8'hcc; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1185 = _T_1184 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1187 = btb_wr_addr == 8'hcd; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1188 = _T_1187 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1190 = btb_wr_addr == 8'hce; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1191 = _T_1190 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1193 = btb_wr_addr == 8'hcf; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1194 = _T_1193 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1196 = btb_wr_addr == 8'hd0; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1197 = _T_1196 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1199 = btb_wr_addr == 8'hd1; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1200 = _T_1199 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1202 = btb_wr_addr == 8'hd2; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1203 = _T_1202 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1205 = btb_wr_addr == 8'hd3; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1206 = _T_1205 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1208 = btb_wr_addr == 8'hd4; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1209 = _T_1208 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1211 = btb_wr_addr == 8'hd5; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1212 = _T_1211 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1214 = btb_wr_addr == 8'hd6; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1215 = _T_1214 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1217 = btb_wr_addr == 8'hd7; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1218 = _T_1217 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1220 = btb_wr_addr == 8'hd8; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1221 = _T_1220 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1223 = btb_wr_addr == 8'hd9; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1224 = _T_1223 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1226 = btb_wr_addr == 8'hda; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1227 = _T_1226 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1229 = btb_wr_addr == 8'hdb; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1230 = _T_1229 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1232 = btb_wr_addr == 8'hdc; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1233 = _T_1232 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1235 = btb_wr_addr == 8'hdd; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1236 = _T_1235 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1238 = btb_wr_addr == 8'hde; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1239 = _T_1238 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1241 = btb_wr_addr == 8'hdf; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1242 = _T_1241 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1244 = btb_wr_addr == 8'he0; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1245 = _T_1244 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1247 = btb_wr_addr == 8'he1; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1248 = _T_1247 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1250 = btb_wr_addr == 8'he2; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1251 = _T_1250 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1253 = btb_wr_addr == 8'he3; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1254 = _T_1253 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1256 = btb_wr_addr == 8'he4; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1257 = _T_1256 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1259 = btb_wr_addr == 8'he5; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1260 = _T_1259 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1262 = btb_wr_addr == 8'he6; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1263 = _T_1262 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1265 = btb_wr_addr == 8'he7; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1266 = _T_1265 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1268 = btb_wr_addr == 8'he8; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1269 = _T_1268 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1271 = btb_wr_addr == 8'he9; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1272 = _T_1271 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1274 = btb_wr_addr == 8'hea; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1275 = _T_1274 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1277 = btb_wr_addr == 8'heb; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1278 = _T_1277 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1280 = btb_wr_addr == 8'hec; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1281 = _T_1280 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1283 = btb_wr_addr == 8'hed; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1284 = _T_1283 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1286 = btb_wr_addr == 8'hee; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1287 = _T_1286 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1289 = btb_wr_addr == 8'hef; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1290 = _T_1289 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1292 = btb_wr_addr == 8'hf0; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1293 = _T_1292 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1295 = btb_wr_addr == 8'hf1; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1296 = _T_1295 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1298 = btb_wr_addr == 8'hf2; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1299 = _T_1298 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1301 = btb_wr_addr == 8'hf3; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1302 = _T_1301 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1304 = btb_wr_addr == 8'hf4; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1305 = _T_1304 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1307 = btb_wr_addr == 8'hf5; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1308 = _T_1307 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1310 = btb_wr_addr == 8'hf6; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1311 = _T_1310 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1313 = btb_wr_addr == 8'hf7; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1314 = _T_1313 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1316 = btb_wr_addr == 8'hf8; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1317 = _T_1316 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1319 = btb_wr_addr == 8'hf9; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1320 = _T_1319 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1322 = btb_wr_addr == 8'hfa; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1323 = _T_1322 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1325 = btb_wr_addr == 8'hfb; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1326 = _T_1325 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1328 = btb_wr_addr == 8'hfc; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1329 = _T_1328 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1331 = btb_wr_addr == 8'hfd; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1332 = _T_1331 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1334 = btb_wr_addr == 8'hfe; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1335 = _T_1334 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1337 = btb_wr_addr == 8'hff; // @[el2_ifu_bp_ctl.scala 366:101]
  wire  _T_1338 = _T_1337 & btb_wr_en_way0; // @[el2_ifu_bp_ctl.scala 366:109]
  wire  _T_1341 = _T_572 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1344 = _T_575 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1347 = _T_578 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1350 = _T_581 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1353 = _T_584 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1356 = _T_587 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1359 = _T_590 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1362 = _T_593 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1365 = _T_596 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1368 = _T_599 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1371 = _T_602 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1374 = _T_605 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1377 = _T_608 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1380 = _T_611 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1383 = _T_614 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1386 = _T_617 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1389 = _T_620 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1392 = _T_623 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1395 = _T_626 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1398 = _T_629 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1401 = _T_632 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1404 = _T_635 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1407 = _T_638 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1410 = _T_641 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1413 = _T_644 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1416 = _T_647 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1419 = _T_650 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1422 = _T_653 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1425 = _T_656 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1428 = _T_659 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1431 = _T_662 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1434 = _T_665 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1437 = _T_668 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1440 = _T_671 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1443 = _T_674 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1446 = _T_677 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1449 = _T_680 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1452 = _T_683 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1455 = _T_686 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1458 = _T_689 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1461 = _T_692 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1464 = _T_695 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1467 = _T_698 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1470 = _T_701 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1473 = _T_704 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1476 = _T_707 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1479 = _T_710 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1482 = _T_713 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1485 = _T_716 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1488 = _T_719 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1491 = _T_722 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1494 = _T_725 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1497 = _T_728 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1500 = _T_731 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1503 = _T_734 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1506 = _T_737 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1509 = _T_740 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1512 = _T_743 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1515 = _T_746 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1518 = _T_749 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1521 = _T_752 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1524 = _T_755 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1527 = _T_758 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1530 = _T_761 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1533 = _T_764 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1536 = _T_767 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1539 = _T_770 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1542 = _T_773 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1545 = _T_776 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1548 = _T_779 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1551 = _T_782 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1554 = _T_785 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1557 = _T_788 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1560 = _T_791 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1563 = _T_794 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1566 = _T_797 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1569 = _T_800 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1572 = _T_803 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1575 = _T_806 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1578 = _T_809 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1581 = _T_812 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1584 = _T_815 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1587 = _T_818 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1590 = _T_821 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1593 = _T_824 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1596 = _T_827 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1599 = _T_830 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1602 = _T_833 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1605 = _T_836 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1608 = _T_839 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1611 = _T_842 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1614 = _T_845 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1617 = _T_848 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1620 = _T_851 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1623 = _T_854 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1626 = _T_857 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1629 = _T_860 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1632 = _T_863 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1635 = _T_866 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1638 = _T_869 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1641 = _T_872 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1644 = _T_875 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1647 = _T_878 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1650 = _T_881 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1653 = _T_884 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1656 = _T_887 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1659 = _T_890 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1662 = _T_893 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1665 = _T_896 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1668 = _T_899 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1671 = _T_902 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1674 = _T_905 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1677 = _T_908 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1680 = _T_911 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1683 = _T_914 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1686 = _T_917 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1689 = _T_920 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1692 = _T_923 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1695 = _T_926 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1698 = _T_929 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1701 = _T_932 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1704 = _T_935 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1707 = _T_938 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1710 = _T_941 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1713 = _T_944 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1716 = _T_947 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1719 = _T_950 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1722 = _T_953 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1725 = _T_956 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1728 = _T_959 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1731 = _T_962 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1734 = _T_965 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1737 = _T_968 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1740 = _T_971 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1743 = _T_974 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1746 = _T_977 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1749 = _T_980 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1752 = _T_983 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1755 = _T_986 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1758 = _T_989 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1761 = _T_992 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1764 = _T_995 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1767 = _T_998 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1770 = _T_1001 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1773 = _T_1004 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1776 = _T_1007 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1779 = _T_1010 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1782 = _T_1013 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1785 = _T_1016 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1788 = _T_1019 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1791 = _T_1022 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1794 = _T_1025 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1797 = _T_1028 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1800 = _T_1031 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1803 = _T_1034 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1806 = _T_1037 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1809 = _T_1040 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1812 = _T_1043 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1815 = _T_1046 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1818 = _T_1049 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1821 = _T_1052 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1824 = _T_1055 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1827 = _T_1058 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1830 = _T_1061 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1833 = _T_1064 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1836 = _T_1067 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1839 = _T_1070 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1842 = _T_1073 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1845 = _T_1076 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1848 = _T_1079 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1851 = _T_1082 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1854 = _T_1085 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1857 = _T_1088 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1860 = _T_1091 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1863 = _T_1094 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1866 = _T_1097 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1869 = _T_1100 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1872 = _T_1103 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1875 = _T_1106 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1878 = _T_1109 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1881 = _T_1112 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1884 = _T_1115 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1887 = _T_1118 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1890 = _T_1121 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1893 = _T_1124 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1896 = _T_1127 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1899 = _T_1130 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1902 = _T_1133 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1905 = _T_1136 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1908 = _T_1139 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1911 = _T_1142 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1914 = _T_1145 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1917 = _T_1148 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1920 = _T_1151 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1923 = _T_1154 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1926 = _T_1157 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1929 = _T_1160 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1932 = _T_1163 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1935 = _T_1166 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1938 = _T_1169 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1941 = _T_1172 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1944 = _T_1175 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1947 = _T_1178 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1950 = _T_1181 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1953 = _T_1184 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1956 = _T_1187 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1959 = _T_1190 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1962 = _T_1193 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1965 = _T_1196 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1968 = _T_1199 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1971 = _T_1202 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1974 = _T_1205 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1977 = _T_1208 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1980 = _T_1211 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1983 = _T_1214 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1986 = _T_1217 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1989 = _T_1220 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1992 = _T_1223 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1995 = _T_1226 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_1998 = _T_1229 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2001 = _T_1232 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2004 = _T_1235 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2007 = _T_1238 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2010 = _T_1241 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2013 = _T_1244 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2016 = _T_1247 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2019 = _T_1250 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2022 = _T_1253 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2025 = _T_1256 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2028 = _T_1259 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2031 = _T_1262 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2034 = _T_1265 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2037 = _T_1268 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2040 = _T_1271 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2043 = _T_1274 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2046 = _T_1277 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2049 = _T_1280 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2052 = _T_1283 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2055 = _T_1286 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2058 = _T_1289 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2061 = _T_1292 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2064 = _T_1295 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2067 = _T_1298 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2070 = _T_1301 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2073 = _T_1304 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2076 = _T_1307 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2079 = _T_1310 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2082 = _T_1313 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2085 = _T_1316 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2088 = _T_1319 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2091 = _T_1322 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2094 = _T_1325 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2097 = _T_1328 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2100 = _T_1331 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2103 = _T_1334 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_2106 = _T_1337 & btb_wr_en_way1; // @[el2_ifu_bp_ctl.scala 367:109]
  wire  _T_6206 = bht_wr_addr2[3:0] == 4'h0; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6207 = bht_wr_en2[0] & _T_6206; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6209 = ~bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_6210 = _T_6207 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6215 = bht_wr_addr2[3:0] == 4'h1; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6216 = bht_wr_en2[0] & _T_6215; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6219 = _T_6216 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6224 = bht_wr_addr2[3:0] == 4'h2; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6225 = bht_wr_en2[0] & _T_6224; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6228 = _T_6225 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6233 = bht_wr_addr2[3:0] == 4'h3; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6234 = bht_wr_en2[0] & _T_6233; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6237 = _T_6234 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6242 = bht_wr_addr2[3:0] == 4'h4; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6243 = bht_wr_en2[0] & _T_6242; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6246 = _T_6243 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6251 = bht_wr_addr2[3:0] == 4'h5; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6252 = bht_wr_en2[0] & _T_6251; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6255 = _T_6252 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6260 = bht_wr_addr2[3:0] == 4'h6; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6261 = bht_wr_en2[0] & _T_6260; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6264 = _T_6261 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6269 = bht_wr_addr2[3:0] == 4'h7; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6270 = bht_wr_en2[0] & _T_6269; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6273 = _T_6270 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6278 = bht_wr_addr2[3:0] == 4'h8; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6279 = bht_wr_en2[0] & _T_6278; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6282 = _T_6279 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6287 = bht_wr_addr2[3:0] == 4'h9; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6288 = bht_wr_en2[0] & _T_6287; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6291 = _T_6288 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6296 = bht_wr_addr2[3:0] == 4'ha; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6297 = bht_wr_en2[0] & _T_6296; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6300 = _T_6297 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6305 = bht_wr_addr2[3:0] == 4'hb; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6306 = bht_wr_en2[0] & _T_6305; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6309 = _T_6306 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6314 = bht_wr_addr2[3:0] == 4'hc; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6315 = bht_wr_en2[0] & _T_6314; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6318 = _T_6315 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6323 = bht_wr_addr2[3:0] == 4'hd; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6324 = bht_wr_en2[0] & _T_6323; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6327 = _T_6324 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6332 = bht_wr_addr2[3:0] == 4'he; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6333 = bht_wr_en2[0] & _T_6332; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6336 = _T_6333 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6341 = bht_wr_addr2[3:0] == 4'hf; // @[el2_ifu_bp_ctl.scala 376:74]
  wire  _T_6342 = bht_wr_en2[0] & _T_6341; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_6345 = _T_6342 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6354 = _T_6207 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6363 = _T_6216 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6372 = _T_6225 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6381 = _T_6234 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6390 = _T_6243 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6399 = _T_6252 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6408 = _T_6261 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6417 = _T_6270 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6426 = _T_6279 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6435 = _T_6288 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6444 = _T_6297 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6453 = _T_6306 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6462 = _T_6315 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6471 = _T_6324 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6480 = _T_6333 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6489 = _T_6342 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire [1:0] _GEN_1040 = {{1'd0}, bht_wr_addr2[4]}; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_6497 = _GEN_1040 == 2'h2; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_6498 = _T_6207 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6507 = _T_6216 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6516 = _T_6225 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6525 = _T_6234 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6534 = _T_6243 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6543 = _T_6252 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6552 = _T_6261 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6561 = _T_6270 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6570 = _T_6279 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6579 = _T_6288 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6588 = _T_6297 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6597 = _T_6306 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6606 = _T_6315 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6615 = _T_6324 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6624 = _T_6333 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6633 = _T_6342 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6641 = _GEN_1040 == 2'h3; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_6642 = _T_6207 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6651 = _T_6216 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6660 = _T_6225 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6669 = _T_6234 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6678 = _T_6243 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6687 = _T_6252 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6696 = _T_6261 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6705 = _T_6270 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6714 = _T_6279 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6723 = _T_6288 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6732 = _T_6297 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6741 = _T_6306 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6750 = _T_6315 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6759 = _T_6324 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6768 = _T_6333 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6777 = _T_6342 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire [2:0] _GEN_1072 = {{2'd0}, bht_wr_addr2[4]}; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_6785 = _GEN_1072 == 3'h4; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_6786 = _T_6207 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6795 = _T_6216 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6804 = _T_6225 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6813 = _T_6234 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6822 = _T_6243 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6831 = _T_6252 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6840 = _T_6261 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6849 = _T_6270 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6858 = _T_6279 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6867 = _T_6288 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6876 = _T_6297 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6885 = _T_6306 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6894 = _T_6315 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6903 = _T_6324 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6912 = _T_6333 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6921 = _T_6342 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6929 = _GEN_1072 == 3'h5; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_6930 = _T_6207 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6939 = _T_6216 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6948 = _T_6225 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6957 = _T_6234 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6966 = _T_6243 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6975 = _T_6252 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6984 = _T_6261 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_6993 = _T_6270 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7002 = _T_6279 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7011 = _T_6288 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7020 = _T_6297 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7029 = _T_6306 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7038 = _T_6315 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7047 = _T_6324 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7056 = _T_6333 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7065 = _T_6342 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7073 = _GEN_1072 == 3'h6; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7074 = _T_6207 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7083 = _T_6216 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7092 = _T_6225 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7101 = _T_6234 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7110 = _T_6243 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7119 = _T_6252 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7128 = _T_6261 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7137 = _T_6270 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7146 = _T_6279 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7155 = _T_6288 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7164 = _T_6297 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7173 = _T_6306 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7182 = _T_6315 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7191 = _T_6324 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7200 = _T_6333 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7209 = _T_6342 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7217 = _GEN_1072 == 3'h7; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7218 = _T_6207 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7227 = _T_6216 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7236 = _T_6225 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7245 = _T_6234 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7254 = _T_6243 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7263 = _T_6252 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7272 = _T_6261 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7281 = _T_6270 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7290 = _T_6279 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7299 = _T_6288 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7308 = _T_6297 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7317 = _T_6306 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7326 = _T_6315 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7335 = _T_6324 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7344 = _T_6333 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7353 = _T_6342 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire [3:0] _GEN_1136 = {{3'd0}, bht_wr_addr2[4]}; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7361 = _GEN_1136 == 4'h8; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7362 = _T_6207 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7371 = _T_6216 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7380 = _T_6225 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7389 = _T_6234 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7398 = _T_6243 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7407 = _T_6252 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7416 = _T_6261 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7425 = _T_6270 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7434 = _T_6279 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7443 = _T_6288 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7452 = _T_6297 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7461 = _T_6306 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7470 = _T_6315 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7479 = _T_6324 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7488 = _T_6333 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7497 = _T_6342 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7505 = _GEN_1136 == 4'h9; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7506 = _T_6207 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7515 = _T_6216 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7524 = _T_6225 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7533 = _T_6234 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7542 = _T_6243 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7551 = _T_6252 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7560 = _T_6261 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7569 = _T_6270 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7578 = _T_6279 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7587 = _T_6288 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7596 = _T_6297 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7605 = _T_6306 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7614 = _T_6315 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7623 = _T_6324 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7632 = _T_6333 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7641 = _T_6342 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7649 = _GEN_1136 == 4'ha; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7650 = _T_6207 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7659 = _T_6216 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7668 = _T_6225 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7677 = _T_6234 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7686 = _T_6243 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7695 = _T_6252 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7704 = _T_6261 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7713 = _T_6270 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7722 = _T_6279 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7731 = _T_6288 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7740 = _T_6297 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7749 = _T_6306 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7758 = _T_6315 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7767 = _T_6324 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7776 = _T_6333 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7785 = _T_6342 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7793 = _GEN_1136 == 4'hb; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7794 = _T_6207 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7803 = _T_6216 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7812 = _T_6225 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7821 = _T_6234 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7830 = _T_6243 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7839 = _T_6252 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7848 = _T_6261 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7857 = _T_6270 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7866 = _T_6279 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7875 = _T_6288 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7884 = _T_6297 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7893 = _T_6306 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7902 = _T_6315 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7911 = _T_6324 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7920 = _T_6333 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7929 = _T_6342 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7937 = _GEN_1136 == 4'hc; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_7938 = _T_6207 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7947 = _T_6216 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7956 = _T_6225 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7965 = _T_6234 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7974 = _T_6243 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7983 = _T_6252 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_7992 = _T_6261 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8001 = _T_6270 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8010 = _T_6279 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8019 = _T_6288 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8028 = _T_6297 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8037 = _T_6306 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8046 = _T_6315 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8055 = _T_6324 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8064 = _T_6333 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8073 = _T_6342 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8081 = _GEN_1136 == 4'hd; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_8082 = _T_6207 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8091 = _T_6216 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8100 = _T_6225 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8109 = _T_6234 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8118 = _T_6243 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8127 = _T_6252 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8136 = _T_6261 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8145 = _T_6270 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8154 = _T_6279 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8163 = _T_6288 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8172 = _T_6297 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8181 = _T_6306 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8190 = _T_6315 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8199 = _T_6324 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8208 = _T_6333 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8217 = _T_6342 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8225 = _GEN_1136 == 4'he; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_8226 = _T_6207 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8235 = _T_6216 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8244 = _T_6225 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8253 = _T_6234 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8262 = _T_6243 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8271 = _T_6252 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8280 = _T_6261 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8289 = _T_6270 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8298 = _T_6279 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8307 = _T_6288 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8316 = _T_6297 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8325 = _T_6306 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8334 = _T_6315 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8343 = _T_6324 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8352 = _T_6333 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8361 = _T_6342 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8369 = _GEN_1136 == 4'hf; // @[el2_ifu_bp_ctl.scala 376:171]
  wire  _T_8370 = _T_6207 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8379 = _T_6216 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8388 = _T_6225 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8397 = _T_6234 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8406 = _T_6243 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8415 = _T_6252 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8424 = _T_6261 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8433 = _T_6270 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8442 = _T_6279 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8451 = _T_6288 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8460 = _T_6297 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8469 = _T_6306 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8478 = _T_6315 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8487 = _T_6324 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8496 = _T_6333 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8505 = _T_6342 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8511 = bht_wr_en2[1] & _T_6206; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8514 = _T_8511 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8520 = bht_wr_en2[1] & _T_6215; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8523 = _T_8520 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8529 = bht_wr_en2[1] & _T_6224; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8532 = _T_8529 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8538 = bht_wr_en2[1] & _T_6233; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8541 = _T_8538 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8547 = bht_wr_en2[1] & _T_6242; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8550 = _T_8547 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8556 = bht_wr_en2[1] & _T_6251; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8559 = _T_8556 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8565 = bht_wr_en2[1] & _T_6260; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8568 = _T_8565 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8574 = bht_wr_en2[1] & _T_6269; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8577 = _T_8574 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8583 = bht_wr_en2[1] & _T_6278; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8586 = _T_8583 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8592 = bht_wr_en2[1] & _T_6287; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8595 = _T_8592 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8601 = bht_wr_en2[1] & _T_6296; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8604 = _T_8601 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8610 = bht_wr_en2[1] & _T_6305; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8613 = _T_8610 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8619 = bht_wr_en2[1] & _T_6314; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8622 = _T_8619 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8628 = bht_wr_en2[1] & _T_6323; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8631 = _T_8628 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8637 = bht_wr_en2[1] & _T_6332; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8640 = _T_8637 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8646 = bht_wr_en2[1] & _T_6341; // @[el2_ifu_bp_ctl.scala 376:23]
  wire  _T_8649 = _T_8646 & _T_6209; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8658 = _T_8511 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8667 = _T_8520 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8676 = _T_8529 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8685 = _T_8538 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8694 = _T_8547 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8703 = _T_8556 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8712 = _T_8565 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8721 = _T_8574 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8730 = _T_8583 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8739 = _T_8592 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8748 = _T_8601 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8757 = _T_8610 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8766 = _T_8619 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8775 = _T_8628 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8784 = _T_8637 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8793 = _T_8646 & bht_wr_addr2[4]; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8802 = _T_8511 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8811 = _T_8520 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8820 = _T_8529 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8829 = _T_8538 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8838 = _T_8547 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8847 = _T_8556 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8856 = _T_8565 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8865 = _T_8574 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8874 = _T_8583 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8883 = _T_8592 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8892 = _T_8601 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8901 = _T_8610 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8910 = _T_8619 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8919 = _T_8628 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8928 = _T_8637 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8937 = _T_8646 & _T_6497; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8946 = _T_8511 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8955 = _T_8520 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8964 = _T_8529 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8973 = _T_8538 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8982 = _T_8547 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_8991 = _T_8556 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9000 = _T_8565 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9009 = _T_8574 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9018 = _T_8583 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9027 = _T_8592 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9036 = _T_8601 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9045 = _T_8610 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9054 = _T_8619 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9063 = _T_8628 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9072 = _T_8637 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9081 = _T_8646 & _T_6641; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9090 = _T_8511 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9099 = _T_8520 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9108 = _T_8529 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9117 = _T_8538 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9126 = _T_8547 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9135 = _T_8556 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9144 = _T_8565 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9153 = _T_8574 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9162 = _T_8583 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9171 = _T_8592 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9180 = _T_8601 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9189 = _T_8610 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9198 = _T_8619 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9207 = _T_8628 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9216 = _T_8637 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9225 = _T_8646 & _T_6785; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9234 = _T_8511 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9243 = _T_8520 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9252 = _T_8529 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9261 = _T_8538 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9270 = _T_8547 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9279 = _T_8556 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9288 = _T_8565 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9297 = _T_8574 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9306 = _T_8583 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9315 = _T_8592 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9324 = _T_8601 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9333 = _T_8610 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9342 = _T_8619 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9351 = _T_8628 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9360 = _T_8637 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9369 = _T_8646 & _T_6929; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9378 = _T_8511 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9387 = _T_8520 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9396 = _T_8529 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9405 = _T_8538 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9414 = _T_8547 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9423 = _T_8556 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9432 = _T_8565 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9441 = _T_8574 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9450 = _T_8583 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9459 = _T_8592 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9468 = _T_8601 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9477 = _T_8610 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9486 = _T_8619 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9495 = _T_8628 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9504 = _T_8637 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9513 = _T_8646 & _T_7073; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9522 = _T_8511 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9531 = _T_8520 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9540 = _T_8529 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9549 = _T_8538 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9558 = _T_8547 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9567 = _T_8556 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9576 = _T_8565 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9585 = _T_8574 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9594 = _T_8583 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9603 = _T_8592 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9612 = _T_8601 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9621 = _T_8610 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9630 = _T_8619 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9639 = _T_8628 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9648 = _T_8637 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9657 = _T_8646 & _T_7217; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9666 = _T_8511 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9675 = _T_8520 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9684 = _T_8529 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9693 = _T_8538 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9702 = _T_8547 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9711 = _T_8556 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9720 = _T_8565 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9729 = _T_8574 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9738 = _T_8583 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9747 = _T_8592 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9756 = _T_8601 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9765 = _T_8610 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9774 = _T_8619 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9783 = _T_8628 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9792 = _T_8637 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9801 = _T_8646 & _T_7361; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9810 = _T_8511 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9819 = _T_8520 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9828 = _T_8529 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9837 = _T_8538 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9846 = _T_8547 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9855 = _T_8556 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9864 = _T_8565 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9873 = _T_8574 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9882 = _T_8583 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9891 = _T_8592 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9900 = _T_8601 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9909 = _T_8610 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9918 = _T_8619 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9927 = _T_8628 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9936 = _T_8637 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9945 = _T_8646 & _T_7505; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9954 = _T_8511 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9963 = _T_8520 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9972 = _T_8529 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9981 = _T_8538 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9990 = _T_8547 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_9999 = _T_8556 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10008 = _T_8565 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10017 = _T_8574 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10026 = _T_8583 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10035 = _T_8592 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10044 = _T_8601 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10053 = _T_8610 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10062 = _T_8619 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10071 = _T_8628 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10080 = _T_8637 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10089 = _T_8646 & _T_7649; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10098 = _T_8511 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10107 = _T_8520 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10116 = _T_8529 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10125 = _T_8538 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10134 = _T_8547 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10143 = _T_8556 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10152 = _T_8565 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10161 = _T_8574 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10170 = _T_8583 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10179 = _T_8592 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10188 = _T_8601 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10197 = _T_8610 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10206 = _T_8619 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10215 = _T_8628 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10224 = _T_8637 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10233 = _T_8646 & _T_7793; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10242 = _T_8511 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10251 = _T_8520 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10260 = _T_8529 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10269 = _T_8538 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10278 = _T_8547 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10287 = _T_8556 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10296 = _T_8565 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10305 = _T_8574 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10314 = _T_8583 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10323 = _T_8592 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10332 = _T_8601 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10341 = _T_8610 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10350 = _T_8619 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10359 = _T_8628 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10368 = _T_8637 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10377 = _T_8646 & _T_7937; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10386 = _T_8511 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10395 = _T_8520 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10404 = _T_8529 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10413 = _T_8538 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10422 = _T_8547 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10431 = _T_8556 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10440 = _T_8565 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10449 = _T_8574 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10458 = _T_8583 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10467 = _T_8592 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10476 = _T_8601 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10485 = _T_8610 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10494 = _T_8619 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10503 = _T_8628 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10512 = _T_8637 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10521 = _T_8646 & _T_8081; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10530 = _T_8511 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10539 = _T_8520 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10548 = _T_8529 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10557 = _T_8538 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10566 = _T_8547 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10575 = _T_8556 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10584 = _T_8565 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10593 = _T_8574 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10602 = _T_8583 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10611 = _T_8592 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10620 = _T_8601 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10629 = _T_8610 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10638 = _T_8619 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10647 = _T_8628 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10656 = _T_8637 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10665 = _T_8646 & _T_8225; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10674 = _T_8511 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10683 = _T_8520 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10692 = _T_8529 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10701 = _T_8538 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10710 = _T_8547 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10719 = _T_8556 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10728 = _T_8565 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10737 = _T_8574 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10746 = _T_8583 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10755 = _T_8592 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10764 = _T_8601 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10773 = _T_8610 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10782 = _T_8619 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10791 = _T_8628 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10800 = _T_8637 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10809 = _T_8646 & _T_8369; // @[el2_ifu_bp_ctl.scala 376:86]
  wire  _T_10814 = bht_wr_addr0[3:0] == 4'h0; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10815 = bht_wr_en0[0] & _T_10814; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10817 = ~bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_10818 = _T_10815 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_0 = _T_10818 | _T_6210; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10830 = bht_wr_addr0[3:0] == 4'h1; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10831 = bht_wr_en0[0] & _T_10830; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10834 = _T_10831 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_1 = _T_10834 | _T_6219; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10846 = bht_wr_addr0[3:0] == 4'h2; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10847 = bht_wr_en0[0] & _T_10846; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10850 = _T_10847 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_2 = _T_10850 | _T_6228; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10862 = bht_wr_addr0[3:0] == 4'h3; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10863 = bht_wr_en0[0] & _T_10862; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10866 = _T_10863 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_3 = _T_10866 | _T_6237; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10878 = bht_wr_addr0[3:0] == 4'h4; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10879 = bht_wr_en0[0] & _T_10878; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10882 = _T_10879 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_4 = _T_10882 | _T_6246; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10894 = bht_wr_addr0[3:0] == 4'h5; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10895 = bht_wr_en0[0] & _T_10894; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10898 = _T_10895 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_5 = _T_10898 | _T_6255; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10910 = bht_wr_addr0[3:0] == 4'h6; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10911 = bht_wr_en0[0] & _T_10910; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10914 = _T_10911 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_6 = _T_10914 | _T_6264; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10926 = bht_wr_addr0[3:0] == 4'h7; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10927 = bht_wr_en0[0] & _T_10926; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10930 = _T_10927 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_7 = _T_10930 | _T_6273; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10942 = bht_wr_addr0[3:0] == 4'h8; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10943 = bht_wr_en0[0] & _T_10942; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10946 = _T_10943 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_8 = _T_10946 | _T_6282; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10958 = bht_wr_addr0[3:0] == 4'h9; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10959 = bht_wr_en0[0] & _T_10958; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10962 = _T_10959 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_9 = _T_10962 | _T_6291; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10974 = bht_wr_addr0[3:0] == 4'ha; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10975 = bht_wr_en0[0] & _T_10974; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10978 = _T_10975 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_10 = _T_10978 | _T_6300; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_10990 = bht_wr_addr0[3:0] == 4'hb; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_10991 = bht_wr_en0[0] & _T_10990; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_10994 = _T_10991 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_11 = _T_10994 | _T_6309; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11006 = bht_wr_addr0[3:0] == 4'hc; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_11007 = bht_wr_en0[0] & _T_11006; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_11010 = _T_11007 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_12 = _T_11010 | _T_6318; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11022 = bht_wr_addr0[3:0] == 4'hd; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_11023 = bht_wr_en0[0] & _T_11022; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_11026 = _T_11023 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_13 = _T_11026 | _T_6327; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11038 = bht_wr_addr0[3:0] == 4'he; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_11039 = bht_wr_en0[0] & _T_11038; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_11042 = _T_11039 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_14 = _T_11042 | _T_6336; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11054 = bht_wr_addr0[3:0] == 4'hf; // @[el2_ifu_bp_ctl.scala 379:69]
  wire  _T_11055 = bht_wr_en0[0] & _T_11054; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_11058 = _T_11055 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_0_15 = _T_11058 | _T_6345; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11074 = _T_10815 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_0 = _T_11074 | _T_6354; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11090 = _T_10831 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_1 = _T_11090 | _T_6363; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11106 = _T_10847 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_2 = _T_11106 | _T_6372; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11122 = _T_10863 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_3 = _T_11122 | _T_6381; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11138 = _T_10879 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_4 = _T_11138 | _T_6390; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11154 = _T_10895 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_5 = _T_11154 | _T_6399; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11170 = _T_10911 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_6 = _T_11170 | _T_6408; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11186 = _T_10927 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_7 = _T_11186 | _T_6417; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11202 = _T_10943 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_8 = _T_11202 | _T_6426; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11218 = _T_10959 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_9 = _T_11218 | _T_6435; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11234 = _T_10975 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_10 = _T_11234 | _T_6444; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11250 = _T_10991 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_11 = _T_11250 | _T_6453; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11266 = _T_11007 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_12 = _T_11266 | _T_6462; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11282 = _T_11023 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_13 = _T_11282 | _T_6471; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11298 = _T_11039 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_14 = _T_11298 | _T_6480; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11314 = _T_11055 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_1_15 = _T_11314 | _T_6489; // @[el2_ifu_bp_ctl.scala 379:204]
  wire [1:0] _GEN_1488 = {{1'd0}, bht_wr_addr0[4]}; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_11329 = _GEN_1488 == 2'h2; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_11330 = _T_10815 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_0 = _T_11330 | _T_6498; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11346 = _T_10831 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_1 = _T_11346 | _T_6507; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11362 = _T_10847 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_2 = _T_11362 | _T_6516; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11378 = _T_10863 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_3 = _T_11378 | _T_6525; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11394 = _T_10879 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_4 = _T_11394 | _T_6534; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11410 = _T_10895 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_5 = _T_11410 | _T_6543; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11426 = _T_10911 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_6 = _T_11426 | _T_6552; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11442 = _T_10927 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_7 = _T_11442 | _T_6561; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11458 = _T_10943 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_8 = _T_11458 | _T_6570; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11474 = _T_10959 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_9 = _T_11474 | _T_6579; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11490 = _T_10975 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_10 = _T_11490 | _T_6588; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11506 = _T_10991 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_11 = _T_11506 | _T_6597; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11522 = _T_11007 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_12 = _T_11522 | _T_6606; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11538 = _T_11023 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_13 = _T_11538 | _T_6615; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11554 = _T_11039 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_14 = _T_11554 | _T_6624; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11570 = _T_11055 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_2_15 = _T_11570 | _T_6633; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11585 = _GEN_1488 == 2'h3; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_11586 = _T_10815 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_0 = _T_11586 | _T_6642; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11602 = _T_10831 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_1 = _T_11602 | _T_6651; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11618 = _T_10847 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_2 = _T_11618 | _T_6660; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11634 = _T_10863 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_3 = _T_11634 | _T_6669; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11650 = _T_10879 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_4 = _T_11650 | _T_6678; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11666 = _T_10895 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_5 = _T_11666 | _T_6687; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11682 = _T_10911 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_6 = _T_11682 | _T_6696; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11698 = _T_10927 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_7 = _T_11698 | _T_6705; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11714 = _T_10943 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_8 = _T_11714 | _T_6714; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11730 = _T_10959 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_9 = _T_11730 | _T_6723; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11746 = _T_10975 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_10 = _T_11746 | _T_6732; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11762 = _T_10991 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_11 = _T_11762 | _T_6741; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11778 = _T_11007 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_12 = _T_11778 | _T_6750; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11794 = _T_11023 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_13 = _T_11794 | _T_6759; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11810 = _T_11039 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_14 = _T_11810 | _T_6768; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11826 = _T_11055 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_3_15 = _T_11826 | _T_6777; // @[el2_ifu_bp_ctl.scala 379:204]
  wire [2:0] _GEN_1552 = {{2'd0}, bht_wr_addr0[4]}; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_11841 = _GEN_1552 == 3'h4; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_11842 = _T_10815 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_0 = _T_11842 | _T_6786; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11858 = _T_10831 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_1 = _T_11858 | _T_6795; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11874 = _T_10847 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_2 = _T_11874 | _T_6804; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11890 = _T_10863 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_3 = _T_11890 | _T_6813; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11906 = _T_10879 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_4 = _T_11906 | _T_6822; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11922 = _T_10895 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_5 = _T_11922 | _T_6831; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11938 = _T_10911 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_6 = _T_11938 | _T_6840; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11954 = _T_10927 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_7 = _T_11954 | _T_6849; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11970 = _T_10943 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_8 = _T_11970 | _T_6858; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_11986 = _T_10959 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_9 = _T_11986 | _T_6867; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12002 = _T_10975 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_10 = _T_12002 | _T_6876; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12018 = _T_10991 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_11 = _T_12018 | _T_6885; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12034 = _T_11007 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_12 = _T_12034 | _T_6894; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12050 = _T_11023 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_13 = _T_12050 | _T_6903; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12066 = _T_11039 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_14 = _T_12066 | _T_6912; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12082 = _T_11055 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_4_15 = _T_12082 | _T_6921; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12097 = _GEN_1552 == 3'h5; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_12098 = _T_10815 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_0 = _T_12098 | _T_6930; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12114 = _T_10831 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_1 = _T_12114 | _T_6939; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12130 = _T_10847 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_2 = _T_12130 | _T_6948; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12146 = _T_10863 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_3 = _T_12146 | _T_6957; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12162 = _T_10879 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_4 = _T_12162 | _T_6966; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12178 = _T_10895 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_5 = _T_12178 | _T_6975; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12194 = _T_10911 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_6 = _T_12194 | _T_6984; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12210 = _T_10927 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_7 = _T_12210 | _T_6993; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12226 = _T_10943 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_8 = _T_12226 | _T_7002; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12242 = _T_10959 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_9 = _T_12242 | _T_7011; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12258 = _T_10975 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_10 = _T_12258 | _T_7020; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12274 = _T_10991 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_11 = _T_12274 | _T_7029; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12290 = _T_11007 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_12 = _T_12290 | _T_7038; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12306 = _T_11023 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_13 = _T_12306 | _T_7047; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12322 = _T_11039 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_14 = _T_12322 | _T_7056; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12338 = _T_11055 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_5_15 = _T_12338 | _T_7065; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12353 = _GEN_1552 == 3'h6; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_12354 = _T_10815 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_0 = _T_12354 | _T_7074; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12370 = _T_10831 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_1 = _T_12370 | _T_7083; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12386 = _T_10847 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_2 = _T_12386 | _T_7092; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12402 = _T_10863 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_3 = _T_12402 | _T_7101; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12418 = _T_10879 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_4 = _T_12418 | _T_7110; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12434 = _T_10895 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_5 = _T_12434 | _T_7119; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12450 = _T_10911 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_6 = _T_12450 | _T_7128; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12466 = _T_10927 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_7 = _T_12466 | _T_7137; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12482 = _T_10943 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_8 = _T_12482 | _T_7146; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12498 = _T_10959 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_9 = _T_12498 | _T_7155; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12514 = _T_10975 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_10 = _T_12514 | _T_7164; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12530 = _T_10991 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_11 = _T_12530 | _T_7173; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12546 = _T_11007 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_12 = _T_12546 | _T_7182; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12562 = _T_11023 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_13 = _T_12562 | _T_7191; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12578 = _T_11039 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_14 = _T_12578 | _T_7200; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12594 = _T_11055 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_6_15 = _T_12594 | _T_7209; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12609 = _GEN_1552 == 3'h7; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_12610 = _T_10815 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_0 = _T_12610 | _T_7218; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12626 = _T_10831 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_1 = _T_12626 | _T_7227; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12642 = _T_10847 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_2 = _T_12642 | _T_7236; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12658 = _T_10863 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_3 = _T_12658 | _T_7245; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12674 = _T_10879 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_4 = _T_12674 | _T_7254; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12690 = _T_10895 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_5 = _T_12690 | _T_7263; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12706 = _T_10911 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_6 = _T_12706 | _T_7272; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12722 = _T_10927 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_7 = _T_12722 | _T_7281; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12738 = _T_10943 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_8 = _T_12738 | _T_7290; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12754 = _T_10959 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_9 = _T_12754 | _T_7299; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12770 = _T_10975 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_10 = _T_12770 | _T_7308; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12786 = _T_10991 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_11 = _T_12786 | _T_7317; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12802 = _T_11007 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_12 = _T_12802 | _T_7326; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12818 = _T_11023 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_13 = _T_12818 | _T_7335; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12834 = _T_11039 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_14 = _T_12834 | _T_7344; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12850 = _T_11055 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_7_15 = _T_12850 | _T_7353; // @[el2_ifu_bp_ctl.scala 379:204]
  wire [3:0] _GEN_1680 = {{3'd0}, bht_wr_addr0[4]}; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_12865 = _GEN_1680 == 4'h8; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_12866 = _T_10815 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_0 = _T_12866 | _T_7362; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12882 = _T_10831 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_1 = _T_12882 | _T_7371; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12898 = _T_10847 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_2 = _T_12898 | _T_7380; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12914 = _T_10863 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_3 = _T_12914 | _T_7389; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12930 = _T_10879 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_4 = _T_12930 | _T_7398; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12946 = _T_10895 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_5 = _T_12946 | _T_7407; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12962 = _T_10911 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_6 = _T_12962 | _T_7416; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12978 = _T_10927 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_7 = _T_12978 | _T_7425; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_12994 = _T_10943 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_8 = _T_12994 | _T_7434; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13010 = _T_10959 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_9 = _T_13010 | _T_7443; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13026 = _T_10975 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_10 = _T_13026 | _T_7452; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13042 = _T_10991 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_11 = _T_13042 | _T_7461; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13058 = _T_11007 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_12 = _T_13058 | _T_7470; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13074 = _T_11023 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_13 = _T_13074 | _T_7479; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13090 = _T_11039 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_14 = _T_13090 | _T_7488; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13106 = _T_11055 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_8_15 = _T_13106 | _T_7497; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13121 = _GEN_1680 == 4'h9; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_13122 = _T_10815 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_0 = _T_13122 | _T_7506; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13138 = _T_10831 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_1 = _T_13138 | _T_7515; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13154 = _T_10847 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_2 = _T_13154 | _T_7524; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13170 = _T_10863 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_3 = _T_13170 | _T_7533; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13186 = _T_10879 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_4 = _T_13186 | _T_7542; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13202 = _T_10895 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_5 = _T_13202 | _T_7551; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13218 = _T_10911 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_6 = _T_13218 | _T_7560; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13234 = _T_10927 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_7 = _T_13234 | _T_7569; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13250 = _T_10943 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_8 = _T_13250 | _T_7578; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13266 = _T_10959 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_9 = _T_13266 | _T_7587; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13282 = _T_10975 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_10 = _T_13282 | _T_7596; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13298 = _T_10991 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_11 = _T_13298 | _T_7605; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13314 = _T_11007 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_12 = _T_13314 | _T_7614; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13330 = _T_11023 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_13 = _T_13330 | _T_7623; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13346 = _T_11039 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_14 = _T_13346 | _T_7632; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13362 = _T_11055 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_9_15 = _T_13362 | _T_7641; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13377 = _GEN_1680 == 4'ha; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_13378 = _T_10815 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_0 = _T_13378 | _T_7650; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13394 = _T_10831 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_1 = _T_13394 | _T_7659; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13410 = _T_10847 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_2 = _T_13410 | _T_7668; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13426 = _T_10863 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_3 = _T_13426 | _T_7677; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13442 = _T_10879 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_4 = _T_13442 | _T_7686; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13458 = _T_10895 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_5 = _T_13458 | _T_7695; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13474 = _T_10911 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_6 = _T_13474 | _T_7704; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13490 = _T_10927 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_7 = _T_13490 | _T_7713; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13506 = _T_10943 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_8 = _T_13506 | _T_7722; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13522 = _T_10959 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_9 = _T_13522 | _T_7731; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13538 = _T_10975 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_10 = _T_13538 | _T_7740; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13554 = _T_10991 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_11 = _T_13554 | _T_7749; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13570 = _T_11007 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_12 = _T_13570 | _T_7758; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13586 = _T_11023 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_13 = _T_13586 | _T_7767; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13602 = _T_11039 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_14 = _T_13602 | _T_7776; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13618 = _T_11055 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_10_15 = _T_13618 | _T_7785; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13633 = _GEN_1680 == 4'hb; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_13634 = _T_10815 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_0 = _T_13634 | _T_7794; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13650 = _T_10831 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_1 = _T_13650 | _T_7803; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13666 = _T_10847 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_2 = _T_13666 | _T_7812; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13682 = _T_10863 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_3 = _T_13682 | _T_7821; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13698 = _T_10879 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_4 = _T_13698 | _T_7830; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13714 = _T_10895 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_5 = _T_13714 | _T_7839; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13730 = _T_10911 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_6 = _T_13730 | _T_7848; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13746 = _T_10927 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_7 = _T_13746 | _T_7857; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13762 = _T_10943 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_8 = _T_13762 | _T_7866; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13778 = _T_10959 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_9 = _T_13778 | _T_7875; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13794 = _T_10975 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_10 = _T_13794 | _T_7884; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13810 = _T_10991 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_11 = _T_13810 | _T_7893; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13826 = _T_11007 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_12 = _T_13826 | _T_7902; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13842 = _T_11023 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_13 = _T_13842 | _T_7911; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13858 = _T_11039 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_14 = _T_13858 | _T_7920; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13874 = _T_11055 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_11_15 = _T_13874 | _T_7929; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13889 = _GEN_1680 == 4'hc; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_13890 = _T_10815 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_0 = _T_13890 | _T_7938; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13906 = _T_10831 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_1 = _T_13906 | _T_7947; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13922 = _T_10847 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_2 = _T_13922 | _T_7956; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13938 = _T_10863 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_3 = _T_13938 | _T_7965; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13954 = _T_10879 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_4 = _T_13954 | _T_7974; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13970 = _T_10895 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_5 = _T_13970 | _T_7983; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_13986 = _T_10911 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_6 = _T_13986 | _T_7992; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14002 = _T_10927 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_7 = _T_14002 | _T_8001; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14018 = _T_10943 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_8 = _T_14018 | _T_8010; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14034 = _T_10959 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_9 = _T_14034 | _T_8019; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14050 = _T_10975 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_10 = _T_14050 | _T_8028; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14066 = _T_10991 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_11 = _T_14066 | _T_8037; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14082 = _T_11007 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_12 = _T_14082 | _T_8046; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14098 = _T_11023 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_13 = _T_14098 | _T_8055; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14114 = _T_11039 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_14 = _T_14114 | _T_8064; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14130 = _T_11055 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_12_15 = _T_14130 | _T_8073; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14145 = _GEN_1680 == 4'hd; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_14146 = _T_10815 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_0 = _T_14146 | _T_8082; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14162 = _T_10831 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_1 = _T_14162 | _T_8091; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14178 = _T_10847 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_2 = _T_14178 | _T_8100; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14194 = _T_10863 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_3 = _T_14194 | _T_8109; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14210 = _T_10879 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_4 = _T_14210 | _T_8118; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14226 = _T_10895 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_5 = _T_14226 | _T_8127; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14242 = _T_10911 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_6 = _T_14242 | _T_8136; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14258 = _T_10927 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_7 = _T_14258 | _T_8145; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14274 = _T_10943 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_8 = _T_14274 | _T_8154; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14290 = _T_10959 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_9 = _T_14290 | _T_8163; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14306 = _T_10975 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_10 = _T_14306 | _T_8172; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14322 = _T_10991 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_11 = _T_14322 | _T_8181; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14338 = _T_11007 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_12 = _T_14338 | _T_8190; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14354 = _T_11023 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_13 = _T_14354 | _T_8199; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14370 = _T_11039 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_14 = _T_14370 | _T_8208; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14386 = _T_11055 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_13_15 = _T_14386 | _T_8217; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14401 = _GEN_1680 == 4'he; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_14402 = _T_10815 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_0 = _T_14402 | _T_8226; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14418 = _T_10831 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_1 = _T_14418 | _T_8235; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14434 = _T_10847 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_2 = _T_14434 | _T_8244; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14450 = _T_10863 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_3 = _T_14450 | _T_8253; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14466 = _T_10879 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_4 = _T_14466 | _T_8262; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14482 = _T_10895 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_5 = _T_14482 | _T_8271; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14498 = _T_10911 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_6 = _T_14498 | _T_8280; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14514 = _T_10927 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_7 = _T_14514 | _T_8289; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14530 = _T_10943 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_8 = _T_14530 | _T_8298; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14546 = _T_10959 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_9 = _T_14546 | _T_8307; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14562 = _T_10975 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_10 = _T_14562 | _T_8316; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14578 = _T_10991 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_11 = _T_14578 | _T_8325; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14594 = _T_11007 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_12 = _T_14594 | _T_8334; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14610 = _T_11023 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_13 = _T_14610 | _T_8343; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14626 = _T_11039 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_14 = _T_14626 | _T_8352; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14642 = _T_11055 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_14_15 = _T_14642 | _T_8361; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14657 = _GEN_1680 == 4'hf; // @[el2_ifu_bp_ctl.scala 379:169]
  wire  _T_14658 = _T_10815 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_0 = _T_14658 | _T_8370; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14674 = _T_10831 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_1 = _T_14674 | _T_8379; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14690 = _T_10847 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_2 = _T_14690 | _T_8388; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14706 = _T_10863 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_3 = _T_14706 | _T_8397; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14722 = _T_10879 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_4 = _T_14722 | _T_8406; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14738 = _T_10895 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_5 = _T_14738 | _T_8415; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14754 = _T_10911 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_6 = _T_14754 | _T_8424; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14770 = _T_10927 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_7 = _T_14770 | _T_8433; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14786 = _T_10943 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_8 = _T_14786 | _T_8442; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14802 = _T_10959 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_9 = _T_14802 | _T_8451; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14818 = _T_10975 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_10 = _T_14818 | _T_8460; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14834 = _T_10991 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_11 = _T_14834 | _T_8469; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14850 = _T_11007 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_12 = _T_14850 | _T_8478; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14866 = _T_11023 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_13 = _T_14866 | _T_8487; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14882 = _T_11039 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_14 = _T_14882 | _T_8496; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14898 = _T_11055 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_0_15_15 = _T_14898 | _T_8505; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14911 = bht_wr_en0[1] & _T_10814; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_14914 = _T_14911 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_0 = _T_14914 | _T_8514; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14927 = bht_wr_en0[1] & _T_10830; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_14930 = _T_14927 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_1 = _T_14930 | _T_8523; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14943 = bht_wr_en0[1] & _T_10846; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_14946 = _T_14943 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_2 = _T_14946 | _T_8532; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14959 = bht_wr_en0[1] & _T_10862; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_14962 = _T_14959 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_3 = _T_14962 | _T_8541; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14975 = bht_wr_en0[1] & _T_10878; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_14978 = _T_14975 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_4 = _T_14978 | _T_8550; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_14991 = bht_wr_en0[1] & _T_10894; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_14994 = _T_14991 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_5 = _T_14994 | _T_8559; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15007 = bht_wr_en0[1] & _T_10910; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15010 = _T_15007 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_6 = _T_15010 | _T_8568; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15023 = bht_wr_en0[1] & _T_10926; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15026 = _T_15023 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_7 = _T_15026 | _T_8577; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15039 = bht_wr_en0[1] & _T_10942; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15042 = _T_15039 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_8 = _T_15042 | _T_8586; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15055 = bht_wr_en0[1] & _T_10958; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15058 = _T_15055 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_9 = _T_15058 | _T_8595; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15071 = bht_wr_en0[1] & _T_10974; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15074 = _T_15071 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_10 = _T_15074 | _T_8604; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15087 = bht_wr_en0[1] & _T_10990; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15090 = _T_15087 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_11 = _T_15090 | _T_8613; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15103 = bht_wr_en0[1] & _T_11006; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15106 = _T_15103 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_12 = _T_15106 | _T_8622; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15119 = bht_wr_en0[1] & _T_11022; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15122 = _T_15119 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_13 = _T_15122 | _T_8631; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15135 = bht_wr_en0[1] & _T_11038; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15138 = _T_15135 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_14 = _T_15138 | _T_8640; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15151 = bht_wr_en0[1] & _T_11054; // @[el2_ifu_bp_ctl.scala 379:17]
  wire  _T_15154 = _T_15151 & _T_10817; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_0_15 = _T_15154 | _T_8649; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15170 = _T_14911 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_0 = _T_15170 | _T_8658; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15186 = _T_14927 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_1 = _T_15186 | _T_8667; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15202 = _T_14943 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_2 = _T_15202 | _T_8676; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15218 = _T_14959 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_3 = _T_15218 | _T_8685; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15234 = _T_14975 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_4 = _T_15234 | _T_8694; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15250 = _T_14991 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_5 = _T_15250 | _T_8703; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15266 = _T_15007 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_6 = _T_15266 | _T_8712; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15282 = _T_15023 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_7 = _T_15282 | _T_8721; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15298 = _T_15039 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_8 = _T_15298 | _T_8730; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15314 = _T_15055 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_9 = _T_15314 | _T_8739; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15330 = _T_15071 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_10 = _T_15330 | _T_8748; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15346 = _T_15087 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_11 = _T_15346 | _T_8757; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15362 = _T_15103 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_12 = _T_15362 | _T_8766; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15378 = _T_15119 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_13 = _T_15378 | _T_8775; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15394 = _T_15135 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_14 = _T_15394 | _T_8784; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15410 = _T_15151 & bht_wr_addr0[4]; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_1_15 = _T_15410 | _T_8793; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15426 = _T_14911 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_0 = _T_15426 | _T_8802; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15442 = _T_14927 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_1 = _T_15442 | _T_8811; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15458 = _T_14943 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_2 = _T_15458 | _T_8820; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15474 = _T_14959 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_3 = _T_15474 | _T_8829; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15490 = _T_14975 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_4 = _T_15490 | _T_8838; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15506 = _T_14991 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_5 = _T_15506 | _T_8847; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15522 = _T_15007 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_6 = _T_15522 | _T_8856; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15538 = _T_15023 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_7 = _T_15538 | _T_8865; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15554 = _T_15039 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_8 = _T_15554 | _T_8874; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15570 = _T_15055 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_9 = _T_15570 | _T_8883; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15586 = _T_15071 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_10 = _T_15586 | _T_8892; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15602 = _T_15087 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_11 = _T_15602 | _T_8901; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15618 = _T_15103 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_12 = _T_15618 | _T_8910; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15634 = _T_15119 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_13 = _T_15634 | _T_8919; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15650 = _T_15135 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_14 = _T_15650 | _T_8928; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15666 = _T_15151 & _T_11329; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_2_15 = _T_15666 | _T_8937; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15682 = _T_14911 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_0 = _T_15682 | _T_8946; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15698 = _T_14927 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_1 = _T_15698 | _T_8955; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15714 = _T_14943 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_2 = _T_15714 | _T_8964; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15730 = _T_14959 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_3 = _T_15730 | _T_8973; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15746 = _T_14975 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_4 = _T_15746 | _T_8982; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15762 = _T_14991 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_5 = _T_15762 | _T_8991; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15778 = _T_15007 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_6 = _T_15778 | _T_9000; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15794 = _T_15023 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_7 = _T_15794 | _T_9009; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15810 = _T_15039 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_8 = _T_15810 | _T_9018; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15826 = _T_15055 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_9 = _T_15826 | _T_9027; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15842 = _T_15071 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_10 = _T_15842 | _T_9036; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15858 = _T_15087 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_11 = _T_15858 | _T_9045; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15874 = _T_15103 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_12 = _T_15874 | _T_9054; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15890 = _T_15119 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_13 = _T_15890 | _T_9063; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15906 = _T_15135 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_14 = _T_15906 | _T_9072; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15922 = _T_15151 & _T_11585; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_3_15 = _T_15922 | _T_9081; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15938 = _T_14911 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_0 = _T_15938 | _T_9090; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15954 = _T_14927 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_1 = _T_15954 | _T_9099; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15970 = _T_14943 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_2 = _T_15970 | _T_9108; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_15986 = _T_14959 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_3 = _T_15986 | _T_9117; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16002 = _T_14975 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_4 = _T_16002 | _T_9126; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16018 = _T_14991 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_5 = _T_16018 | _T_9135; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16034 = _T_15007 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_6 = _T_16034 | _T_9144; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16050 = _T_15023 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_7 = _T_16050 | _T_9153; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16066 = _T_15039 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_8 = _T_16066 | _T_9162; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16082 = _T_15055 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_9 = _T_16082 | _T_9171; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16098 = _T_15071 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_10 = _T_16098 | _T_9180; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16114 = _T_15087 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_11 = _T_16114 | _T_9189; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16130 = _T_15103 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_12 = _T_16130 | _T_9198; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16146 = _T_15119 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_13 = _T_16146 | _T_9207; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16162 = _T_15135 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_14 = _T_16162 | _T_9216; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16178 = _T_15151 & _T_11841; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_4_15 = _T_16178 | _T_9225; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16194 = _T_14911 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_0 = _T_16194 | _T_9234; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16210 = _T_14927 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_1 = _T_16210 | _T_9243; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16226 = _T_14943 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_2 = _T_16226 | _T_9252; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16242 = _T_14959 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_3 = _T_16242 | _T_9261; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16258 = _T_14975 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_4 = _T_16258 | _T_9270; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16274 = _T_14991 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_5 = _T_16274 | _T_9279; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16290 = _T_15007 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_6 = _T_16290 | _T_9288; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16306 = _T_15023 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_7 = _T_16306 | _T_9297; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16322 = _T_15039 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_8 = _T_16322 | _T_9306; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16338 = _T_15055 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_9 = _T_16338 | _T_9315; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16354 = _T_15071 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_10 = _T_16354 | _T_9324; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16370 = _T_15087 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_11 = _T_16370 | _T_9333; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16386 = _T_15103 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_12 = _T_16386 | _T_9342; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16402 = _T_15119 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_13 = _T_16402 | _T_9351; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16418 = _T_15135 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_14 = _T_16418 | _T_9360; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16434 = _T_15151 & _T_12097; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_5_15 = _T_16434 | _T_9369; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16450 = _T_14911 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_0 = _T_16450 | _T_9378; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16466 = _T_14927 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_1 = _T_16466 | _T_9387; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16482 = _T_14943 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_2 = _T_16482 | _T_9396; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16498 = _T_14959 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_3 = _T_16498 | _T_9405; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16514 = _T_14975 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_4 = _T_16514 | _T_9414; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16530 = _T_14991 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_5 = _T_16530 | _T_9423; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16546 = _T_15007 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_6 = _T_16546 | _T_9432; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16562 = _T_15023 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_7 = _T_16562 | _T_9441; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16578 = _T_15039 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_8 = _T_16578 | _T_9450; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16594 = _T_15055 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_9 = _T_16594 | _T_9459; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16610 = _T_15071 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_10 = _T_16610 | _T_9468; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16626 = _T_15087 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_11 = _T_16626 | _T_9477; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16642 = _T_15103 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_12 = _T_16642 | _T_9486; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16658 = _T_15119 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_13 = _T_16658 | _T_9495; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16674 = _T_15135 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_14 = _T_16674 | _T_9504; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16690 = _T_15151 & _T_12353; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_6_15 = _T_16690 | _T_9513; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16706 = _T_14911 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_0 = _T_16706 | _T_9522; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16722 = _T_14927 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_1 = _T_16722 | _T_9531; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16738 = _T_14943 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_2 = _T_16738 | _T_9540; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16754 = _T_14959 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_3 = _T_16754 | _T_9549; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16770 = _T_14975 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_4 = _T_16770 | _T_9558; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16786 = _T_14991 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_5 = _T_16786 | _T_9567; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16802 = _T_15007 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_6 = _T_16802 | _T_9576; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16818 = _T_15023 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_7 = _T_16818 | _T_9585; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16834 = _T_15039 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_8 = _T_16834 | _T_9594; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16850 = _T_15055 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_9 = _T_16850 | _T_9603; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16866 = _T_15071 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_10 = _T_16866 | _T_9612; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16882 = _T_15087 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_11 = _T_16882 | _T_9621; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16898 = _T_15103 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_12 = _T_16898 | _T_9630; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16914 = _T_15119 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_13 = _T_16914 | _T_9639; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16930 = _T_15135 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_14 = _T_16930 | _T_9648; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16946 = _T_15151 & _T_12609; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_7_15 = _T_16946 | _T_9657; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16962 = _T_14911 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_0 = _T_16962 | _T_9666; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16978 = _T_14927 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_1 = _T_16978 | _T_9675; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_16994 = _T_14943 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_2 = _T_16994 | _T_9684; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17010 = _T_14959 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_3 = _T_17010 | _T_9693; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17026 = _T_14975 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_4 = _T_17026 | _T_9702; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17042 = _T_14991 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_5 = _T_17042 | _T_9711; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17058 = _T_15007 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_6 = _T_17058 | _T_9720; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17074 = _T_15023 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_7 = _T_17074 | _T_9729; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17090 = _T_15039 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_8 = _T_17090 | _T_9738; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17106 = _T_15055 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_9 = _T_17106 | _T_9747; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17122 = _T_15071 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_10 = _T_17122 | _T_9756; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17138 = _T_15087 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_11 = _T_17138 | _T_9765; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17154 = _T_15103 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_12 = _T_17154 | _T_9774; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17170 = _T_15119 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_13 = _T_17170 | _T_9783; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17186 = _T_15135 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_14 = _T_17186 | _T_9792; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17202 = _T_15151 & _T_12865; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_8_15 = _T_17202 | _T_9801; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17218 = _T_14911 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_0 = _T_17218 | _T_9810; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17234 = _T_14927 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_1 = _T_17234 | _T_9819; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17250 = _T_14943 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_2 = _T_17250 | _T_9828; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17266 = _T_14959 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_3 = _T_17266 | _T_9837; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17282 = _T_14975 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_4 = _T_17282 | _T_9846; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17298 = _T_14991 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_5 = _T_17298 | _T_9855; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17314 = _T_15007 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_6 = _T_17314 | _T_9864; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17330 = _T_15023 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_7 = _T_17330 | _T_9873; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17346 = _T_15039 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_8 = _T_17346 | _T_9882; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17362 = _T_15055 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_9 = _T_17362 | _T_9891; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17378 = _T_15071 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_10 = _T_17378 | _T_9900; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17394 = _T_15087 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_11 = _T_17394 | _T_9909; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17410 = _T_15103 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_12 = _T_17410 | _T_9918; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17426 = _T_15119 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_13 = _T_17426 | _T_9927; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17442 = _T_15135 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_14 = _T_17442 | _T_9936; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17458 = _T_15151 & _T_13121; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_9_15 = _T_17458 | _T_9945; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17474 = _T_14911 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_0 = _T_17474 | _T_9954; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17490 = _T_14927 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_1 = _T_17490 | _T_9963; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17506 = _T_14943 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_2 = _T_17506 | _T_9972; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17522 = _T_14959 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_3 = _T_17522 | _T_9981; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17538 = _T_14975 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_4 = _T_17538 | _T_9990; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17554 = _T_14991 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_5 = _T_17554 | _T_9999; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17570 = _T_15007 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_6 = _T_17570 | _T_10008; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17586 = _T_15023 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_7 = _T_17586 | _T_10017; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17602 = _T_15039 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_8 = _T_17602 | _T_10026; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17618 = _T_15055 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_9 = _T_17618 | _T_10035; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17634 = _T_15071 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_10 = _T_17634 | _T_10044; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17650 = _T_15087 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_11 = _T_17650 | _T_10053; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17666 = _T_15103 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_12 = _T_17666 | _T_10062; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17682 = _T_15119 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_13 = _T_17682 | _T_10071; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17698 = _T_15135 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_14 = _T_17698 | _T_10080; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17714 = _T_15151 & _T_13377; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_10_15 = _T_17714 | _T_10089; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17730 = _T_14911 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_0 = _T_17730 | _T_10098; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17746 = _T_14927 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_1 = _T_17746 | _T_10107; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17762 = _T_14943 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_2 = _T_17762 | _T_10116; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17778 = _T_14959 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_3 = _T_17778 | _T_10125; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17794 = _T_14975 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_4 = _T_17794 | _T_10134; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17810 = _T_14991 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_5 = _T_17810 | _T_10143; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17826 = _T_15007 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_6 = _T_17826 | _T_10152; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17842 = _T_15023 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_7 = _T_17842 | _T_10161; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17858 = _T_15039 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_8 = _T_17858 | _T_10170; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17874 = _T_15055 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_9 = _T_17874 | _T_10179; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17890 = _T_15071 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_10 = _T_17890 | _T_10188; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17906 = _T_15087 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_11 = _T_17906 | _T_10197; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17922 = _T_15103 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_12 = _T_17922 | _T_10206; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17938 = _T_15119 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_13 = _T_17938 | _T_10215; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17954 = _T_15135 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_14 = _T_17954 | _T_10224; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17970 = _T_15151 & _T_13633; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_11_15 = _T_17970 | _T_10233; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_17986 = _T_14911 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_0 = _T_17986 | _T_10242; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18002 = _T_14927 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_1 = _T_18002 | _T_10251; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18018 = _T_14943 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_2 = _T_18018 | _T_10260; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18034 = _T_14959 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_3 = _T_18034 | _T_10269; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18050 = _T_14975 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_4 = _T_18050 | _T_10278; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18066 = _T_14991 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_5 = _T_18066 | _T_10287; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18082 = _T_15007 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_6 = _T_18082 | _T_10296; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18098 = _T_15023 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_7 = _T_18098 | _T_10305; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18114 = _T_15039 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_8 = _T_18114 | _T_10314; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18130 = _T_15055 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_9 = _T_18130 | _T_10323; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18146 = _T_15071 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_10 = _T_18146 | _T_10332; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18162 = _T_15087 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_11 = _T_18162 | _T_10341; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18178 = _T_15103 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_12 = _T_18178 | _T_10350; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18194 = _T_15119 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_13 = _T_18194 | _T_10359; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18210 = _T_15135 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_14 = _T_18210 | _T_10368; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18226 = _T_15151 & _T_13889; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_12_15 = _T_18226 | _T_10377; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18242 = _T_14911 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_0 = _T_18242 | _T_10386; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18258 = _T_14927 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_1 = _T_18258 | _T_10395; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18274 = _T_14943 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_2 = _T_18274 | _T_10404; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18290 = _T_14959 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_3 = _T_18290 | _T_10413; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18306 = _T_14975 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_4 = _T_18306 | _T_10422; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18322 = _T_14991 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_5 = _T_18322 | _T_10431; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18338 = _T_15007 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_6 = _T_18338 | _T_10440; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18354 = _T_15023 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_7 = _T_18354 | _T_10449; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18370 = _T_15039 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_8 = _T_18370 | _T_10458; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18386 = _T_15055 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_9 = _T_18386 | _T_10467; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18402 = _T_15071 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_10 = _T_18402 | _T_10476; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18418 = _T_15087 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_11 = _T_18418 | _T_10485; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18434 = _T_15103 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_12 = _T_18434 | _T_10494; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18450 = _T_15119 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_13 = _T_18450 | _T_10503; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18466 = _T_15135 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_14 = _T_18466 | _T_10512; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18482 = _T_15151 & _T_14145; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_13_15 = _T_18482 | _T_10521; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18498 = _T_14911 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_0 = _T_18498 | _T_10530; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18514 = _T_14927 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_1 = _T_18514 | _T_10539; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18530 = _T_14943 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_2 = _T_18530 | _T_10548; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18546 = _T_14959 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_3 = _T_18546 | _T_10557; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18562 = _T_14975 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_4 = _T_18562 | _T_10566; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18578 = _T_14991 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_5 = _T_18578 | _T_10575; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18594 = _T_15007 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_6 = _T_18594 | _T_10584; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18610 = _T_15023 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_7 = _T_18610 | _T_10593; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18626 = _T_15039 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_8 = _T_18626 | _T_10602; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18642 = _T_15055 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_9 = _T_18642 | _T_10611; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18658 = _T_15071 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_10 = _T_18658 | _T_10620; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18674 = _T_15087 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_11 = _T_18674 | _T_10629; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18690 = _T_15103 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_12 = _T_18690 | _T_10638; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18706 = _T_15119 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_13 = _T_18706 | _T_10647; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18722 = _T_15135 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_14 = _T_18722 | _T_10656; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18738 = _T_15151 & _T_14401; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_14_15 = _T_18738 | _T_10665; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18754 = _T_14911 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_0 = _T_18754 | _T_10674; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18770 = _T_14927 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_1 = _T_18770 | _T_10683; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18786 = _T_14943 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_2 = _T_18786 | _T_10692; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18802 = _T_14959 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_3 = _T_18802 | _T_10701; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18818 = _T_14975 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_4 = _T_18818 | _T_10710; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18834 = _T_14991 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_5 = _T_18834 | _T_10719; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18850 = _T_15007 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_6 = _T_18850 | _T_10728; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18866 = _T_15023 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_7 = _T_18866 | _T_10737; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18882 = _T_15039 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_8 = _T_18882 | _T_10746; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18898 = _T_15055 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_9 = _T_18898 | _T_10755; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18914 = _T_15071 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_10 = _T_18914 | _T_10764; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18930 = _T_15087 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_11 = _T_18930 | _T_10773; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18946 = _T_15103 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_12 = _T_18946 | _T_10782; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18962 = _T_15119 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_13 = _T_18962 | _T_10791; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18978 = _T_15135 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_14 = _T_18978 | _T_10800; // @[el2_ifu_bp_ctl.scala 379:204]
  wire  _T_18994 = _T_15151 & _T_14657; // @[el2_ifu_bp_ctl.scala 379:82]
  wire  bht_bank_sel_1_15_15 = _T_18994 | _T_10809; // @[el2_ifu_bp_ctl.scala 379:204]
  assign io_ifu_bp_hit_taken_f = _T_236 & _T_237; // @[el2_ifu_bp_ctl.scala 234:25]
  assign io_ifu_bp_btb_target_f = _T_425 ? rets_out_0[31:1] : bp_btb_target_adder_f[31:1]; // @[el2_ifu_bp_ctl.scala 316:26]
  assign io_ifu_bp_inst_mask_f = _T_273 | _T_274; // @[el2_ifu_bp_ctl.scala 254:25]
  assign io_ifu_bp_fghr_f = fghr; // @[el2_ifu_bp_ctl.scala 286:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_212; // @[el2_ifu_bp_ctl.scala 288:19]
  assign io_ifu_bp_ret_f = {_T_293,_T_299}; // @[el2_ifu_bp_ctl.scala 294:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_278; // @[el2_ifu_bp_ctl.scala 289:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[el2_ifu_bp_ctl.scala 290:21]
  assign io_ifu_bp_pc4_f = {_T_284,_T_287}; // @[el2_ifu_bp_ctl.scala 291:19]
  assign io_ifu_bp_valid_f = bht_valid_f & _T_342; // @[el2_ifu_bp_ctl.scala 293:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[el2_ifu_bp_ctl.scala 306:23]
  assign io_test_hash = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[el2_ifu_bp_ctl.scala 101:16]
  assign io_test_hash_p1 = _T_11 ^ _T_8[24:17]; // @[el2_ifu_bp_ctl.scala 106:19]
  assign io_test = _T_160 & _T_162; // @[el2_ifu_bp_ctl.scala 192:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_0 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_1 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_2 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_3 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_4 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_5 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_6 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_7 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_8 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_9 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_10 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_11 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_12 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_13 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_14 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_15 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_16 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_17 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_18 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_19 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_20 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_21 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_22 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_23 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_24 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_25 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_26 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_27 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_28 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_29 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_30 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_31 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_32 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_33 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_34 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_35 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_36 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_37 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_38 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_39 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_40 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_41 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_42 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_43 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_44 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_45 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_46 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_47 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_48 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_49 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_50 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_51 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_52 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_53 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_54 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_55 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_56 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_57 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_58 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_59 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_60 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_61 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_62 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_63 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_64 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_65 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_66 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_67 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_68 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_69 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_70 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_71 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_72 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_73 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_74 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_75 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_76 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_77 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_78 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_79 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_80 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_81 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_82 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_83 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_84 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_85 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_86 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_87 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_88 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_89 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_90 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_91 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_92 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_93 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_94 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_95 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_96 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_97 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_98 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_99 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_100 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_101 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_102 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_103 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_104 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_105 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_106 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_107 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_108 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_109 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_110 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_111 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_112 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_113 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_114 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_115 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_116 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_117 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_118 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_119 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_120 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_121 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_122 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_123 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_124 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_125 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_126 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_127 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_128 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_129 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_130 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_131 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_132 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_133 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_134 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_135 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_136 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_137 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_138 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_139 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_140 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_141 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_142 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_143 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_144 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_145 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_146 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_147 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_148 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_149 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_150 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_151 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_152 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_153 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_154 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_155 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_156 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_157 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_158 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_159 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_160 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_161 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_162 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_163 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_164 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_165 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_166 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_167 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_168 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_169 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_170 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_171 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_172 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_173 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_174 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_175 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_176 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_177 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_178 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_179 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_180 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_181 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_182 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_183 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_184 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_185 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_186 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_187 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_188 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_189 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_190 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_191 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_192 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_193 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_194 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_195 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_196 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_197 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_198 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_199 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_200 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_201 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_202 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_203 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_204 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_205 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_206 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_207 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_208 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_209 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_210 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_211 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_212 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_213 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_214 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_215 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_216 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_217 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_218 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_219 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_220 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_221 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_222 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_223 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_224 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_225 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_226 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_227 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_228 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_229 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_230 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_231 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_232 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_233 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_234 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_235 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_236 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_237 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_238 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_239 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_240 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_241 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_242 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_243 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_244 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_245 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_246 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_247 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_248 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_249 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_250 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_251 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_252 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_253 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_254 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_255 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  dec_tlu_way_wb_f = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_0 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_1 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_2 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_3 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_4 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_5 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_6 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_7 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_8 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_9 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_10 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_11 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_12 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_13 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_14 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_15 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_16 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_17 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_18 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_19 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_20 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_21 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_22 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_23 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_24 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_25 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_26 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_27 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_28 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_29 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_30 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_31 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_32 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_33 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_34 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_35 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_36 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_37 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_38 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_39 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_40 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_41 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_42 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_43 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_44 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_45 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_46 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_47 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_48 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_49 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_50 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_51 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_52 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_53 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_54 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_55 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_56 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_57 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_58 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_59 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_60 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_61 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_62 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_63 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_64 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_65 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_66 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_67 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_68 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_69 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_70 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_71 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_72 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_73 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_74 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_75 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_76 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_77 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_78 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_79 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_80 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_81 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_82 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_83 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_84 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_85 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_86 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_87 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_88 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_89 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_90 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_91 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_92 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_93 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_94 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_95 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_96 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_97 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_98 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_99 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_100 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_101 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_102 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_103 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_104 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_105 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_106 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_107 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_108 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_109 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_110 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_111 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_112 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_113 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_114 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_115 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_116 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_117 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_118 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_119 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_120 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_121 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_122 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_123 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_124 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_125 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_126 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_127 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_128 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_129 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_130 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_131 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_132 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_133 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_134 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_135 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_136 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_137 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_138 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_139 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_140 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_141 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_142 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_143 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_144 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_145 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_146 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_147 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_148 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_149 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_150 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_151 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_152 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_153 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_154 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_155 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_156 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_157 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_158 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_159 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_160 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_161 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_162 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_163 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_164 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_165 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_166 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_167 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_168 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_169 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_170 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_171 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_172 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_173 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_174 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_175 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_176 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_177 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_178 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_179 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_180 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_181 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_182 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_183 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_184 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_185 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_186 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_187 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_188 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_189 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_190 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_191 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_192 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_193 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_194 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_195 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_196 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_197 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_198 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_199 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_200 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_201 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_202 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_203 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_204 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_205 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_206 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_207 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_208 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_209 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_210 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_211 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_212 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_213 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_214 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_215 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_216 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_217 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_218 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_219 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_220 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_221 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_222 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_223 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_224 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_225 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_226 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_227 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_228 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_229 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_230 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_231 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_232 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_233 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_234 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_235 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_236 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_237 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_238 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_239 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_240 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_241 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_242 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_243 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_244 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_245 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_246 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_247 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_248 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_249 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_250 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_251 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_252 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_253 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_254 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_255 = _RAND_513[21:0];
  _RAND_514 = {1{`RANDOM}};
  fghr = _RAND_514[7:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1026[1:0];
  _RAND_1027 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1027[0:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1029[255:0];
  _RAND_1030 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1030[30:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_0 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_1 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_2 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_3 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_4 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_5 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_6 = _RAND_1037[31:0];
  _RAND_1038 = {1{`RANDOM}};
  rets_out_7 = _RAND_1038[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else begin
      leak_one_f_d1 <= leak_one_f;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_0 <= 22'h0;
    end else if (_T_573) begin
      btb_bank0_rd_data_way0_out_0 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_1 <= 22'h0;
    end else if (_T_576) begin
      btb_bank0_rd_data_way0_out_1 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_2 <= 22'h0;
    end else if (_T_579) begin
      btb_bank0_rd_data_way0_out_2 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_3 <= 22'h0;
    end else if (_T_582) begin
      btb_bank0_rd_data_way0_out_3 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_4 <= 22'h0;
    end else if (_T_585) begin
      btb_bank0_rd_data_way0_out_4 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_5 <= 22'h0;
    end else if (_T_588) begin
      btb_bank0_rd_data_way0_out_5 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_6 <= 22'h0;
    end else if (_T_591) begin
      btb_bank0_rd_data_way0_out_6 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_7 <= 22'h0;
    end else if (_T_594) begin
      btb_bank0_rd_data_way0_out_7 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_8 <= 22'h0;
    end else if (_T_597) begin
      btb_bank0_rd_data_way0_out_8 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_9 <= 22'h0;
    end else if (_T_600) begin
      btb_bank0_rd_data_way0_out_9 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_10 <= 22'h0;
    end else if (_T_603) begin
      btb_bank0_rd_data_way0_out_10 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_11 <= 22'h0;
    end else if (_T_606) begin
      btb_bank0_rd_data_way0_out_11 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_12 <= 22'h0;
    end else if (_T_609) begin
      btb_bank0_rd_data_way0_out_12 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_13 <= 22'h0;
    end else if (_T_612) begin
      btb_bank0_rd_data_way0_out_13 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_14 <= 22'h0;
    end else if (_T_615) begin
      btb_bank0_rd_data_way0_out_14 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_15 <= 22'h0;
    end else if (_T_618) begin
      btb_bank0_rd_data_way0_out_15 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_16 <= 22'h0;
    end else if (_T_621) begin
      btb_bank0_rd_data_way0_out_16 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_17 <= 22'h0;
    end else if (_T_624) begin
      btb_bank0_rd_data_way0_out_17 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_18 <= 22'h0;
    end else if (_T_627) begin
      btb_bank0_rd_data_way0_out_18 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_19 <= 22'h0;
    end else if (_T_630) begin
      btb_bank0_rd_data_way0_out_19 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_20 <= 22'h0;
    end else if (_T_633) begin
      btb_bank0_rd_data_way0_out_20 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_21 <= 22'h0;
    end else if (_T_636) begin
      btb_bank0_rd_data_way0_out_21 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_22 <= 22'h0;
    end else if (_T_639) begin
      btb_bank0_rd_data_way0_out_22 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_23 <= 22'h0;
    end else if (_T_642) begin
      btb_bank0_rd_data_way0_out_23 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_24 <= 22'h0;
    end else if (_T_645) begin
      btb_bank0_rd_data_way0_out_24 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_25 <= 22'h0;
    end else if (_T_648) begin
      btb_bank0_rd_data_way0_out_25 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_26 <= 22'h0;
    end else if (_T_651) begin
      btb_bank0_rd_data_way0_out_26 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_27 <= 22'h0;
    end else if (_T_654) begin
      btb_bank0_rd_data_way0_out_27 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_28 <= 22'h0;
    end else if (_T_657) begin
      btb_bank0_rd_data_way0_out_28 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_29 <= 22'h0;
    end else if (_T_660) begin
      btb_bank0_rd_data_way0_out_29 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_30 <= 22'h0;
    end else if (_T_663) begin
      btb_bank0_rd_data_way0_out_30 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_31 <= 22'h0;
    end else if (_T_666) begin
      btb_bank0_rd_data_way0_out_31 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_32 <= 22'h0;
    end else if (_T_669) begin
      btb_bank0_rd_data_way0_out_32 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_33 <= 22'h0;
    end else if (_T_672) begin
      btb_bank0_rd_data_way0_out_33 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_34 <= 22'h0;
    end else if (_T_675) begin
      btb_bank0_rd_data_way0_out_34 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_35 <= 22'h0;
    end else if (_T_678) begin
      btb_bank0_rd_data_way0_out_35 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_36 <= 22'h0;
    end else if (_T_681) begin
      btb_bank0_rd_data_way0_out_36 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_37 <= 22'h0;
    end else if (_T_684) begin
      btb_bank0_rd_data_way0_out_37 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_38 <= 22'h0;
    end else if (_T_687) begin
      btb_bank0_rd_data_way0_out_38 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_39 <= 22'h0;
    end else if (_T_690) begin
      btb_bank0_rd_data_way0_out_39 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_40 <= 22'h0;
    end else if (_T_693) begin
      btb_bank0_rd_data_way0_out_40 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_41 <= 22'h0;
    end else if (_T_696) begin
      btb_bank0_rd_data_way0_out_41 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_42 <= 22'h0;
    end else if (_T_699) begin
      btb_bank0_rd_data_way0_out_42 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_43 <= 22'h0;
    end else if (_T_702) begin
      btb_bank0_rd_data_way0_out_43 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_44 <= 22'h0;
    end else if (_T_705) begin
      btb_bank0_rd_data_way0_out_44 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_45 <= 22'h0;
    end else if (_T_708) begin
      btb_bank0_rd_data_way0_out_45 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_46 <= 22'h0;
    end else if (_T_711) begin
      btb_bank0_rd_data_way0_out_46 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_47 <= 22'h0;
    end else if (_T_714) begin
      btb_bank0_rd_data_way0_out_47 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_48 <= 22'h0;
    end else if (_T_717) begin
      btb_bank0_rd_data_way0_out_48 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_49 <= 22'h0;
    end else if (_T_720) begin
      btb_bank0_rd_data_way0_out_49 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_50 <= 22'h0;
    end else if (_T_723) begin
      btb_bank0_rd_data_way0_out_50 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_51 <= 22'h0;
    end else if (_T_726) begin
      btb_bank0_rd_data_way0_out_51 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_52 <= 22'h0;
    end else if (_T_729) begin
      btb_bank0_rd_data_way0_out_52 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_53 <= 22'h0;
    end else if (_T_732) begin
      btb_bank0_rd_data_way0_out_53 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_54 <= 22'h0;
    end else if (_T_735) begin
      btb_bank0_rd_data_way0_out_54 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_55 <= 22'h0;
    end else if (_T_738) begin
      btb_bank0_rd_data_way0_out_55 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_56 <= 22'h0;
    end else if (_T_741) begin
      btb_bank0_rd_data_way0_out_56 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_57 <= 22'h0;
    end else if (_T_744) begin
      btb_bank0_rd_data_way0_out_57 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_58 <= 22'h0;
    end else if (_T_747) begin
      btb_bank0_rd_data_way0_out_58 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_59 <= 22'h0;
    end else if (_T_750) begin
      btb_bank0_rd_data_way0_out_59 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_60 <= 22'h0;
    end else if (_T_753) begin
      btb_bank0_rd_data_way0_out_60 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_61 <= 22'h0;
    end else if (_T_756) begin
      btb_bank0_rd_data_way0_out_61 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_62 <= 22'h0;
    end else if (_T_759) begin
      btb_bank0_rd_data_way0_out_62 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_63 <= 22'h0;
    end else if (_T_762) begin
      btb_bank0_rd_data_way0_out_63 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_64 <= 22'h0;
    end else if (_T_765) begin
      btb_bank0_rd_data_way0_out_64 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_65 <= 22'h0;
    end else if (_T_768) begin
      btb_bank0_rd_data_way0_out_65 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_66 <= 22'h0;
    end else if (_T_771) begin
      btb_bank0_rd_data_way0_out_66 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_67 <= 22'h0;
    end else if (_T_774) begin
      btb_bank0_rd_data_way0_out_67 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_68 <= 22'h0;
    end else if (_T_777) begin
      btb_bank0_rd_data_way0_out_68 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_69 <= 22'h0;
    end else if (_T_780) begin
      btb_bank0_rd_data_way0_out_69 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_70 <= 22'h0;
    end else if (_T_783) begin
      btb_bank0_rd_data_way0_out_70 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_71 <= 22'h0;
    end else if (_T_786) begin
      btb_bank0_rd_data_way0_out_71 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_72 <= 22'h0;
    end else if (_T_789) begin
      btb_bank0_rd_data_way0_out_72 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_73 <= 22'h0;
    end else if (_T_792) begin
      btb_bank0_rd_data_way0_out_73 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_74 <= 22'h0;
    end else if (_T_795) begin
      btb_bank0_rd_data_way0_out_74 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_75 <= 22'h0;
    end else if (_T_798) begin
      btb_bank0_rd_data_way0_out_75 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_76 <= 22'h0;
    end else if (_T_801) begin
      btb_bank0_rd_data_way0_out_76 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_77 <= 22'h0;
    end else if (_T_804) begin
      btb_bank0_rd_data_way0_out_77 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_78 <= 22'h0;
    end else if (_T_807) begin
      btb_bank0_rd_data_way0_out_78 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_79 <= 22'h0;
    end else if (_T_810) begin
      btb_bank0_rd_data_way0_out_79 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_80 <= 22'h0;
    end else if (_T_813) begin
      btb_bank0_rd_data_way0_out_80 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_81 <= 22'h0;
    end else if (_T_816) begin
      btb_bank0_rd_data_way0_out_81 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_82 <= 22'h0;
    end else if (_T_819) begin
      btb_bank0_rd_data_way0_out_82 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_83 <= 22'h0;
    end else if (_T_822) begin
      btb_bank0_rd_data_way0_out_83 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_84 <= 22'h0;
    end else if (_T_825) begin
      btb_bank0_rd_data_way0_out_84 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_85 <= 22'h0;
    end else if (_T_828) begin
      btb_bank0_rd_data_way0_out_85 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_86 <= 22'h0;
    end else if (_T_831) begin
      btb_bank0_rd_data_way0_out_86 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_87 <= 22'h0;
    end else if (_T_834) begin
      btb_bank0_rd_data_way0_out_87 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_88 <= 22'h0;
    end else if (_T_837) begin
      btb_bank0_rd_data_way0_out_88 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_89 <= 22'h0;
    end else if (_T_840) begin
      btb_bank0_rd_data_way0_out_89 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_90 <= 22'h0;
    end else if (_T_843) begin
      btb_bank0_rd_data_way0_out_90 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_91 <= 22'h0;
    end else if (_T_846) begin
      btb_bank0_rd_data_way0_out_91 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_92 <= 22'h0;
    end else if (_T_849) begin
      btb_bank0_rd_data_way0_out_92 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_93 <= 22'h0;
    end else if (_T_852) begin
      btb_bank0_rd_data_way0_out_93 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_94 <= 22'h0;
    end else if (_T_855) begin
      btb_bank0_rd_data_way0_out_94 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_95 <= 22'h0;
    end else if (_T_858) begin
      btb_bank0_rd_data_way0_out_95 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_96 <= 22'h0;
    end else if (_T_861) begin
      btb_bank0_rd_data_way0_out_96 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_97 <= 22'h0;
    end else if (_T_864) begin
      btb_bank0_rd_data_way0_out_97 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_98 <= 22'h0;
    end else if (_T_867) begin
      btb_bank0_rd_data_way0_out_98 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_99 <= 22'h0;
    end else if (_T_870) begin
      btb_bank0_rd_data_way0_out_99 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_100 <= 22'h0;
    end else if (_T_873) begin
      btb_bank0_rd_data_way0_out_100 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_101 <= 22'h0;
    end else if (_T_876) begin
      btb_bank0_rd_data_way0_out_101 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_102 <= 22'h0;
    end else if (_T_879) begin
      btb_bank0_rd_data_way0_out_102 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_103 <= 22'h0;
    end else if (_T_882) begin
      btb_bank0_rd_data_way0_out_103 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_104 <= 22'h0;
    end else if (_T_885) begin
      btb_bank0_rd_data_way0_out_104 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_105 <= 22'h0;
    end else if (_T_888) begin
      btb_bank0_rd_data_way0_out_105 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_106 <= 22'h0;
    end else if (_T_891) begin
      btb_bank0_rd_data_way0_out_106 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_107 <= 22'h0;
    end else if (_T_894) begin
      btb_bank0_rd_data_way0_out_107 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_108 <= 22'h0;
    end else if (_T_897) begin
      btb_bank0_rd_data_way0_out_108 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_109 <= 22'h0;
    end else if (_T_900) begin
      btb_bank0_rd_data_way0_out_109 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_110 <= 22'h0;
    end else if (_T_903) begin
      btb_bank0_rd_data_way0_out_110 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_111 <= 22'h0;
    end else if (_T_906) begin
      btb_bank0_rd_data_way0_out_111 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_112 <= 22'h0;
    end else if (_T_909) begin
      btb_bank0_rd_data_way0_out_112 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_113 <= 22'h0;
    end else if (_T_912) begin
      btb_bank0_rd_data_way0_out_113 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_114 <= 22'h0;
    end else if (_T_915) begin
      btb_bank0_rd_data_way0_out_114 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_115 <= 22'h0;
    end else if (_T_918) begin
      btb_bank0_rd_data_way0_out_115 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_116 <= 22'h0;
    end else if (_T_921) begin
      btb_bank0_rd_data_way0_out_116 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_117 <= 22'h0;
    end else if (_T_924) begin
      btb_bank0_rd_data_way0_out_117 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_118 <= 22'h0;
    end else if (_T_927) begin
      btb_bank0_rd_data_way0_out_118 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_119 <= 22'h0;
    end else if (_T_930) begin
      btb_bank0_rd_data_way0_out_119 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_120 <= 22'h0;
    end else if (_T_933) begin
      btb_bank0_rd_data_way0_out_120 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_121 <= 22'h0;
    end else if (_T_936) begin
      btb_bank0_rd_data_way0_out_121 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_122 <= 22'h0;
    end else if (_T_939) begin
      btb_bank0_rd_data_way0_out_122 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_123 <= 22'h0;
    end else if (_T_942) begin
      btb_bank0_rd_data_way0_out_123 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_124 <= 22'h0;
    end else if (_T_945) begin
      btb_bank0_rd_data_way0_out_124 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_125 <= 22'h0;
    end else if (_T_948) begin
      btb_bank0_rd_data_way0_out_125 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_126 <= 22'h0;
    end else if (_T_951) begin
      btb_bank0_rd_data_way0_out_126 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_127 <= 22'h0;
    end else if (_T_954) begin
      btb_bank0_rd_data_way0_out_127 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_128 <= 22'h0;
    end else if (_T_957) begin
      btb_bank0_rd_data_way0_out_128 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_129 <= 22'h0;
    end else if (_T_960) begin
      btb_bank0_rd_data_way0_out_129 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_130 <= 22'h0;
    end else if (_T_963) begin
      btb_bank0_rd_data_way0_out_130 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_131 <= 22'h0;
    end else if (_T_966) begin
      btb_bank0_rd_data_way0_out_131 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_132 <= 22'h0;
    end else if (_T_969) begin
      btb_bank0_rd_data_way0_out_132 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_133 <= 22'h0;
    end else if (_T_972) begin
      btb_bank0_rd_data_way0_out_133 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_134 <= 22'h0;
    end else if (_T_975) begin
      btb_bank0_rd_data_way0_out_134 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_135 <= 22'h0;
    end else if (_T_978) begin
      btb_bank0_rd_data_way0_out_135 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_136 <= 22'h0;
    end else if (_T_981) begin
      btb_bank0_rd_data_way0_out_136 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_137 <= 22'h0;
    end else if (_T_984) begin
      btb_bank0_rd_data_way0_out_137 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_138 <= 22'h0;
    end else if (_T_987) begin
      btb_bank0_rd_data_way0_out_138 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_139 <= 22'h0;
    end else if (_T_990) begin
      btb_bank0_rd_data_way0_out_139 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_140 <= 22'h0;
    end else if (_T_993) begin
      btb_bank0_rd_data_way0_out_140 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_141 <= 22'h0;
    end else if (_T_996) begin
      btb_bank0_rd_data_way0_out_141 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_142 <= 22'h0;
    end else if (_T_999) begin
      btb_bank0_rd_data_way0_out_142 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_143 <= 22'h0;
    end else if (_T_1002) begin
      btb_bank0_rd_data_way0_out_143 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_144 <= 22'h0;
    end else if (_T_1005) begin
      btb_bank0_rd_data_way0_out_144 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_145 <= 22'h0;
    end else if (_T_1008) begin
      btb_bank0_rd_data_way0_out_145 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_146 <= 22'h0;
    end else if (_T_1011) begin
      btb_bank0_rd_data_way0_out_146 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_147 <= 22'h0;
    end else if (_T_1014) begin
      btb_bank0_rd_data_way0_out_147 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_148 <= 22'h0;
    end else if (_T_1017) begin
      btb_bank0_rd_data_way0_out_148 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_149 <= 22'h0;
    end else if (_T_1020) begin
      btb_bank0_rd_data_way0_out_149 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_150 <= 22'h0;
    end else if (_T_1023) begin
      btb_bank0_rd_data_way0_out_150 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_151 <= 22'h0;
    end else if (_T_1026) begin
      btb_bank0_rd_data_way0_out_151 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_152 <= 22'h0;
    end else if (_T_1029) begin
      btb_bank0_rd_data_way0_out_152 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_153 <= 22'h0;
    end else if (_T_1032) begin
      btb_bank0_rd_data_way0_out_153 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_154 <= 22'h0;
    end else if (_T_1035) begin
      btb_bank0_rd_data_way0_out_154 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_155 <= 22'h0;
    end else if (_T_1038) begin
      btb_bank0_rd_data_way0_out_155 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_156 <= 22'h0;
    end else if (_T_1041) begin
      btb_bank0_rd_data_way0_out_156 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_157 <= 22'h0;
    end else if (_T_1044) begin
      btb_bank0_rd_data_way0_out_157 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_158 <= 22'h0;
    end else if (_T_1047) begin
      btb_bank0_rd_data_way0_out_158 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_159 <= 22'h0;
    end else if (_T_1050) begin
      btb_bank0_rd_data_way0_out_159 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_160 <= 22'h0;
    end else if (_T_1053) begin
      btb_bank0_rd_data_way0_out_160 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_161 <= 22'h0;
    end else if (_T_1056) begin
      btb_bank0_rd_data_way0_out_161 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_162 <= 22'h0;
    end else if (_T_1059) begin
      btb_bank0_rd_data_way0_out_162 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_163 <= 22'h0;
    end else if (_T_1062) begin
      btb_bank0_rd_data_way0_out_163 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_164 <= 22'h0;
    end else if (_T_1065) begin
      btb_bank0_rd_data_way0_out_164 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_165 <= 22'h0;
    end else if (_T_1068) begin
      btb_bank0_rd_data_way0_out_165 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_166 <= 22'h0;
    end else if (_T_1071) begin
      btb_bank0_rd_data_way0_out_166 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_167 <= 22'h0;
    end else if (_T_1074) begin
      btb_bank0_rd_data_way0_out_167 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_168 <= 22'h0;
    end else if (_T_1077) begin
      btb_bank0_rd_data_way0_out_168 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_169 <= 22'h0;
    end else if (_T_1080) begin
      btb_bank0_rd_data_way0_out_169 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_170 <= 22'h0;
    end else if (_T_1083) begin
      btb_bank0_rd_data_way0_out_170 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_171 <= 22'h0;
    end else if (_T_1086) begin
      btb_bank0_rd_data_way0_out_171 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_172 <= 22'h0;
    end else if (_T_1089) begin
      btb_bank0_rd_data_way0_out_172 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_173 <= 22'h0;
    end else if (_T_1092) begin
      btb_bank0_rd_data_way0_out_173 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_174 <= 22'h0;
    end else if (_T_1095) begin
      btb_bank0_rd_data_way0_out_174 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_175 <= 22'h0;
    end else if (_T_1098) begin
      btb_bank0_rd_data_way0_out_175 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_176 <= 22'h0;
    end else if (_T_1101) begin
      btb_bank0_rd_data_way0_out_176 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_177 <= 22'h0;
    end else if (_T_1104) begin
      btb_bank0_rd_data_way0_out_177 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_178 <= 22'h0;
    end else if (_T_1107) begin
      btb_bank0_rd_data_way0_out_178 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_179 <= 22'h0;
    end else if (_T_1110) begin
      btb_bank0_rd_data_way0_out_179 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_180 <= 22'h0;
    end else if (_T_1113) begin
      btb_bank0_rd_data_way0_out_180 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_181 <= 22'h0;
    end else if (_T_1116) begin
      btb_bank0_rd_data_way0_out_181 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_182 <= 22'h0;
    end else if (_T_1119) begin
      btb_bank0_rd_data_way0_out_182 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_183 <= 22'h0;
    end else if (_T_1122) begin
      btb_bank0_rd_data_way0_out_183 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_184 <= 22'h0;
    end else if (_T_1125) begin
      btb_bank0_rd_data_way0_out_184 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_185 <= 22'h0;
    end else if (_T_1128) begin
      btb_bank0_rd_data_way0_out_185 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_186 <= 22'h0;
    end else if (_T_1131) begin
      btb_bank0_rd_data_way0_out_186 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_187 <= 22'h0;
    end else if (_T_1134) begin
      btb_bank0_rd_data_way0_out_187 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_188 <= 22'h0;
    end else if (_T_1137) begin
      btb_bank0_rd_data_way0_out_188 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_189 <= 22'h0;
    end else if (_T_1140) begin
      btb_bank0_rd_data_way0_out_189 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_190 <= 22'h0;
    end else if (_T_1143) begin
      btb_bank0_rd_data_way0_out_190 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_191 <= 22'h0;
    end else if (_T_1146) begin
      btb_bank0_rd_data_way0_out_191 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_192 <= 22'h0;
    end else if (_T_1149) begin
      btb_bank0_rd_data_way0_out_192 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_193 <= 22'h0;
    end else if (_T_1152) begin
      btb_bank0_rd_data_way0_out_193 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_194 <= 22'h0;
    end else if (_T_1155) begin
      btb_bank0_rd_data_way0_out_194 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_195 <= 22'h0;
    end else if (_T_1158) begin
      btb_bank0_rd_data_way0_out_195 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_196 <= 22'h0;
    end else if (_T_1161) begin
      btb_bank0_rd_data_way0_out_196 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_197 <= 22'h0;
    end else if (_T_1164) begin
      btb_bank0_rd_data_way0_out_197 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_198 <= 22'h0;
    end else if (_T_1167) begin
      btb_bank0_rd_data_way0_out_198 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_199 <= 22'h0;
    end else if (_T_1170) begin
      btb_bank0_rd_data_way0_out_199 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_200 <= 22'h0;
    end else if (_T_1173) begin
      btb_bank0_rd_data_way0_out_200 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_201 <= 22'h0;
    end else if (_T_1176) begin
      btb_bank0_rd_data_way0_out_201 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_202 <= 22'h0;
    end else if (_T_1179) begin
      btb_bank0_rd_data_way0_out_202 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_203 <= 22'h0;
    end else if (_T_1182) begin
      btb_bank0_rd_data_way0_out_203 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_204 <= 22'h0;
    end else if (_T_1185) begin
      btb_bank0_rd_data_way0_out_204 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_205 <= 22'h0;
    end else if (_T_1188) begin
      btb_bank0_rd_data_way0_out_205 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_206 <= 22'h0;
    end else if (_T_1191) begin
      btb_bank0_rd_data_way0_out_206 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_207 <= 22'h0;
    end else if (_T_1194) begin
      btb_bank0_rd_data_way0_out_207 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_208 <= 22'h0;
    end else if (_T_1197) begin
      btb_bank0_rd_data_way0_out_208 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_209 <= 22'h0;
    end else if (_T_1200) begin
      btb_bank0_rd_data_way0_out_209 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_210 <= 22'h0;
    end else if (_T_1203) begin
      btb_bank0_rd_data_way0_out_210 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_211 <= 22'h0;
    end else if (_T_1206) begin
      btb_bank0_rd_data_way0_out_211 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_212 <= 22'h0;
    end else if (_T_1209) begin
      btb_bank0_rd_data_way0_out_212 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_213 <= 22'h0;
    end else if (_T_1212) begin
      btb_bank0_rd_data_way0_out_213 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_214 <= 22'h0;
    end else if (_T_1215) begin
      btb_bank0_rd_data_way0_out_214 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_215 <= 22'h0;
    end else if (_T_1218) begin
      btb_bank0_rd_data_way0_out_215 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_216 <= 22'h0;
    end else if (_T_1221) begin
      btb_bank0_rd_data_way0_out_216 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_217 <= 22'h0;
    end else if (_T_1224) begin
      btb_bank0_rd_data_way0_out_217 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_218 <= 22'h0;
    end else if (_T_1227) begin
      btb_bank0_rd_data_way0_out_218 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_219 <= 22'h0;
    end else if (_T_1230) begin
      btb_bank0_rd_data_way0_out_219 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_220 <= 22'h0;
    end else if (_T_1233) begin
      btb_bank0_rd_data_way0_out_220 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_221 <= 22'h0;
    end else if (_T_1236) begin
      btb_bank0_rd_data_way0_out_221 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_222 <= 22'h0;
    end else if (_T_1239) begin
      btb_bank0_rd_data_way0_out_222 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_223 <= 22'h0;
    end else if (_T_1242) begin
      btb_bank0_rd_data_way0_out_223 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_224 <= 22'h0;
    end else if (_T_1245) begin
      btb_bank0_rd_data_way0_out_224 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_225 <= 22'h0;
    end else if (_T_1248) begin
      btb_bank0_rd_data_way0_out_225 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_226 <= 22'h0;
    end else if (_T_1251) begin
      btb_bank0_rd_data_way0_out_226 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_227 <= 22'h0;
    end else if (_T_1254) begin
      btb_bank0_rd_data_way0_out_227 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_228 <= 22'h0;
    end else if (_T_1257) begin
      btb_bank0_rd_data_way0_out_228 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_229 <= 22'h0;
    end else if (_T_1260) begin
      btb_bank0_rd_data_way0_out_229 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_230 <= 22'h0;
    end else if (_T_1263) begin
      btb_bank0_rd_data_way0_out_230 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_231 <= 22'h0;
    end else if (_T_1266) begin
      btb_bank0_rd_data_way0_out_231 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_232 <= 22'h0;
    end else if (_T_1269) begin
      btb_bank0_rd_data_way0_out_232 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_233 <= 22'h0;
    end else if (_T_1272) begin
      btb_bank0_rd_data_way0_out_233 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_234 <= 22'h0;
    end else if (_T_1275) begin
      btb_bank0_rd_data_way0_out_234 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_235 <= 22'h0;
    end else if (_T_1278) begin
      btb_bank0_rd_data_way0_out_235 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_236 <= 22'h0;
    end else if (_T_1281) begin
      btb_bank0_rd_data_way0_out_236 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_237 <= 22'h0;
    end else if (_T_1284) begin
      btb_bank0_rd_data_way0_out_237 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_238 <= 22'h0;
    end else if (_T_1287) begin
      btb_bank0_rd_data_way0_out_238 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_239 <= 22'h0;
    end else if (_T_1290) begin
      btb_bank0_rd_data_way0_out_239 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_240 <= 22'h0;
    end else if (_T_1293) begin
      btb_bank0_rd_data_way0_out_240 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_241 <= 22'h0;
    end else if (_T_1296) begin
      btb_bank0_rd_data_way0_out_241 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_242 <= 22'h0;
    end else if (_T_1299) begin
      btb_bank0_rd_data_way0_out_242 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_243 <= 22'h0;
    end else if (_T_1302) begin
      btb_bank0_rd_data_way0_out_243 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_244 <= 22'h0;
    end else if (_T_1305) begin
      btb_bank0_rd_data_way0_out_244 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_245 <= 22'h0;
    end else if (_T_1308) begin
      btb_bank0_rd_data_way0_out_245 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_246 <= 22'h0;
    end else if (_T_1311) begin
      btb_bank0_rd_data_way0_out_246 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_247 <= 22'h0;
    end else if (_T_1314) begin
      btb_bank0_rd_data_way0_out_247 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_248 <= 22'h0;
    end else if (_T_1317) begin
      btb_bank0_rd_data_way0_out_248 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_249 <= 22'h0;
    end else if (_T_1320) begin
      btb_bank0_rd_data_way0_out_249 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_250 <= 22'h0;
    end else if (_T_1323) begin
      btb_bank0_rd_data_way0_out_250 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_251 <= 22'h0;
    end else if (_T_1326) begin
      btb_bank0_rd_data_way0_out_251 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_252 <= 22'h0;
    end else if (_T_1329) begin
      btb_bank0_rd_data_way0_out_252 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_253 <= 22'h0;
    end else if (_T_1332) begin
      btb_bank0_rd_data_way0_out_253 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_254 <= 22'h0;
    end else if (_T_1335) begin
      btb_bank0_rd_data_way0_out_254 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way0_out_255 <= 22'h0;
    end else if (_T_1338) begin
      btb_bank0_rd_data_way0_out_255 <= btb_wr_data;
    end
    if (reset) begin
      dec_tlu_way_wb_f <= 1'h0;
    end else begin
      dec_tlu_way_wb_f <= io_dec_tlu_br0_r_pkt_way;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_0 <= 22'h0;
    end else if (_T_1341) begin
      btb_bank0_rd_data_way1_out_0 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_1 <= 22'h0;
    end else if (_T_1344) begin
      btb_bank0_rd_data_way1_out_1 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_2 <= 22'h0;
    end else if (_T_1347) begin
      btb_bank0_rd_data_way1_out_2 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_3 <= 22'h0;
    end else if (_T_1350) begin
      btb_bank0_rd_data_way1_out_3 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_4 <= 22'h0;
    end else if (_T_1353) begin
      btb_bank0_rd_data_way1_out_4 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_5 <= 22'h0;
    end else if (_T_1356) begin
      btb_bank0_rd_data_way1_out_5 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_6 <= 22'h0;
    end else if (_T_1359) begin
      btb_bank0_rd_data_way1_out_6 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_7 <= 22'h0;
    end else if (_T_1362) begin
      btb_bank0_rd_data_way1_out_7 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_8 <= 22'h0;
    end else if (_T_1365) begin
      btb_bank0_rd_data_way1_out_8 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_9 <= 22'h0;
    end else if (_T_1368) begin
      btb_bank0_rd_data_way1_out_9 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_10 <= 22'h0;
    end else if (_T_1371) begin
      btb_bank0_rd_data_way1_out_10 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_11 <= 22'h0;
    end else if (_T_1374) begin
      btb_bank0_rd_data_way1_out_11 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_12 <= 22'h0;
    end else if (_T_1377) begin
      btb_bank0_rd_data_way1_out_12 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_13 <= 22'h0;
    end else if (_T_1380) begin
      btb_bank0_rd_data_way1_out_13 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_14 <= 22'h0;
    end else if (_T_1383) begin
      btb_bank0_rd_data_way1_out_14 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_15 <= 22'h0;
    end else if (_T_1386) begin
      btb_bank0_rd_data_way1_out_15 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_16 <= 22'h0;
    end else if (_T_1389) begin
      btb_bank0_rd_data_way1_out_16 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_17 <= 22'h0;
    end else if (_T_1392) begin
      btb_bank0_rd_data_way1_out_17 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_18 <= 22'h0;
    end else if (_T_1395) begin
      btb_bank0_rd_data_way1_out_18 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_19 <= 22'h0;
    end else if (_T_1398) begin
      btb_bank0_rd_data_way1_out_19 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_20 <= 22'h0;
    end else if (_T_1401) begin
      btb_bank0_rd_data_way1_out_20 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_21 <= 22'h0;
    end else if (_T_1404) begin
      btb_bank0_rd_data_way1_out_21 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_22 <= 22'h0;
    end else if (_T_1407) begin
      btb_bank0_rd_data_way1_out_22 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_23 <= 22'h0;
    end else if (_T_1410) begin
      btb_bank0_rd_data_way1_out_23 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_24 <= 22'h0;
    end else if (_T_1413) begin
      btb_bank0_rd_data_way1_out_24 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_25 <= 22'h0;
    end else if (_T_1416) begin
      btb_bank0_rd_data_way1_out_25 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_26 <= 22'h0;
    end else if (_T_1419) begin
      btb_bank0_rd_data_way1_out_26 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_27 <= 22'h0;
    end else if (_T_1422) begin
      btb_bank0_rd_data_way1_out_27 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_28 <= 22'h0;
    end else if (_T_1425) begin
      btb_bank0_rd_data_way1_out_28 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_29 <= 22'h0;
    end else if (_T_1428) begin
      btb_bank0_rd_data_way1_out_29 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_30 <= 22'h0;
    end else if (_T_1431) begin
      btb_bank0_rd_data_way1_out_30 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_31 <= 22'h0;
    end else if (_T_1434) begin
      btb_bank0_rd_data_way1_out_31 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_32 <= 22'h0;
    end else if (_T_1437) begin
      btb_bank0_rd_data_way1_out_32 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_33 <= 22'h0;
    end else if (_T_1440) begin
      btb_bank0_rd_data_way1_out_33 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_34 <= 22'h0;
    end else if (_T_1443) begin
      btb_bank0_rd_data_way1_out_34 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_35 <= 22'h0;
    end else if (_T_1446) begin
      btb_bank0_rd_data_way1_out_35 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_36 <= 22'h0;
    end else if (_T_1449) begin
      btb_bank0_rd_data_way1_out_36 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_37 <= 22'h0;
    end else if (_T_1452) begin
      btb_bank0_rd_data_way1_out_37 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_38 <= 22'h0;
    end else if (_T_1455) begin
      btb_bank0_rd_data_way1_out_38 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_39 <= 22'h0;
    end else if (_T_1458) begin
      btb_bank0_rd_data_way1_out_39 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_40 <= 22'h0;
    end else if (_T_1461) begin
      btb_bank0_rd_data_way1_out_40 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_41 <= 22'h0;
    end else if (_T_1464) begin
      btb_bank0_rd_data_way1_out_41 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_42 <= 22'h0;
    end else if (_T_1467) begin
      btb_bank0_rd_data_way1_out_42 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_43 <= 22'h0;
    end else if (_T_1470) begin
      btb_bank0_rd_data_way1_out_43 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_44 <= 22'h0;
    end else if (_T_1473) begin
      btb_bank0_rd_data_way1_out_44 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_45 <= 22'h0;
    end else if (_T_1476) begin
      btb_bank0_rd_data_way1_out_45 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_46 <= 22'h0;
    end else if (_T_1479) begin
      btb_bank0_rd_data_way1_out_46 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_47 <= 22'h0;
    end else if (_T_1482) begin
      btb_bank0_rd_data_way1_out_47 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_48 <= 22'h0;
    end else if (_T_1485) begin
      btb_bank0_rd_data_way1_out_48 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_49 <= 22'h0;
    end else if (_T_1488) begin
      btb_bank0_rd_data_way1_out_49 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_50 <= 22'h0;
    end else if (_T_1491) begin
      btb_bank0_rd_data_way1_out_50 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_51 <= 22'h0;
    end else if (_T_1494) begin
      btb_bank0_rd_data_way1_out_51 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_52 <= 22'h0;
    end else if (_T_1497) begin
      btb_bank0_rd_data_way1_out_52 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_53 <= 22'h0;
    end else if (_T_1500) begin
      btb_bank0_rd_data_way1_out_53 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_54 <= 22'h0;
    end else if (_T_1503) begin
      btb_bank0_rd_data_way1_out_54 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_55 <= 22'h0;
    end else if (_T_1506) begin
      btb_bank0_rd_data_way1_out_55 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_56 <= 22'h0;
    end else if (_T_1509) begin
      btb_bank0_rd_data_way1_out_56 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_57 <= 22'h0;
    end else if (_T_1512) begin
      btb_bank0_rd_data_way1_out_57 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_58 <= 22'h0;
    end else if (_T_1515) begin
      btb_bank0_rd_data_way1_out_58 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_59 <= 22'h0;
    end else if (_T_1518) begin
      btb_bank0_rd_data_way1_out_59 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_60 <= 22'h0;
    end else if (_T_1521) begin
      btb_bank0_rd_data_way1_out_60 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_61 <= 22'h0;
    end else if (_T_1524) begin
      btb_bank0_rd_data_way1_out_61 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_62 <= 22'h0;
    end else if (_T_1527) begin
      btb_bank0_rd_data_way1_out_62 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_63 <= 22'h0;
    end else if (_T_1530) begin
      btb_bank0_rd_data_way1_out_63 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_64 <= 22'h0;
    end else if (_T_1533) begin
      btb_bank0_rd_data_way1_out_64 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_65 <= 22'h0;
    end else if (_T_1536) begin
      btb_bank0_rd_data_way1_out_65 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_66 <= 22'h0;
    end else if (_T_1539) begin
      btb_bank0_rd_data_way1_out_66 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_67 <= 22'h0;
    end else if (_T_1542) begin
      btb_bank0_rd_data_way1_out_67 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_68 <= 22'h0;
    end else if (_T_1545) begin
      btb_bank0_rd_data_way1_out_68 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_69 <= 22'h0;
    end else if (_T_1548) begin
      btb_bank0_rd_data_way1_out_69 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_70 <= 22'h0;
    end else if (_T_1551) begin
      btb_bank0_rd_data_way1_out_70 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_71 <= 22'h0;
    end else if (_T_1554) begin
      btb_bank0_rd_data_way1_out_71 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_72 <= 22'h0;
    end else if (_T_1557) begin
      btb_bank0_rd_data_way1_out_72 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_73 <= 22'h0;
    end else if (_T_1560) begin
      btb_bank0_rd_data_way1_out_73 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_74 <= 22'h0;
    end else if (_T_1563) begin
      btb_bank0_rd_data_way1_out_74 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_75 <= 22'h0;
    end else if (_T_1566) begin
      btb_bank0_rd_data_way1_out_75 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_76 <= 22'h0;
    end else if (_T_1569) begin
      btb_bank0_rd_data_way1_out_76 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_77 <= 22'h0;
    end else if (_T_1572) begin
      btb_bank0_rd_data_way1_out_77 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_78 <= 22'h0;
    end else if (_T_1575) begin
      btb_bank0_rd_data_way1_out_78 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_79 <= 22'h0;
    end else if (_T_1578) begin
      btb_bank0_rd_data_way1_out_79 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_80 <= 22'h0;
    end else if (_T_1581) begin
      btb_bank0_rd_data_way1_out_80 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_81 <= 22'h0;
    end else if (_T_1584) begin
      btb_bank0_rd_data_way1_out_81 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_82 <= 22'h0;
    end else if (_T_1587) begin
      btb_bank0_rd_data_way1_out_82 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_83 <= 22'h0;
    end else if (_T_1590) begin
      btb_bank0_rd_data_way1_out_83 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_84 <= 22'h0;
    end else if (_T_1593) begin
      btb_bank0_rd_data_way1_out_84 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_85 <= 22'h0;
    end else if (_T_1596) begin
      btb_bank0_rd_data_way1_out_85 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_86 <= 22'h0;
    end else if (_T_1599) begin
      btb_bank0_rd_data_way1_out_86 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_87 <= 22'h0;
    end else if (_T_1602) begin
      btb_bank0_rd_data_way1_out_87 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_88 <= 22'h0;
    end else if (_T_1605) begin
      btb_bank0_rd_data_way1_out_88 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_89 <= 22'h0;
    end else if (_T_1608) begin
      btb_bank0_rd_data_way1_out_89 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_90 <= 22'h0;
    end else if (_T_1611) begin
      btb_bank0_rd_data_way1_out_90 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_91 <= 22'h0;
    end else if (_T_1614) begin
      btb_bank0_rd_data_way1_out_91 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_92 <= 22'h0;
    end else if (_T_1617) begin
      btb_bank0_rd_data_way1_out_92 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_93 <= 22'h0;
    end else if (_T_1620) begin
      btb_bank0_rd_data_way1_out_93 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_94 <= 22'h0;
    end else if (_T_1623) begin
      btb_bank0_rd_data_way1_out_94 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_95 <= 22'h0;
    end else if (_T_1626) begin
      btb_bank0_rd_data_way1_out_95 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_96 <= 22'h0;
    end else if (_T_1629) begin
      btb_bank0_rd_data_way1_out_96 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_97 <= 22'h0;
    end else if (_T_1632) begin
      btb_bank0_rd_data_way1_out_97 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_98 <= 22'h0;
    end else if (_T_1635) begin
      btb_bank0_rd_data_way1_out_98 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_99 <= 22'h0;
    end else if (_T_1638) begin
      btb_bank0_rd_data_way1_out_99 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_100 <= 22'h0;
    end else if (_T_1641) begin
      btb_bank0_rd_data_way1_out_100 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_101 <= 22'h0;
    end else if (_T_1644) begin
      btb_bank0_rd_data_way1_out_101 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_102 <= 22'h0;
    end else if (_T_1647) begin
      btb_bank0_rd_data_way1_out_102 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_103 <= 22'h0;
    end else if (_T_1650) begin
      btb_bank0_rd_data_way1_out_103 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_104 <= 22'h0;
    end else if (_T_1653) begin
      btb_bank0_rd_data_way1_out_104 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_105 <= 22'h0;
    end else if (_T_1656) begin
      btb_bank0_rd_data_way1_out_105 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_106 <= 22'h0;
    end else if (_T_1659) begin
      btb_bank0_rd_data_way1_out_106 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_107 <= 22'h0;
    end else if (_T_1662) begin
      btb_bank0_rd_data_way1_out_107 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_108 <= 22'h0;
    end else if (_T_1665) begin
      btb_bank0_rd_data_way1_out_108 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_109 <= 22'h0;
    end else if (_T_1668) begin
      btb_bank0_rd_data_way1_out_109 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_110 <= 22'h0;
    end else if (_T_1671) begin
      btb_bank0_rd_data_way1_out_110 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_111 <= 22'h0;
    end else if (_T_1674) begin
      btb_bank0_rd_data_way1_out_111 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_112 <= 22'h0;
    end else if (_T_1677) begin
      btb_bank0_rd_data_way1_out_112 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_113 <= 22'h0;
    end else if (_T_1680) begin
      btb_bank0_rd_data_way1_out_113 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_114 <= 22'h0;
    end else if (_T_1683) begin
      btb_bank0_rd_data_way1_out_114 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_115 <= 22'h0;
    end else if (_T_1686) begin
      btb_bank0_rd_data_way1_out_115 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_116 <= 22'h0;
    end else if (_T_1689) begin
      btb_bank0_rd_data_way1_out_116 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_117 <= 22'h0;
    end else if (_T_1692) begin
      btb_bank0_rd_data_way1_out_117 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_118 <= 22'h0;
    end else if (_T_1695) begin
      btb_bank0_rd_data_way1_out_118 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_119 <= 22'h0;
    end else if (_T_1698) begin
      btb_bank0_rd_data_way1_out_119 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_120 <= 22'h0;
    end else if (_T_1701) begin
      btb_bank0_rd_data_way1_out_120 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_121 <= 22'h0;
    end else if (_T_1704) begin
      btb_bank0_rd_data_way1_out_121 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_122 <= 22'h0;
    end else if (_T_1707) begin
      btb_bank0_rd_data_way1_out_122 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_123 <= 22'h0;
    end else if (_T_1710) begin
      btb_bank0_rd_data_way1_out_123 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_124 <= 22'h0;
    end else if (_T_1713) begin
      btb_bank0_rd_data_way1_out_124 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_125 <= 22'h0;
    end else if (_T_1716) begin
      btb_bank0_rd_data_way1_out_125 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_126 <= 22'h0;
    end else if (_T_1719) begin
      btb_bank0_rd_data_way1_out_126 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_127 <= 22'h0;
    end else if (_T_1722) begin
      btb_bank0_rd_data_way1_out_127 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_128 <= 22'h0;
    end else if (_T_1725) begin
      btb_bank0_rd_data_way1_out_128 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_129 <= 22'h0;
    end else if (_T_1728) begin
      btb_bank0_rd_data_way1_out_129 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_130 <= 22'h0;
    end else if (_T_1731) begin
      btb_bank0_rd_data_way1_out_130 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_131 <= 22'h0;
    end else if (_T_1734) begin
      btb_bank0_rd_data_way1_out_131 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_132 <= 22'h0;
    end else if (_T_1737) begin
      btb_bank0_rd_data_way1_out_132 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_133 <= 22'h0;
    end else if (_T_1740) begin
      btb_bank0_rd_data_way1_out_133 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_134 <= 22'h0;
    end else if (_T_1743) begin
      btb_bank0_rd_data_way1_out_134 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_135 <= 22'h0;
    end else if (_T_1746) begin
      btb_bank0_rd_data_way1_out_135 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_136 <= 22'h0;
    end else if (_T_1749) begin
      btb_bank0_rd_data_way1_out_136 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_137 <= 22'h0;
    end else if (_T_1752) begin
      btb_bank0_rd_data_way1_out_137 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_138 <= 22'h0;
    end else if (_T_1755) begin
      btb_bank0_rd_data_way1_out_138 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_139 <= 22'h0;
    end else if (_T_1758) begin
      btb_bank0_rd_data_way1_out_139 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_140 <= 22'h0;
    end else if (_T_1761) begin
      btb_bank0_rd_data_way1_out_140 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_141 <= 22'h0;
    end else if (_T_1764) begin
      btb_bank0_rd_data_way1_out_141 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_142 <= 22'h0;
    end else if (_T_1767) begin
      btb_bank0_rd_data_way1_out_142 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_143 <= 22'h0;
    end else if (_T_1770) begin
      btb_bank0_rd_data_way1_out_143 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_144 <= 22'h0;
    end else if (_T_1773) begin
      btb_bank0_rd_data_way1_out_144 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_145 <= 22'h0;
    end else if (_T_1776) begin
      btb_bank0_rd_data_way1_out_145 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_146 <= 22'h0;
    end else if (_T_1779) begin
      btb_bank0_rd_data_way1_out_146 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_147 <= 22'h0;
    end else if (_T_1782) begin
      btb_bank0_rd_data_way1_out_147 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_148 <= 22'h0;
    end else if (_T_1785) begin
      btb_bank0_rd_data_way1_out_148 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_149 <= 22'h0;
    end else if (_T_1788) begin
      btb_bank0_rd_data_way1_out_149 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_150 <= 22'h0;
    end else if (_T_1791) begin
      btb_bank0_rd_data_way1_out_150 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_151 <= 22'h0;
    end else if (_T_1794) begin
      btb_bank0_rd_data_way1_out_151 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_152 <= 22'h0;
    end else if (_T_1797) begin
      btb_bank0_rd_data_way1_out_152 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_153 <= 22'h0;
    end else if (_T_1800) begin
      btb_bank0_rd_data_way1_out_153 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_154 <= 22'h0;
    end else if (_T_1803) begin
      btb_bank0_rd_data_way1_out_154 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_155 <= 22'h0;
    end else if (_T_1806) begin
      btb_bank0_rd_data_way1_out_155 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_156 <= 22'h0;
    end else if (_T_1809) begin
      btb_bank0_rd_data_way1_out_156 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_157 <= 22'h0;
    end else if (_T_1812) begin
      btb_bank0_rd_data_way1_out_157 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_158 <= 22'h0;
    end else if (_T_1815) begin
      btb_bank0_rd_data_way1_out_158 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_159 <= 22'h0;
    end else if (_T_1818) begin
      btb_bank0_rd_data_way1_out_159 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_160 <= 22'h0;
    end else if (_T_1821) begin
      btb_bank0_rd_data_way1_out_160 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_161 <= 22'h0;
    end else if (_T_1824) begin
      btb_bank0_rd_data_way1_out_161 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_162 <= 22'h0;
    end else if (_T_1827) begin
      btb_bank0_rd_data_way1_out_162 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_163 <= 22'h0;
    end else if (_T_1830) begin
      btb_bank0_rd_data_way1_out_163 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_164 <= 22'h0;
    end else if (_T_1833) begin
      btb_bank0_rd_data_way1_out_164 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_165 <= 22'h0;
    end else if (_T_1836) begin
      btb_bank0_rd_data_way1_out_165 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_166 <= 22'h0;
    end else if (_T_1839) begin
      btb_bank0_rd_data_way1_out_166 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_167 <= 22'h0;
    end else if (_T_1842) begin
      btb_bank0_rd_data_way1_out_167 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_168 <= 22'h0;
    end else if (_T_1845) begin
      btb_bank0_rd_data_way1_out_168 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_169 <= 22'h0;
    end else if (_T_1848) begin
      btb_bank0_rd_data_way1_out_169 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_170 <= 22'h0;
    end else if (_T_1851) begin
      btb_bank0_rd_data_way1_out_170 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_171 <= 22'h0;
    end else if (_T_1854) begin
      btb_bank0_rd_data_way1_out_171 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_172 <= 22'h0;
    end else if (_T_1857) begin
      btb_bank0_rd_data_way1_out_172 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_173 <= 22'h0;
    end else if (_T_1860) begin
      btb_bank0_rd_data_way1_out_173 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_174 <= 22'h0;
    end else if (_T_1863) begin
      btb_bank0_rd_data_way1_out_174 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_175 <= 22'h0;
    end else if (_T_1866) begin
      btb_bank0_rd_data_way1_out_175 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_176 <= 22'h0;
    end else if (_T_1869) begin
      btb_bank0_rd_data_way1_out_176 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_177 <= 22'h0;
    end else if (_T_1872) begin
      btb_bank0_rd_data_way1_out_177 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_178 <= 22'h0;
    end else if (_T_1875) begin
      btb_bank0_rd_data_way1_out_178 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_179 <= 22'h0;
    end else if (_T_1878) begin
      btb_bank0_rd_data_way1_out_179 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_180 <= 22'h0;
    end else if (_T_1881) begin
      btb_bank0_rd_data_way1_out_180 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_181 <= 22'h0;
    end else if (_T_1884) begin
      btb_bank0_rd_data_way1_out_181 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_182 <= 22'h0;
    end else if (_T_1887) begin
      btb_bank0_rd_data_way1_out_182 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_183 <= 22'h0;
    end else if (_T_1890) begin
      btb_bank0_rd_data_way1_out_183 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_184 <= 22'h0;
    end else if (_T_1893) begin
      btb_bank0_rd_data_way1_out_184 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_185 <= 22'h0;
    end else if (_T_1896) begin
      btb_bank0_rd_data_way1_out_185 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_186 <= 22'h0;
    end else if (_T_1899) begin
      btb_bank0_rd_data_way1_out_186 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_187 <= 22'h0;
    end else if (_T_1902) begin
      btb_bank0_rd_data_way1_out_187 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_188 <= 22'h0;
    end else if (_T_1905) begin
      btb_bank0_rd_data_way1_out_188 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_189 <= 22'h0;
    end else if (_T_1908) begin
      btb_bank0_rd_data_way1_out_189 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_190 <= 22'h0;
    end else if (_T_1911) begin
      btb_bank0_rd_data_way1_out_190 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_191 <= 22'h0;
    end else if (_T_1914) begin
      btb_bank0_rd_data_way1_out_191 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_192 <= 22'h0;
    end else if (_T_1917) begin
      btb_bank0_rd_data_way1_out_192 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_193 <= 22'h0;
    end else if (_T_1920) begin
      btb_bank0_rd_data_way1_out_193 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_194 <= 22'h0;
    end else if (_T_1923) begin
      btb_bank0_rd_data_way1_out_194 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_195 <= 22'h0;
    end else if (_T_1926) begin
      btb_bank0_rd_data_way1_out_195 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_196 <= 22'h0;
    end else if (_T_1929) begin
      btb_bank0_rd_data_way1_out_196 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_197 <= 22'h0;
    end else if (_T_1932) begin
      btb_bank0_rd_data_way1_out_197 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_198 <= 22'h0;
    end else if (_T_1935) begin
      btb_bank0_rd_data_way1_out_198 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_199 <= 22'h0;
    end else if (_T_1938) begin
      btb_bank0_rd_data_way1_out_199 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_200 <= 22'h0;
    end else if (_T_1941) begin
      btb_bank0_rd_data_way1_out_200 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_201 <= 22'h0;
    end else if (_T_1944) begin
      btb_bank0_rd_data_way1_out_201 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_202 <= 22'h0;
    end else if (_T_1947) begin
      btb_bank0_rd_data_way1_out_202 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_203 <= 22'h0;
    end else if (_T_1950) begin
      btb_bank0_rd_data_way1_out_203 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_204 <= 22'h0;
    end else if (_T_1953) begin
      btb_bank0_rd_data_way1_out_204 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_205 <= 22'h0;
    end else if (_T_1956) begin
      btb_bank0_rd_data_way1_out_205 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_206 <= 22'h0;
    end else if (_T_1959) begin
      btb_bank0_rd_data_way1_out_206 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_207 <= 22'h0;
    end else if (_T_1962) begin
      btb_bank0_rd_data_way1_out_207 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_208 <= 22'h0;
    end else if (_T_1965) begin
      btb_bank0_rd_data_way1_out_208 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_209 <= 22'h0;
    end else if (_T_1968) begin
      btb_bank0_rd_data_way1_out_209 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_210 <= 22'h0;
    end else if (_T_1971) begin
      btb_bank0_rd_data_way1_out_210 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_211 <= 22'h0;
    end else if (_T_1974) begin
      btb_bank0_rd_data_way1_out_211 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_212 <= 22'h0;
    end else if (_T_1977) begin
      btb_bank0_rd_data_way1_out_212 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_213 <= 22'h0;
    end else if (_T_1980) begin
      btb_bank0_rd_data_way1_out_213 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_214 <= 22'h0;
    end else if (_T_1983) begin
      btb_bank0_rd_data_way1_out_214 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_215 <= 22'h0;
    end else if (_T_1986) begin
      btb_bank0_rd_data_way1_out_215 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_216 <= 22'h0;
    end else if (_T_1989) begin
      btb_bank0_rd_data_way1_out_216 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_217 <= 22'h0;
    end else if (_T_1992) begin
      btb_bank0_rd_data_way1_out_217 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_218 <= 22'h0;
    end else if (_T_1995) begin
      btb_bank0_rd_data_way1_out_218 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_219 <= 22'h0;
    end else if (_T_1998) begin
      btb_bank0_rd_data_way1_out_219 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_220 <= 22'h0;
    end else if (_T_2001) begin
      btb_bank0_rd_data_way1_out_220 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_221 <= 22'h0;
    end else if (_T_2004) begin
      btb_bank0_rd_data_way1_out_221 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_222 <= 22'h0;
    end else if (_T_2007) begin
      btb_bank0_rd_data_way1_out_222 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_223 <= 22'h0;
    end else if (_T_2010) begin
      btb_bank0_rd_data_way1_out_223 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_224 <= 22'h0;
    end else if (_T_2013) begin
      btb_bank0_rd_data_way1_out_224 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_225 <= 22'h0;
    end else if (_T_2016) begin
      btb_bank0_rd_data_way1_out_225 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_226 <= 22'h0;
    end else if (_T_2019) begin
      btb_bank0_rd_data_way1_out_226 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_227 <= 22'h0;
    end else if (_T_2022) begin
      btb_bank0_rd_data_way1_out_227 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_228 <= 22'h0;
    end else if (_T_2025) begin
      btb_bank0_rd_data_way1_out_228 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_229 <= 22'h0;
    end else if (_T_2028) begin
      btb_bank0_rd_data_way1_out_229 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_230 <= 22'h0;
    end else if (_T_2031) begin
      btb_bank0_rd_data_way1_out_230 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_231 <= 22'h0;
    end else if (_T_2034) begin
      btb_bank0_rd_data_way1_out_231 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_232 <= 22'h0;
    end else if (_T_2037) begin
      btb_bank0_rd_data_way1_out_232 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_233 <= 22'h0;
    end else if (_T_2040) begin
      btb_bank0_rd_data_way1_out_233 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_234 <= 22'h0;
    end else if (_T_2043) begin
      btb_bank0_rd_data_way1_out_234 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_235 <= 22'h0;
    end else if (_T_2046) begin
      btb_bank0_rd_data_way1_out_235 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_236 <= 22'h0;
    end else if (_T_2049) begin
      btb_bank0_rd_data_way1_out_236 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_237 <= 22'h0;
    end else if (_T_2052) begin
      btb_bank0_rd_data_way1_out_237 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_238 <= 22'h0;
    end else if (_T_2055) begin
      btb_bank0_rd_data_way1_out_238 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_239 <= 22'h0;
    end else if (_T_2058) begin
      btb_bank0_rd_data_way1_out_239 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_240 <= 22'h0;
    end else if (_T_2061) begin
      btb_bank0_rd_data_way1_out_240 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_241 <= 22'h0;
    end else if (_T_2064) begin
      btb_bank0_rd_data_way1_out_241 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_242 <= 22'h0;
    end else if (_T_2067) begin
      btb_bank0_rd_data_way1_out_242 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_243 <= 22'h0;
    end else if (_T_2070) begin
      btb_bank0_rd_data_way1_out_243 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_244 <= 22'h0;
    end else if (_T_2073) begin
      btb_bank0_rd_data_way1_out_244 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_245 <= 22'h0;
    end else if (_T_2076) begin
      btb_bank0_rd_data_way1_out_245 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_246 <= 22'h0;
    end else if (_T_2079) begin
      btb_bank0_rd_data_way1_out_246 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_247 <= 22'h0;
    end else if (_T_2082) begin
      btb_bank0_rd_data_way1_out_247 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_248 <= 22'h0;
    end else if (_T_2085) begin
      btb_bank0_rd_data_way1_out_248 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_249 <= 22'h0;
    end else if (_T_2088) begin
      btb_bank0_rd_data_way1_out_249 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_250 <= 22'h0;
    end else if (_T_2091) begin
      btb_bank0_rd_data_way1_out_250 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_251 <= 22'h0;
    end else if (_T_2094) begin
      btb_bank0_rd_data_way1_out_251 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_252 <= 22'h0;
    end else if (_T_2097) begin
      btb_bank0_rd_data_way1_out_252 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_253 <= 22'h0;
    end else if (_T_2100) begin
      btb_bank0_rd_data_way1_out_253 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_254 <= 22'h0;
    end else if (_T_2103) begin
      btb_bank0_rd_data_way1_out_254 <= btb_wr_data;
    end
    if (reset) begin
      btb_bank0_rd_data_way1_out_255 <= 22'h0;
    end else if (_T_2106) begin
      btb_bank0_rd_data_way1_out_255 <= btb_wr_data;
    end
    if (reset) begin
      fghr <= 8'h0;
    end else begin
      fghr <= fghr_ns;
    end
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_8514) begin
        bht_bank_rd_data_out_1_0 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_8658) begin
        bht_bank_rd_data_out_1_1 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_8802) begin
        bht_bank_rd_data_out_1_2 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_8946) begin
        bht_bank_rd_data_out_1_3 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_9090) begin
        bht_bank_rd_data_out_1_4 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_9234) begin
        bht_bank_rd_data_out_1_5 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_9378) begin
        bht_bank_rd_data_out_1_6 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_9522) begin
        bht_bank_rd_data_out_1_7 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_9666) begin
        bht_bank_rd_data_out_1_8 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_9810) begin
        bht_bank_rd_data_out_1_9 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_9954) begin
        bht_bank_rd_data_out_1_10 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_10098) begin
        bht_bank_rd_data_out_1_11 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_10242) begin
        bht_bank_rd_data_out_1_12 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_10386) begin
        bht_bank_rd_data_out_1_13 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_10530) begin
        bht_bank_rd_data_out_1_14 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_10674) begin
        bht_bank_rd_data_out_1_15 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_8523) begin
        bht_bank_rd_data_out_1_16 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_8667) begin
        bht_bank_rd_data_out_1_17 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_8811) begin
        bht_bank_rd_data_out_1_18 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_8955) begin
        bht_bank_rd_data_out_1_19 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_9099) begin
        bht_bank_rd_data_out_1_20 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_9243) begin
        bht_bank_rd_data_out_1_21 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_9387) begin
        bht_bank_rd_data_out_1_22 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_9531) begin
        bht_bank_rd_data_out_1_23 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_9675) begin
        bht_bank_rd_data_out_1_24 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_9819) begin
        bht_bank_rd_data_out_1_25 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_9963) begin
        bht_bank_rd_data_out_1_26 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_10107) begin
        bht_bank_rd_data_out_1_27 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_10251) begin
        bht_bank_rd_data_out_1_28 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_10395) begin
        bht_bank_rd_data_out_1_29 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_10539) begin
        bht_bank_rd_data_out_1_30 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_10683) begin
        bht_bank_rd_data_out_1_31 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_8532) begin
        bht_bank_rd_data_out_1_32 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_8676) begin
        bht_bank_rd_data_out_1_33 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_8820) begin
        bht_bank_rd_data_out_1_34 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_8964) begin
        bht_bank_rd_data_out_1_35 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_9108) begin
        bht_bank_rd_data_out_1_36 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_9252) begin
        bht_bank_rd_data_out_1_37 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_9396) begin
        bht_bank_rd_data_out_1_38 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_9540) begin
        bht_bank_rd_data_out_1_39 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_9684) begin
        bht_bank_rd_data_out_1_40 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_9828) begin
        bht_bank_rd_data_out_1_41 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_9972) begin
        bht_bank_rd_data_out_1_42 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_10116) begin
        bht_bank_rd_data_out_1_43 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_10260) begin
        bht_bank_rd_data_out_1_44 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_10404) begin
        bht_bank_rd_data_out_1_45 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_10548) begin
        bht_bank_rd_data_out_1_46 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_10692) begin
        bht_bank_rd_data_out_1_47 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_8541) begin
        bht_bank_rd_data_out_1_48 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_8685) begin
        bht_bank_rd_data_out_1_49 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_8829) begin
        bht_bank_rd_data_out_1_50 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_8973) begin
        bht_bank_rd_data_out_1_51 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_9117) begin
        bht_bank_rd_data_out_1_52 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_9261) begin
        bht_bank_rd_data_out_1_53 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_9405) begin
        bht_bank_rd_data_out_1_54 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_9549) begin
        bht_bank_rd_data_out_1_55 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_9693) begin
        bht_bank_rd_data_out_1_56 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_9837) begin
        bht_bank_rd_data_out_1_57 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_9981) begin
        bht_bank_rd_data_out_1_58 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_10125) begin
        bht_bank_rd_data_out_1_59 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_10269) begin
        bht_bank_rd_data_out_1_60 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_10413) begin
        bht_bank_rd_data_out_1_61 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_10557) begin
        bht_bank_rd_data_out_1_62 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_10701) begin
        bht_bank_rd_data_out_1_63 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_8550) begin
        bht_bank_rd_data_out_1_64 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_8694) begin
        bht_bank_rd_data_out_1_65 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_8838) begin
        bht_bank_rd_data_out_1_66 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_8982) begin
        bht_bank_rd_data_out_1_67 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_9126) begin
        bht_bank_rd_data_out_1_68 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_9270) begin
        bht_bank_rd_data_out_1_69 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_9414) begin
        bht_bank_rd_data_out_1_70 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_9558) begin
        bht_bank_rd_data_out_1_71 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_9702) begin
        bht_bank_rd_data_out_1_72 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_9846) begin
        bht_bank_rd_data_out_1_73 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_9990) begin
        bht_bank_rd_data_out_1_74 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_10134) begin
        bht_bank_rd_data_out_1_75 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_10278) begin
        bht_bank_rd_data_out_1_76 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_10422) begin
        bht_bank_rd_data_out_1_77 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_10566) begin
        bht_bank_rd_data_out_1_78 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_10710) begin
        bht_bank_rd_data_out_1_79 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_8559) begin
        bht_bank_rd_data_out_1_80 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_8703) begin
        bht_bank_rd_data_out_1_81 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_8847) begin
        bht_bank_rd_data_out_1_82 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_8991) begin
        bht_bank_rd_data_out_1_83 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_9135) begin
        bht_bank_rd_data_out_1_84 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_9279) begin
        bht_bank_rd_data_out_1_85 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_9423) begin
        bht_bank_rd_data_out_1_86 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_9567) begin
        bht_bank_rd_data_out_1_87 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_9711) begin
        bht_bank_rd_data_out_1_88 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_9855) begin
        bht_bank_rd_data_out_1_89 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_9999) begin
        bht_bank_rd_data_out_1_90 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_10143) begin
        bht_bank_rd_data_out_1_91 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_10287) begin
        bht_bank_rd_data_out_1_92 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_10431) begin
        bht_bank_rd_data_out_1_93 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_10575) begin
        bht_bank_rd_data_out_1_94 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_10719) begin
        bht_bank_rd_data_out_1_95 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_8568) begin
        bht_bank_rd_data_out_1_96 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_8712) begin
        bht_bank_rd_data_out_1_97 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_8856) begin
        bht_bank_rd_data_out_1_98 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9000) begin
        bht_bank_rd_data_out_1_99 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_9144) begin
        bht_bank_rd_data_out_1_100 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_9288) begin
        bht_bank_rd_data_out_1_101 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_9432) begin
        bht_bank_rd_data_out_1_102 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_9576) begin
        bht_bank_rd_data_out_1_103 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_9720) begin
        bht_bank_rd_data_out_1_104 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_9864) begin
        bht_bank_rd_data_out_1_105 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10008) begin
        bht_bank_rd_data_out_1_106 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_10152) begin
        bht_bank_rd_data_out_1_107 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_10296) begin
        bht_bank_rd_data_out_1_108 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_10440) begin
        bht_bank_rd_data_out_1_109 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_10584) begin
        bht_bank_rd_data_out_1_110 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_10728) begin
        bht_bank_rd_data_out_1_111 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_8577) begin
        bht_bank_rd_data_out_1_112 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_8721) begin
        bht_bank_rd_data_out_1_113 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_8865) begin
        bht_bank_rd_data_out_1_114 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9009) begin
        bht_bank_rd_data_out_1_115 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_9153) begin
        bht_bank_rd_data_out_1_116 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_9297) begin
        bht_bank_rd_data_out_1_117 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_9441) begin
        bht_bank_rd_data_out_1_118 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_9585) begin
        bht_bank_rd_data_out_1_119 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_9729) begin
        bht_bank_rd_data_out_1_120 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_9873) begin
        bht_bank_rd_data_out_1_121 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10017) begin
        bht_bank_rd_data_out_1_122 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_10161) begin
        bht_bank_rd_data_out_1_123 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_10305) begin
        bht_bank_rd_data_out_1_124 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_10449) begin
        bht_bank_rd_data_out_1_125 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_10593) begin
        bht_bank_rd_data_out_1_126 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_10737) begin
        bht_bank_rd_data_out_1_127 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_8586) begin
        bht_bank_rd_data_out_1_128 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_8730) begin
        bht_bank_rd_data_out_1_129 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_8874) begin
        bht_bank_rd_data_out_1_130 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9018) begin
        bht_bank_rd_data_out_1_131 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_9162) begin
        bht_bank_rd_data_out_1_132 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_9306) begin
        bht_bank_rd_data_out_1_133 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_9450) begin
        bht_bank_rd_data_out_1_134 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_9594) begin
        bht_bank_rd_data_out_1_135 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_9738) begin
        bht_bank_rd_data_out_1_136 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_9882) begin
        bht_bank_rd_data_out_1_137 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10026) begin
        bht_bank_rd_data_out_1_138 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_10170) begin
        bht_bank_rd_data_out_1_139 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_10314) begin
        bht_bank_rd_data_out_1_140 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_10458) begin
        bht_bank_rd_data_out_1_141 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_10602) begin
        bht_bank_rd_data_out_1_142 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_10746) begin
        bht_bank_rd_data_out_1_143 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_8595) begin
        bht_bank_rd_data_out_1_144 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_8739) begin
        bht_bank_rd_data_out_1_145 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_8883) begin
        bht_bank_rd_data_out_1_146 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9027) begin
        bht_bank_rd_data_out_1_147 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_9171) begin
        bht_bank_rd_data_out_1_148 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_9315) begin
        bht_bank_rd_data_out_1_149 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_9459) begin
        bht_bank_rd_data_out_1_150 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_9603) begin
        bht_bank_rd_data_out_1_151 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_9747) begin
        bht_bank_rd_data_out_1_152 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_9891) begin
        bht_bank_rd_data_out_1_153 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10035) begin
        bht_bank_rd_data_out_1_154 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_10179) begin
        bht_bank_rd_data_out_1_155 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_10323) begin
        bht_bank_rd_data_out_1_156 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_10467) begin
        bht_bank_rd_data_out_1_157 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_10611) begin
        bht_bank_rd_data_out_1_158 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_10755) begin
        bht_bank_rd_data_out_1_159 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_8604) begin
        bht_bank_rd_data_out_1_160 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_8748) begin
        bht_bank_rd_data_out_1_161 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_8892) begin
        bht_bank_rd_data_out_1_162 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9036) begin
        bht_bank_rd_data_out_1_163 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_9180) begin
        bht_bank_rd_data_out_1_164 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_9324) begin
        bht_bank_rd_data_out_1_165 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_9468) begin
        bht_bank_rd_data_out_1_166 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_9612) begin
        bht_bank_rd_data_out_1_167 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_9756) begin
        bht_bank_rd_data_out_1_168 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_9900) begin
        bht_bank_rd_data_out_1_169 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10044) begin
        bht_bank_rd_data_out_1_170 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_10188) begin
        bht_bank_rd_data_out_1_171 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_10332) begin
        bht_bank_rd_data_out_1_172 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_10476) begin
        bht_bank_rd_data_out_1_173 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_10620) begin
        bht_bank_rd_data_out_1_174 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_10764) begin
        bht_bank_rd_data_out_1_175 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_8613) begin
        bht_bank_rd_data_out_1_176 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_8757) begin
        bht_bank_rd_data_out_1_177 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_8901) begin
        bht_bank_rd_data_out_1_178 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9045) begin
        bht_bank_rd_data_out_1_179 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_9189) begin
        bht_bank_rd_data_out_1_180 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_9333) begin
        bht_bank_rd_data_out_1_181 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_9477) begin
        bht_bank_rd_data_out_1_182 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_9621) begin
        bht_bank_rd_data_out_1_183 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_9765) begin
        bht_bank_rd_data_out_1_184 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_9909) begin
        bht_bank_rd_data_out_1_185 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10053) begin
        bht_bank_rd_data_out_1_186 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_10197) begin
        bht_bank_rd_data_out_1_187 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_10341) begin
        bht_bank_rd_data_out_1_188 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_10485) begin
        bht_bank_rd_data_out_1_189 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_10629) begin
        bht_bank_rd_data_out_1_190 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_10773) begin
        bht_bank_rd_data_out_1_191 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_8622) begin
        bht_bank_rd_data_out_1_192 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_8766) begin
        bht_bank_rd_data_out_1_193 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_8910) begin
        bht_bank_rd_data_out_1_194 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9054) begin
        bht_bank_rd_data_out_1_195 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_9198) begin
        bht_bank_rd_data_out_1_196 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_9342) begin
        bht_bank_rd_data_out_1_197 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_9486) begin
        bht_bank_rd_data_out_1_198 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_9630) begin
        bht_bank_rd_data_out_1_199 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_9774) begin
        bht_bank_rd_data_out_1_200 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_9918) begin
        bht_bank_rd_data_out_1_201 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10062) begin
        bht_bank_rd_data_out_1_202 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_10206) begin
        bht_bank_rd_data_out_1_203 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_10350) begin
        bht_bank_rd_data_out_1_204 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_10494) begin
        bht_bank_rd_data_out_1_205 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_10638) begin
        bht_bank_rd_data_out_1_206 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_10782) begin
        bht_bank_rd_data_out_1_207 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_8631) begin
        bht_bank_rd_data_out_1_208 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_8775) begin
        bht_bank_rd_data_out_1_209 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_8919) begin
        bht_bank_rd_data_out_1_210 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9063) begin
        bht_bank_rd_data_out_1_211 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_9207) begin
        bht_bank_rd_data_out_1_212 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_9351) begin
        bht_bank_rd_data_out_1_213 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_9495) begin
        bht_bank_rd_data_out_1_214 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_9639) begin
        bht_bank_rd_data_out_1_215 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_9783) begin
        bht_bank_rd_data_out_1_216 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_9927) begin
        bht_bank_rd_data_out_1_217 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_10071) begin
        bht_bank_rd_data_out_1_218 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_10215) begin
        bht_bank_rd_data_out_1_219 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_10359) begin
        bht_bank_rd_data_out_1_220 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_10503) begin
        bht_bank_rd_data_out_1_221 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_10647) begin
        bht_bank_rd_data_out_1_222 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_10791) begin
        bht_bank_rd_data_out_1_223 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_8640) begin
        bht_bank_rd_data_out_1_224 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_8784) begin
        bht_bank_rd_data_out_1_225 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_8928) begin
        bht_bank_rd_data_out_1_226 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_9072) begin
        bht_bank_rd_data_out_1_227 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_9216) begin
        bht_bank_rd_data_out_1_228 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_9360) begin
        bht_bank_rd_data_out_1_229 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_9504) begin
        bht_bank_rd_data_out_1_230 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_9648) begin
        bht_bank_rd_data_out_1_231 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_9792) begin
        bht_bank_rd_data_out_1_232 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_9936) begin
        bht_bank_rd_data_out_1_233 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_10080) begin
        bht_bank_rd_data_out_1_234 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_10224) begin
        bht_bank_rd_data_out_1_235 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_10368) begin
        bht_bank_rd_data_out_1_236 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_10512) begin
        bht_bank_rd_data_out_1_237 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_10656) begin
        bht_bank_rd_data_out_1_238 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_10800) begin
        bht_bank_rd_data_out_1_239 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_8649) begin
        bht_bank_rd_data_out_1_240 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_8793) begin
        bht_bank_rd_data_out_1_241 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_8937) begin
        bht_bank_rd_data_out_1_242 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_9081) begin
        bht_bank_rd_data_out_1_243 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_9225) begin
        bht_bank_rd_data_out_1_244 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_9369) begin
        bht_bank_rd_data_out_1_245 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_9513) begin
        bht_bank_rd_data_out_1_246 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_9657) begin
        bht_bank_rd_data_out_1_247 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_9801) begin
        bht_bank_rd_data_out_1_248 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_9945) begin
        bht_bank_rd_data_out_1_249 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_10089) begin
        bht_bank_rd_data_out_1_250 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_10233) begin
        bht_bank_rd_data_out_1_251 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_10377) begin
        bht_bank_rd_data_out_1_252 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_10521) begin
        bht_bank_rd_data_out_1_253 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_10665) begin
        bht_bank_rd_data_out_1_254 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_10809) begin
        bht_bank_rd_data_out_1_255 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_6210) begin
        bht_bank_rd_data_out_0_0 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_6354) begin
        bht_bank_rd_data_out_0_1 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_6498) begin
        bht_bank_rd_data_out_0_2 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_6642) begin
        bht_bank_rd_data_out_0_3 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_6786) begin
        bht_bank_rd_data_out_0_4 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_6930) begin
        bht_bank_rd_data_out_0_5 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_7074) begin
        bht_bank_rd_data_out_0_6 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_7218) begin
        bht_bank_rd_data_out_0_7 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_7362) begin
        bht_bank_rd_data_out_0_8 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_7506) begin
        bht_bank_rd_data_out_0_9 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_7650) begin
        bht_bank_rd_data_out_0_10 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_7794) begin
        bht_bank_rd_data_out_0_11 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_7938) begin
        bht_bank_rd_data_out_0_12 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_8082) begin
        bht_bank_rd_data_out_0_13 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_8226) begin
        bht_bank_rd_data_out_0_14 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_8370) begin
        bht_bank_rd_data_out_0_15 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_6219) begin
        bht_bank_rd_data_out_0_16 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_6363) begin
        bht_bank_rd_data_out_0_17 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_6507) begin
        bht_bank_rd_data_out_0_18 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_6651) begin
        bht_bank_rd_data_out_0_19 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_6795) begin
        bht_bank_rd_data_out_0_20 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_6939) begin
        bht_bank_rd_data_out_0_21 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_7083) begin
        bht_bank_rd_data_out_0_22 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_7227) begin
        bht_bank_rd_data_out_0_23 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_7371) begin
        bht_bank_rd_data_out_0_24 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_7515) begin
        bht_bank_rd_data_out_0_25 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_7659) begin
        bht_bank_rd_data_out_0_26 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_7803) begin
        bht_bank_rd_data_out_0_27 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_7947) begin
        bht_bank_rd_data_out_0_28 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_8091) begin
        bht_bank_rd_data_out_0_29 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_8235) begin
        bht_bank_rd_data_out_0_30 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_8379) begin
        bht_bank_rd_data_out_0_31 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_6228) begin
        bht_bank_rd_data_out_0_32 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_6372) begin
        bht_bank_rd_data_out_0_33 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_6516) begin
        bht_bank_rd_data_out_0_34 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_6660) begin
        bht_bank_rd_data_out_0_35 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_6804) begin
        bht_bank_rd_data_out_0_36 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_6948) begin
        bht_bank_rd_data_out_0_37 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_7092) begin
        bht_bank_rd_data_out_0_38 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_7236) begin
        bht_bank_rd_data_out_0_39 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_7380) begin
        bht_bank_rd_data_out_0_40 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_7524) begin
        bht_bank_rd_data_out_0_41 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_7668) begin
        bht_bank_rd_data_out_0_42 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_7812) begin
        bht_bank_rd_data_out_0_43 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_7956) begin
        bht_bank_rd_data_out_0_44 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_8100) begin
        bht_bank_rd_data_out_0_45 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_8244) begin
        bht_bank_rd_data_out_0_46 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_8388) begin
        bht_bank_rd_data_out_0_47 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_6237) begin
        bht_bank_rd_data_out_0_48 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_6381) begin
        bht_bank_rd_data_out_0_49 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_6525) begin
        bht_bank_rd_data_out_0_50 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_6669) begin
        bht_bank_rd_data_out_0_51 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_6813) begin
        bht_bank_rd_data_out_0_52 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_6957) begin
        bht_bank_rd_data_out_0_53 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_7101) begin
        bht_bank_rd_data_out_0_54 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_7245) begin
        bht_bank_rd_data_out_0_55 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_7389) begin
        bht_bank_rd_data_out_0_56 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_7533) begin
        bht_bank_rd_data_out_0_57 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_7677) begin
        bht_bank_rd_data_out_0_58 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_7821) begin
        bht_bank_rd_data_out_0_59 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_7965) begin
        bht_bank_rd_data_out_0_60 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_8109) begin
        bht_bank_rd_data_out_0_61 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_8253) begin
        bht_bank_rd_data_out_0_62 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_8397) begin
        bht_bank_rd_data_out_0_63 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_6246) begin
        bht_bank_rd_data_out_0_64 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_6390) begin
        bht_bank_rd_data_out_0_65 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_6534) begin
        bht_bank_rd_data_out_0_66 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_6678) begin
        bht_bank_rd_data_out_0_67 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_6822) begin
        bht_bank_rd_data_out_0_68 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_6966) begin
        bht_bank_rd_data_out_0_69 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_7110) begin
        bht_bank_rd_data_out_0_70 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_7254) begin
        bht_bank_rd_data_out_0_71 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_7398) begin
        bht_bank_rd_data_out_0_72 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_7542) begin
        bht_bank_rd_data_out_0_73 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_7686) begin
        bht_bank_rd_data_out_0_74 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_7830) begin
        bht_bank_rd_data_out_0_75 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_7974) begin
        bht_bank_rd_data_out_0_76 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_8118) begin
        bht_bank_rd_data_out_0_77 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_8262) begin
        bht_bank_rd_data_out_0_78 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_8406) begin
        bht_bank_rd_data_out_0_79 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_6255) begin
        bht_bank_rd_data_out_0_80 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_6399) begin
        bht_bank_rd_data_out_0_81 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_6543) begin
        bht_bank_rd_data_out_0_82 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_6687) begin
        bht_bank_rd_data_out_0_83 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_6831) begin
        bht_bank_rd_data_out_0_84 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_6975) begin
        bht_bank_rd_data_out_0_85 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_7119) begin
        bht_bank_rd_data_out_0_86 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_7263) begin
        bht_bank_rd_data_out_0_87 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_7407) begin
        bht_bank_rd_data_out_0_88 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_7551) begin
        bht_bank_rd_data_out_0_89 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_7695) begin
        bht_bank_rd_data_out_0_90 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_7839) begin
        bht_bank_rd_data_out_0_91 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_7983) begin
        bht_bank_rd_data_out_0_92 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_8127) begin
        bht_bank_rd_data_out_0_93 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_8271) begin
        bht_bank_rd_data_out_0_94 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_8415) begin
        bht_bank_rd_data_out_0_95 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_6264) begin
        bht_bank_rd_data_out_0_96 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_6408) begin
        bht_bank_rd_data_out_0_97 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_6552) begin
        bht_bank_rd_data_out_0_98 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_6696) begin
        bht_bank_rd_data_out_0_99 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_6840) begin
        bht_bank_rd_data_out_0_100 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_6984) begin
        bht_bank_rd_data_out_0_101 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_7128) begin
        bht_bank_rd_data_out_0_102 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_7272) begin
        bht_bank_rd_data_out_0_103 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_7416) begin
        bht_bank_rd_data_out_0_104 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_7560) begin
        bht_bank_rd_data_out_0_105 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_7704) begin
        bht_bank_rd_data_out_0_106 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_7848) begin
        bht_bank_rd_data_out_0_107 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_7992) begin
        bht_bank_rd_data_out_0_108 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_8136) begin
        bht_bank_rd_data_out_0_109 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_8280) begin
        bht_bank_rd_data_out_0_110 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_8424) begin
        bht_bank_rd_data_out_0_111 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_6273) begin
        bht_bank_rd_data_out_0_112 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_6417) begin
        bht_bank_rd_data_out_0_113 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_6561) begin
        bht_bank_rd_data_out_0_114 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_6705) begin
        bht_bank_rd_data_out_0_115 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_6849) begin
        bht_bank_rd_data_out_0_116 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_6993) begin
        bht_bank_rd_data_out_0_117 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_7137) begin
        bht_bank_rd_data_out_0_118 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_7281) begin
        bht_bank_rd_data_out_0_119 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_7425) begin
        bht_bank_rd_data_out_0_120 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_7569) begin
        bht_bank_rd_data_out_0_121 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_7713) begin
        bht_bank_rd_data_out_0_122 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_7857) begin
        bht_bank_rd_data_out_0_123 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8001) begin
        bht_bank_rd_data_out_0_124 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_8145) begin
        bht_bank_rd_data_out_0_125 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_8289) begin
        bht_bank_rd_data_out_0_126 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_8433) begin
        bht_bank_rd_data_out_0_127 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_6282) begin
        bht_bank_rd_data_out_0_128 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_6426) begin
        bht_bank_rd_data_out_0_129 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_6570) begin
        bht_bank_rd_data_out_0_130 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_6714) begin
        bht_bank_rd_data_out_0_131 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_6858) begin
        bht_bank_rd_data_out_0_132 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7002) begin
        bht_bank_rd_data_out_0_133 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_7146) begin
        bht_bank_rd_data_out_0_134 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_7290) begin
        bht_bank_rd_data_out_0_135 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_7434) begin
        bht_bank_rd_data_out_0_136 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_7578) begin
        bht_bank_rd_data_out_0_137 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_7722) begin
        bht_bank_rd_data_out_0_138 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_7866) begin
        bht_bank_rd_data_out_0_139 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8010) begin
        bht_bank_rd_data_out_0_140 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_8154) begin
        bht_bank_rd_data_out_0_141 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_8298) begin
        bht_bank_rd_data_out_0_142 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_8442) begin
        bht_bank_rd_data_out_0_143 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_6291) begin
        bht_bank_rd_data_out_0_144 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_6435) begin
        bht_bank_rd_data_out_0_145 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_6579) begin
        bht_bank_rd_data_out_0_146 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_6723) begin
        bht_bank_rd_data_out_0_147 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_6867) begin
        bht_bank_rd_data_out_0_148 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7011) begin
        bht_bank_rd_data_out_0_149 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_7155) begin
        bht_bank_rd_data_out_0_150 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_7299) begin
        bht_bank_rd_data_out_0_151 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_7443) begin
        bht_bank_rd_data_out_0_152 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_7587) begin
        bht_bank_rd_data_out_0_153 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_7731) begin
        bht_bank_rd_data_out_0_154 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_7875) begin
        bht_bank_rd_data_out_0_155 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8019) begin
        bht_bank_rd_data_out_0_156 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_8163) begin
        bht_bank_rd_data_out_0_157 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_8307) begin
        bht_bank_rd_data_out_0_158 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_8451) begin
        bht_bank_rd_data_out_0_159 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_6300) begin
        bht_bank_rd_data_out_0_160 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_6444) begin
        bht_bank_rd_data_out_0_161 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_6588) begin
        bht_bank_rd_data_out_0_162 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_6732) begin
        bht_bank_rd_data_out_0_163 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_6876) begin
        bht_bank_rd_data_out_0_164 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7020) begin
        bht_bank_rd_data_out_0_165 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_7164) begin
        bht_bank_rd_data_out_0_166 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_7308) begin
        bht_bank_rd_data_out_0_167 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_7452) begin
        bht_bank_rd_data_out_0_168 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_7596) begin
        bht_bank_rd_data_out_0_169 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_7740) begin
        bht_bank_rd_data_out_0_170 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_7884) begin
        bht_bank_rd_data_out_0_171 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8028) begin
        bht_bank_rd_data_out_0_172 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_8172) begin
        bht_bank_rd_data_out_0_173 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_8316) begin
        bht_bank_rd_data_out_0_174 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_8460) begin
        bht_bank_rd_data_out_0_175 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_6309) begin
        bht_bank_rd_data_out_0_176 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_6453) begin
        bht_bank_rd_data_out_0_177 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_6597) begin
        bht_bank_rd_data_out_0_178 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_6741) begin
        bht_bank_rd_data_out_0_179 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_6885) begin
        bht_bank_rd_data_out_0_180 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7029) begin
        bht_bank_rd_data_out_0_181 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_7173) begin
        bht_bank_rd_data_out_0_182 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_7317) begin
        bht_bank_rd_data_out_0_183 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_7461) begin
        bht_bank_rd_data_out_0_184 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_7605) begin
        bht_bank_rd_data_out_0_185 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_7749) begin
        bht_bank_rd_data_out_0_186 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_7893) begin
        bht_bank_rd_data_out_0_187 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8037) begin
        bht_bank_rd_data_out_0_188 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_8181) begin
        bht_bank_rd_data_out_0_189 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_8325) begin
        bht_bank_rd_data_out_0_190 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_8469) begin
        bht_bank_rd_data_out_0_191 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_6318) begin
        bht_bank_rd_data_out_0_192 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_6462) begin
        bht_bank_rd_data_out_0_193 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_6606) begin
        bht_bank_rd_data_out_0_194 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_6750) begin
        bht_bank_rd_data_out_0_195 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_6894) begin
        bht_bank_rd_data_out_0_196 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7038) begin
        bht_bank_rd_data_out_0_197 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_7182) begin
        bht_bank_rd_data_out_0_198 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_7326) begin
        bht_bank_rd_data_out_0_199 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_7470) begin
        bht_bank_rd_data_out_0_200 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_7614) begin
        bht_bank_rd_data_out_0_201 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_7758) begin
        bht_bank_rd_data_out_0_202 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_7902) begin
        bht_bank_rd_data_out_0_203 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8046) begin
        bht_bank_rd_data_out_0_204 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_8190) begin
        bht_bank_rd_data_out_0_205 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_8334) begin
        bht_bank_rd_data_out_0_206 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_8478) begin
        bht_bank_rd_data_out_0_207 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_6327) begin
        bht_bank_rd_data_out_0_208 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_6471) begin
        bht_bank_rd_data_out_0_209 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_6615) begin
        bht_bank_rd_data_out_0_210 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_6759) begin
        bht_bank_rd_data_out_0_211 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_6903) begin
        bht_bank_rd_data_out_0_212 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7047) begin
        bht_bank_rd_data_out_0_213 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_7191) begin
        bht_bank_rd_data_out_0_214 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_7335) begin
        bht_bank_rd_data_out_0_215 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_7479) begin
        bht_bank_rd_data_out_0_216 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_7623) begin
        bht_bank_rd_data_out_0_217 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_7767) begin
        bht_bank_rd_data_out_0_218 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_7911) begin
        bht_bank_rd_data_out_0_219 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8055) begin
        bht_bank_rd_data_out_0_220 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_8199) begin
        bht_bank_rd_data_out_0_221 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_8343) begin
        bht_bank_rd_data_out_0_222 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_8487) begin
        bht_bank_rd_data_out_0_223 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_6336) begin
        bht_bank_rd_data_out_0_224 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_6480) begin
        bht_bank_rd_data_out_0_225 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_6624) begin
        bht_bank_rd_data_out_0_226 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_6768) begin
        bht_bank_rd_data_out_0_227 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_6912) begin
        bht_bank_rd_data_out_0_228 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7056) begin
        bht_bank_rd_data_out_0_229 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_7200) begin
        bht_bank_rd_data_out_0_230 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_7344) begin
        bht_bank_rd_data_out_0_231 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_7488) begin
        bht_bank_rd_data_out_0_232 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_7632) begin
        bht_bank_rd_data_out_0_233 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_7776) begin
        bht_bank_rd_data_out_0_234 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_7920) begin
        bht_bank_rd_data_out_0_235 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8064) begin
        bht_bank_rd_data_out_0_236 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_8208) begin
        bht_bank_rd_data_out_0_237 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_8352) begin
        bht_bank_rd_data_out_0_238 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_8496) begin
        bht_bank_rd_data_out_0_239 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_6345) begin
        bht_bank_rd_data_out_0_240 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_6489) begin
        bht_bank_rd_data_out_0_241 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_6633) begin
        bht_bank_rd_data_out_0_242 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_6777) begin
        bht_bank_rd_data_out_0_243 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_6921) begin
        bht_bank_rd_data_out_0_244 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_7065) begin
        bht_bank_rd_data_out_0_245 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_7209) begin
        bht_bank_rd_data_out_0_246 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_7353) begin
        bht_bank_rd_data_out_0_247 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_7497) begin
        bht_bank_rd_data_out_0_248 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_7641) begin
        bht_bank_rd_data_out_0_249 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_7785) begin
        bht_bank_rd_data_out_0_250 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_7929) begin
        bht_bank_rd_data_out_0_251 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_8073) begin
        bht_bank_rd_data_out_0_252 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_8217) begin
        bht_bank_rd_data_out_0_253 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_8361) begin
        bht_bank_rd_data_out_0_254 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_8505) begin
        bht_bank_rd_data_out_0_255 <= io_dec_tlu_br0_r_pkt_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_mp_pkt_hist;
      end
    end
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else begin
      exu_mp_way_f <= io_exu_mp_pkt_way;
    end
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else if (_T_213) begin
      btb_lru_b0_f <= btb_lru_b0_ns;
    end
    if (reset) begin
      ifc_fetch_adder_prior <= 31'h0;
    end else if (_T_373) begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f;
    end
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else if (rsenable_0) begin
      rets_out_0 <= rets_in_0;
    end
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_1 <= rets_in_1;
    end
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_2 <= rets_in_2;
    end
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_3 <= rets_in_3;
    end
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_4 <= rets_in_4;
    end
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_5 <= rets_in_5;
    end
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_6 <= rets_in_6;
    end
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else if (rs_push) begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
