module rvecc_encode_64(
  input  [63:0] io_din,
  output [6:0]  io_ecc_out
);
  wire  w0_0 = io_din[0]; // @[el2_lib.scala 343:39]
  wire  w0_1 = io_din[1]; // @[el2_lib.scala 343:39]
  wire  w1_1 = io_din[2]; // @[el2_lib.scala 344:39]
  wire  w0_2 = io_din[3]; // @[el2_lib.scala 343:39]
  wire  w0_3 = io_din[4]; // @[el2_lib.scala 343:39]
  wire  w1_3 = io_din[5]; // @[el2_lib.scala 344:39]
  wire  w0_4 = io_din[6]; // @[el2_lib.scala 343:39]
  wire  w2_3 = io_din[7]; // @[el2_lib.scala 345:39]
  wire  w0_5 = io_din[8]; // @[el2_lib.scala 343:39]
  wire  w1_5 = io_din[9]; // @[el2_lib.scala 344:39]
  wire  w0_6 = io_din[10]; // @[el2_lib.scala 343:39]
  wire  w0_7 = io_din[11]; // @[el2_lib.scala 343:39]
  wire  w1_7 = io_din[12]; // @[el2_lib.scala 344:39]
  wire  w0_8 = io_din[13]; // @[el2_lib.scala 343:39]
  wire  w2_7 = io_din[14]; // @[el2_lib.scala 345:39]
  wire  w0_9 = io_din[15]; // @[el2_lib.scala 343:39]
  wire  w1_9 = io_din[16]; // @[el2_lib.scala 344:39]
  wire  w0_10 = io_din[17]; // @[el2_lib.scala 343:39]
  wire  w3_7 = io_din[18]; // @[el2_lib.scala 346:39]
  wire  w0_11 = io_din[19]; // @[el2_lib.scala 343:39]
  wire  w1_11 = io_din[20]; // @[el2_lib.scala 344:39]
  wire  w0_12 = io_din[21]; // @[el2_lib.scala 343:39]
  wire  w2_11 = io_din[22]; // @[el2_lib.scala 345:39]
  wire  w0_13 = io_din[23]; // @[el2_lib.scala 343:39]
  wire  w1_13 = io_din[24]; // @[el2_lib.scala 344:39]
  wire  w0_14 = io_din[25]; // @[el2_lib.scala 343:39]
  wire  w0_15 = io_din[26]; // @[el2_lib.scala 343:39]
  wire  w1_15 = io_din[27]; // @[el2_lib.scala 344:39]
  wire  w0_16 = io_din[28]; // @[el2_lib.scala 343:39]
  wire  w2_15 = io_din[29]; // @[el2_lib.scala 345:39]
  wire  w0_17 = io_din[30]; // @[el2_lib.scala 343:39]
  wire  w1_17 = io_din[31]; // @[el2_lib.scala 344:39]
  wire  w0_18 = io_din[32]; // @[el2_lib.scala 343:39]
  wire  w3_15 = io_din[33]; // @[el2_lib.scala 346:39]
  wire  w0_19 = io_din[34]; // @[el2_lib.scala 343:39]
  wire  w1_19 = io_din[35]; // @[el2_lib.scala 344:39]
  wire  w0_20 = io_din[36]; // @[el2_lib.scala 343:39]
  wire  w2_19 = io_din[37]; // @[el2_lib.scala 345:39]
  wire  w0_21 = io_din[38]; // @[el2_lib.scala 343:39]
  wire  w1_21 = io_din[39]; // @[el2_lib.scala 344:39]
  wire  w0_22 = io_din[40]; // @[el2_lib.scala 343:39]
  wire  w4_15 = io_din[41]; // @[el2_lib.scala 347:39]
  wire  w0_23 = io_din[42]; // @[el2_lib.scala 343:39]
  wire  w1_23 = io_din[43]; // @[el2_lib.scala 344:39]
  wire  w0_24 = io_din[44]; // @[el2_lib.scala 343:39]
  wire  w2_23 = io_din[45]; // @[el2_lib.scala 345:39]
  wire  w0_25 = io_din[46]; // @[el2_lib.scala 343:39]
  wire  w1_25 = io_din[47]; // @[el2_lib.scala 344:39]
  wire  w0_26 = io_din[48]; // @[el2_lib.scala 343:39]
  wire  w3_23 = io_din[49]; // @[el2_lib.scala 346:39]
  wire  w0_27 = io_din[50]; // @[el2_lib.scala 343:39]
  wire  w1_27 = io_din[51]; // @[el2_lib.scala 344:39]
  wire  w0_28 = io_din[52]; // @[el2_lib.scala 343:39]
  wire  w2_27 = io_din[53]; // @[el2_lib.scala 345:39]
  wire  w0_29 = io_din[54]; // @[el2_lib.scala 343:39]
  wire  w1_29 = io_din[55]; // @[el2_lib.scala 344:39]
  wire  w0_30 = io_din[56]; // @[el2_lib.scala 343:39]
  wire  w0_31 = io_din[57]; // @[el2_lib.scala 343:39]
  wire  w1_31 = io_din[58]; // @[el2_lib.scala 344:39]
  wire  w0_32 = io_din[59]; // @[el2_lib.scala 343:39]
  wire  w2_31 = io_din[60]; // @[el2_lib.scala 345:39]
  wire  w0_33 = io_din[61]; // @[el2_lib.scala 343:39]
  wire  w1_33 = io_din[62]; // @[el2_lib.scala 344:39]
  wire  w0_34 = io_din[63]; // @[el2_lib.scala 343:39]
  wire [6:0] _T_210 = {w0_34,w1_33,w0_33,w2_31,w0_32,w1_31,w0_31}; // @[el2_lib.scala 351:27]
  wire  _T_211 = ^_T_210; // @[el2_lib.scala 351:34]
  wire [6:0] _T_217 = {w0_18,w1_17,w0_17,w2_15,w0_16,w1_15,w0_15}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_224 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15}; // @[el2_lib.scala 351:44]
  wire [14:0] _T_225 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15,_T_217}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_232 = {w0_26,w1_25,w0_25,w2_23,w0_24,w1_23,w0_23,w4_15}; // @[el2_lib.scala 351:44]
  wire [30:0] _T_241 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_225}; // @[el2_lib.scala 351:44]
  wire  _T_242 = ^_T_241; // @[el2_lib.scala 351:51]
  wire [6:0] _T_248 = {w0_10,w1_9,w0_9,w2_7,w0_8,w1_7,w0_7}; // @[el2_lib.scala 351:61]
  wire [14:0] _T_256 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_248}; // @[el2_lib.scala 351:61]
  wire [30:0] _T_272 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_256}; // @[el2_lib.scala 351:61]
  wire  _T_273 = ^_T_272; // @[el2_lib.scala 351:68]
  wire [6:0] _T_279 = {w0_6,w1_5,w0_5,w2_3,w0_4,w1_3,w0_3}; // @[el2_lib.scala 351:78]
  wire [14:0] _T_287 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_279}; // @[el2_lib.scala 351:78]
  wire [30:0] _T_303 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_224,_T_287}; // @[el2_lib.scala 351:78]
  wire  _T_304 = ^_T_303; // @[el2_lib.scala 351:85]
  wire [7:0] _T_311 = {w2_7,w0_6,w1_5,w0_5,w2_3,w0_2,w1_1,w0_1}; // @[el2_lib.scala 351:95]
  wire [16:0] _T_320 = {w0_17,w2_15,w0_14,w1_13,w0_13,w2_11,w0_10,w1_9,w0_9,_T_311}; // @[el2_lib.scala 351:95]
  wire [8:0] _T_328 = {w1_25,w0_25,w2_23,w0_22,w1_21,w0_21,w2_19,w0_18,w1_17}; // @[el2_lib.scala 351:95]
  wire [17:0] _T_337 = {w0_34,w1_33,w0_33,w2_31,w0_30,w1_29,w0_29,w2_27,w0_26,_T_328}; // @[el2_lib.scala 351:95]
  wire [34:0] _T_338 = {_T_337,_T_320}; // @[el2_lib.scala 351:95]
  wire  _T_339 = ^_T_338; // @[el2_lib.scala 351:102]
  wire [7:0] _T_346 = {w1_7,w0_6,w1_5,w0_4,w1_3,w0_2,w1_1,w0_0}; // @[el2_lib.scala 351:112]
  wire [16:0] _T_355 = {w0_16,w1_15,w0_14,w1_13,w0_12,w1_11,w0_10,w1_9,w0_8,_T_346}; // @[el2_lib.scala 351:112]
  wire [8:0] _T_363 = {w1_25,w0_24,w1_23,w0_22,w1_21,w0_20,w1_19,w0_18,w1_17}; // @[el2_lib.scala 351:112]
  wire [17:0] _T_372 = {w0_34,w1_33,w0_32,w1_31,w0_30,w1_29,w0_28,w1_27,w0_26,_T_363}; // @[el2_lib.scala 351:112]
  wire [34:0] _T_373 = {_T_372,_T_355}; // @[el2_lib.scala 351:112]
  wire  _T_374 = ^_T_373; // @[el2_lib.scala 351:119]
  wire [7:0] _T_381 = {w0_7,w0_6,w0_5,w0_4,w0_3,w0_2,w0_1,w0_0}; // @[el2_lib.scala 351:129]
  wire [16:0] _T_390 = {w0_16,w0_15,w0_14,w0_13,w0_12,w0_11,w0_10,w0_9,w0_8,_T_381}; // @[el2_lib.scala 351:129]
  wire [8:0] _T_398 = {w0_25,w0_24,w0_23,w0_22,w0_21,w0_20,w0_19,w0_18,w0_17}; // @[el2_lib.scala 351:129]
  wire [17:0] _T_407 = {w0_34,w0_33,w0_32,w0_31,w0_30,w0_29,w0_28,w0_27,w0_26,_T_398}; // @[el2_lib.scala 351:129]
  wire [34:0] _T_408 = {_T_407,_T_390}; // @[el2_lib.scala 351:129]
  wire  _T_409 = ^_T_408; // @[el2_lib.scala 351:136]
  wire [2:0] _T_411 = {_T_339,_T_374,_T_409}; // @[Cat.scala 29:58]
  wire [3:0] _T_414 = {_T_211,_T_242,_T_273,_T_304}; // @[Cat.scala 29:58]
  assign io_ecc_out = {_T_414,_T_411}; // @[el2_lib.scala 351:16]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode,
  output [6:0]  io_ic_miss_buff_ecc,
  output [6:0]  io_ic_wr_ecc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] m1_io_din; // @[el2_ifu_mem_ctl.scala 343:18]
  wire [6:0] m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 343:18]
  wire [63:0] m2_io_din; // @[el2_ifu_mem_ctl.scala 344:18]
  wire [6:0] m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 344:18]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 185:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 321:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 322:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 322:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 254:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 556:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 558:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 187:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 309:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 673:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 673:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 676:91]
  wire [1:0] _T_2239 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 676:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 323:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 276:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 676:113]
  wire [1:0] _T_2240 = _T_2239 & _GEN_465; // @[el2_ifu_mem_ctl.scala 676:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 662:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 676:130]
  wire [1:0] _T_2241 = _T_2240 | _GEN_466; // @[el2_ifu_mem_ctl.scala 676:130]
  wire  _T_2242 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 676:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_2242}; // @[el2_ifu_mem_ctl.scala 676:152]
  wire [1:0] _T_2243 = _T_2241 & _GEN_467; // @[el2_ifu_mem_ctl.scala 676:152]
  wire [1:0] _T_2232 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 676:91]
  wire [1:0] _T_2233 = _T_2232 & _GEN_465; // @[el2_ifu_mem_ctl.scala 676:113]
  wire [1:0] _T_2234 = _T_2233 | _GEN_466; // @[el2_ifu_mem_ctl.scala 676:130]
  wire [1:0] _T_2236 = _T_2234 & _GEN_467; // @[el2_ifu_mem_ctl.scala 676:152]
  wire [3:0] iccm_ecc_word_enable = {_T_2243,_T_2236}; // @[Cat.scala 29:58]
  wire  _T_2343 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_2344 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_2345 = _T_2343 ^ _T_2344; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2353 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_2354 = ^_T_2353; // @[el2_lib.scala 301:83]
  wire  _T_2355 = io_iccm_rd_data_ecc[37] ^ _T_2354; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2362 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2370 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2362}; // @[el2_lib.scala 301:103]
  wire  _T_2371 = ^_T_2370; // @[el2_lib.scala 301:110]
  wire  _T_2372 = io_iccm_rd_data_ecc[36] ^ _T_2371; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2379 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2387 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2379}; // @[el2_lib.scala 301:130]
  wire  _T_2388 = ^_T_2387; // @[el2_lib.scala 301:137]
  wire  _T_2389 = io_iccm_rd_data_ecc[35] ^ _T_2388; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2398 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2407 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2398}; // @[el2_lib.scala 301:157]
  wire  _T_2408 = ^_T_2407; // @[el2_lib.scala 301:164]
  wire  _T_2409 = io_iccm_rd_data_ecc[34] ^ _T_2408; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2418 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2427 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2418}; // @[el2_lib.scala 301:184]
  wire  _T_2428 = ^_T_2427; // @[el2_lib.scala 301:191]
  wire  _T_2429 = io_iccm_rd_data_ecc[33] ^ _T_2428; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2438 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2447 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_2438}; // @[el2_lib.scala 301:211]
  wire  _T_2448 = ^_T_2447; // @[el2_lib.scala 301:218]
  wire  _T_2449 = io_iccm_rd_data_ecc[32] ^ _T_2448; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2455 = {_T_2345,_T_2355,_T_2372,_T_2389,_T_2409,_T_2429,_T_2449}; // @[Cat.scala 29:58]
  wire  _T_2456 = _T_2455 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2457 = iccm_ecc_word_enable[0] & _T_2456; // @[el2_lib.scala 302:32]
  wire  _T_2459 = _T_2457 & _T_2455[6]; // @[el2_lib.scala 302:53]
  wire  _T_2728 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_2729 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_2730 = _T_2728 ^ _T_2729; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2738 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_2739 = ^_T_2738; // @[el2_lib.scala 301:83]
  wire  _T_2740 = io_iccm_rd_data_ecc[76] ^ _T_2739; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2747 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2755 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2747}; // @[el2_lib.scala 301:103]
  wire  _T_2756 = ^_T_2755; // @[el2_lib.scala 301:110]
  wire  _T_2757 = io_iccm_rd_data_ecc[75] ^ _T_2756; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2764 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2772 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2764}; // @[el2_lib.scala 301:130]
  wire  _T_2773 = ^_T_2772; // @[el2_lib.scala 301:137]
  wire  _T_2774 = io_iccm_rd_data_ecc[74] ^ _T_2773; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2783 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2792 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2783}; // @[el2_lib.scala 301:157]
  wire  _T_2793 = ^_T_2792; // @[el2_lib.scala 301:164]
  wire  _T_2794 = io_iccm_rd_data_ecc[73] ^ _T_2793; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2803 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2812 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2803}; // @[el2_lib.scala 301:184]
  wire  _T_2813 = ^_T_2812; // @[el2_lib.scala 301:191]
  wire  _T_2814 = io_iccm_rd_data_ecc[72] ^ _T_2813; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2823 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2832 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_2823}; // @[el2_lib.scala 301:211]
  wire  _T_2833 = ^_T_2832; // @[el2_lib.scala 301:218]
  wire  _T_2834 = io_iccm_rd_data_ecc[71] ^ _T_2833; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2840 = {_T_2730,_T_2740,_T_2757,_T_2774,_T_2794,_T_2814,_T_2834}; // @[Cat.scala 29:58]
  wire  _T_2841 = _T_2840 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2842 = iccm_ecc_word_enable[1] & _T_2841; // @[el2_lib.scala 302:32]
  wire  _T_2844 = _T_2842 & _T_2840[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_2459,_T_2844}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 190:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 640:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 192:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 485:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 192:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 192:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 192:72]
  wire  _T_1608 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1613 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1633 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 535:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 401:42]
  wire  _T_1635 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 535:79]
  wire  _T_1636 = _T_1633 | _T_1635; // @[el2_ifu_mem_ctl.scala 535:56]
  wire  _T_1637 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 535:122]
  wire  _T_1638 = ~_T_1637; // @[el2_ifu_mem_ctl.scala 535:101]
  wire  _T_1639 = _T_1636 & _T_1638; // @[el2_ifu_mem_ctl.scala 535:99]
  wire  _T_1640 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1654 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 542:45]
  wire  _T_1655 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 542:69]
  wire  _T_1656 = _T_1654 & _T_1655; // @[el2_ifu_mem_ctl.scala 542:67]
  wire  _T_1657 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_1640 ? _T_1656 : _T_1657; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_1613 ? _T_1639 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_1608 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 192:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 194:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 194:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 284:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 284:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 708:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 275:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 325:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 275:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 275:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 284:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 284:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 284:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 284:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 555:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 597:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 624:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 311:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 605:56]
  wire  _T_1759 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 622:69]
  wire  _T_1760 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 622:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_1759 : _T_1760; // @[el2_ifu_mem_ctl.scala 622:28]
  wire  _T_1706 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 601:68]
  wire  _T_1707 = ic_act_miss_f | _T_1706; // @[el2_ifu_mem_ctl.scala 601:48]
  wire  bus_reset_data_beat_cnt = _T_1707 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 601:91]
  wire  _T_1703 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 600:50]
  wire  _T_1704 = bus_ifu_wr_en_ff & _T_1703; // @[el2_ifu_mem_ctl.scala 600:48]
  wire  _T_1705 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 600:72]
  wire  bus_inc_data_beat_cnt = _T_1704 & _T_1705; // @[el2_ifu_mem_ctl.scala 600:70]
  wire [2:0] _T_1711 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 604:115]
  wire [2:0] _T_1713 = bus_inc_data_beat_cnt ? _T_1711 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_1708 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 602:32]
  wire  _T_1709 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 602:57]
  wire  bus_hold_data_beat_cnt = _T_1708 & _T_1709; // @[el2_ifu_mem_ctl.scala 602:55]
  wire [2:0] _T_1714 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_1713 | _T_1714; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 194:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 195:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 194:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 195:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 201:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 437:45]
  wire  _T_1278 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 458:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 414:60]
  wire  _T_1309 = _T_1278 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1282 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1310 = _T_1282 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1317 = _T_1309 | _T_1310; // @[Mux.scala 27:72]
  wire  _T_1286 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1311 = _T_1286 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1318 = _T_1317 | _T_1311; // @[Mux.scala 27:72]
  wire  _T_1290 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1312 = _T_1290 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1319 = _T_1318 | _T_1312; // @[Mux.scala 27:72]
  wire  _T_1294 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1313 = _T_1294 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1320 = _T_1319 | _T_1313; // @[Mux.scala 27:72]
  wire  _T_1298 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1314 = _T_1298 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1321 = _T_1320 | _T_1314; // @[Mux.scala 27:72]
  wire  _T_1302 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1315 = _T_1302 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1322 = _T_1321 | _T_1315; // @[Mux.scala 27:72]
  wire  _T_1306 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1316 = _T_1306 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_1322 | _T_1316; // @[Mux.scala 27:72]
  wire  _T_1364 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 460:69]
  wire  _T_1365 = ic_miss_buff_data_valid_bypass_index & _T_1364; // @[el2_ifu_mem_ctl.scala 460:67]
  wire  _T_1367 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 460:91]
  wire  _T_1368 = _T_1365 & _T_1367; // @[el2_ifu_mem_ctl.scala 460:89]
  wire  _T_1373 = _T_1365 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 461:65]
  wire  _T_1374 = _T_1368 | _T_1373; // @[el2_ifu_mem_ctl.scala 460:112]
  wire  _T_1376 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 462:43]
  wire  _T_1379 = _T_1376 & _T_1367; // @[el2_ifu_mem_ctl.scala 462:65]
  wire  _T_1380 = _T_1374 | _T_1379; // @[el2_ifu_mem_ctl.scala 461:88]
  wire  _T_1384 = _T_1376 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 463:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 440:75]
  wire  _T_1324 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1348 = _T_1324 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1327 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1349 = _T_1327 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1356 = _T_1348 | _T_1349; // @[Mux.scala 27:72]
  wire  _T_1330 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1350 = _T_1330 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1357 = _T_1356 | _T_1350; // @[Mux.scala 27:72]
  wire  _T_1333 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1351 = _T_1333 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1358 = _T_1357 | _T_1351; // @[Mux.scala 27:72]
  wire  _T_1336 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1352 = _T_1336 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1359 = _T_1358 | _T_1352; // @[Mux.scala 27:72]
  wire  _T_1339 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1353 = _T_1339 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1360 = _T_1359 | _T_1353; // @[Mux.scala 27:72]
  wire  _T_1342 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1354 = _T_1342 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1361 = _T_1360 | _T_1354; // @[Mux.scala 27:72]
  wire  _T_1345 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1355 = _T_1345 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_1361 | _T_1355; // @[Mux.scala 27:72]
  wire  _T_1385 = _T_1384 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 463:87]
  wire  _T_1386 = _T_1380 | _T_1385; // @[el2_ifu_mem_ctl.scala 462:88]
  wire  _T_1390 = ic_miss_buff_data_valid_bypass_index & _T_1306; // @[el2_ifu_mem_ctl.scala 464:43]
  wire  miss_buff_hit_unq_f = _T_1386 | _T_1390; // @[el2_ifu_mem_ctl.scala 463:131]
  wire  _T_1406 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 469:55]
  wire  _T_1407 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 469:87]
  wire  _T_1408 = _T_1406 | _T_1407; // @[el2_ifu_mem_ctl.scala 469:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_1408; // @[el2_ifu_mem_ctl.scala 469:41]
  wire  _T_1391 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 466:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 312:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 457:51]
  wire  _T_1392 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 466:68]
  wire  _T_1393 = miss_buff_hit_unq_f & _T_1392; // @[el2_ifu_mem_ctl.scala 466:66]
  wire  stream_hit_f = _T_1391 & _T_1393; // @[el2_ifu_mem_ctl.scala 466:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 279:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 279:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 607:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 634:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 205:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 205:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 205:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 205:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 207:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 208:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 209:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 209:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 209:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 197:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 209:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 209:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 210:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 210:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 210:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 210:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 211:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 212:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 209:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 208:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 207:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 206:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_1403 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 468:60]
  wire  _T_1404 = _T_1403 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 468:92]
  wire  stream_eol_f = _T_1404 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 468:110]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 220:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 220:87]
  wire  _T_113 = _T_111 & _T_1705; // @[el2_ifu_mem_ctl.scala 220:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 220:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 224:48]
  wire  _T_126 = _T_124 & _T_1705; // @[el2_ifu_mem_ctl.scala 224:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 285:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 285:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 285:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 285:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 285:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 285:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 286:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 339:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 286:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 286:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 286:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:50]
  wire  _T_137 = _T_135 & _T_1705; // @[el2_ifu_mem_ctl.scala 228:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 287:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 288:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 288:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 287:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:35]
  wire  _T_143 = _T_141 & _T_1705; // @[el2_ifu_mem_ctl.scala 229:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 234:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 233:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 238:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 238:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 195:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 195:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 195:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 195:91]
  wire  _T_30 = ic_act_miss_f & _T_1705; // @[el2_ifu_mem_ctl.scala 202:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 213:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 213:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 213:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 213:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 217:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 217:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 221:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 225:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 230:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 235:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 235:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 255:95]
  wire  _T_175 = _T_1406 & _T_174; // @[el2_ifu_mem_ctl.scala 255:93]
  wire  crit_wd_byp_ok_ff = _T_1407 | _T_175; // @[el2_ifu_mem_ctl.scala 255:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 256:36]
  wire  _T_180 = _T_1406 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 256:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 256:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 256:70]
  wire  _T_184 = _T_1406 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 257:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 257:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 256:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 257:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 258:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 258:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 257:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 260:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:35]
  reg [6:0] _T_4284; // @[el2_ifu_mem_ctl.scala 736:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_4284[5:0]; // @[el2_ifu_mem_ctl.scala 735:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 732:121]
  wire  _T_4149 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4151 = _T_4149 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3640; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_3640[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4152 = _T_4151 & _GEN_473; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4145 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4147 = _T_4145 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3636; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_3636[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4148 = _T_4147 & _GEN_475; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4141 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4143 = _T_4141 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3632; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_3632[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4144 = _T_4143 & _GEN_477; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4137 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4139 = _T_4137 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3628; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_3628[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4140 = _T_4139 & _GEN_479; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4133 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4135 = _T_4133 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3624; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_3624[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4136 = _T_4135 & _GEN_481; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4129 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4131 = _T_4129 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3620; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_3620[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4132 = _T_4131 & _GEN_483; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4125 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4127 = _T_4125 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3616; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_3616[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4128 = _T_4127 & _GEN_485; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4121 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4123 = _T_4121 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3612; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_3612[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4124 = _T_4123 & _GEN_487; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4117 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4119 = _T_4117 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3608; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_3608[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4120 = _T_4119 & _GEN_489; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4113 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4115 = _T_4113 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3604; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_3604[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4116 = _T_4115 & _GEN_491; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [59:0] _T_4161 = {_T_4152,_T_4148,_T_4144,_T_4140,_T_4136,_T_4132,_T_4128,_T_4124,_T_4120,_T_4116}; // @[Cat.scala 29:58]
  wire  _T_4109 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4111 = _T_4109 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3600; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_3600[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4112 = _T_4111 & _GEN_493; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4105 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4107 = _T_4105 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3596; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_3596[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4108 = _T_4107 & _GEN_495; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4101 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4103 = _T_4101 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3592; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_3592[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4104 = _T_4103 & _GEN_497; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4097 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4099 = _T_4097 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3588; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_3588[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4100 = _T_4099 & _GEN_499; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4093 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4095 = _T_4093 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3584; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_3584[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4096 = _T_4095 & _GEN_501; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4089 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4091 = _T_4089 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3580; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_3580[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4092 = _T_4091 & _GEN_503; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4085 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4087 = _T_4085 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3576; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_3576[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4088 = _T_4087 & _GEN_505; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4081 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4083 = _T_4081 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3572; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_3572[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4084 = _T_4083 & _GEN_507; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4077 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4079 = _T_4077 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3568; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_3568[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4080 = _T_4079 & _GEN_509; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [113:0] _T_4170 = {_T_4161,_T_4112,_T_4108,_T_4104,_T_4100,_T_4096,_T_4092,_T_4088,_T_4084,_T_4080}; // @[Cat.scala 29:58]
  wire  _T_4073 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4075 = _T_4073 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3564; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_3564[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4076 = _T_4075 & _GEN_511; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4069 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4071 = _T_4069 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3560; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_3560[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4072 = _T_4071 & _GEN_513; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4065 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4067 = _T_4065 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3556; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_3556[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4068 = _T_4067 & _GEN_515; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4061 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4063 = _T_4061 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3552; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_3552[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4064 = _T_4063 & _GEN_517; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4057 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4059 = _T_4057 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3548; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_3548[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4060 = _T_4059 & _GEN_519; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4053 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4055 = _T_4053 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3544; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_3544[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4056 = _T_4055 & _GEN_521; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4049 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4051 = _T_4049 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3540; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_3540[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4052 = _T_4051 & _GEN_523; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4045 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4047 = _T_4045 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3536; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_3536[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4048 = _T_4047 & _GEN_525; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4041 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4043 = _T_4041 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3532; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_3532[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4044 = _T_4043 & _GEN_527; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [167:0] _T_4179 = {_T_4170,_T_4076,_T_4072,_T_4068,_T_4064,_T_4060,_T_4056,_T_4052,_T_4048,_T_4044}; // @[Cat.scala 29:58]
  wire  _T_4037 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4039 = _T_4037 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3528; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_3528[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4040 = _T_4039 & _GEN_529; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4033 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4035 = _T_4033 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3524; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_3524[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4036 = _T_4035 & _GEN_531; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4029 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4031 = _T_4029 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3520; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_3520[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4032 = _T_4031 & _GEN_533; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4025 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4027 = _T_4025 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3516; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_3516[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4028 = _T_4027 & _GEN_535; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4021 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4023 = _T_4021 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3512; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_3512[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4024 = _T_4023 & _GEN_537; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4017 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4019 = _T_4017 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3508; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_3508[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4020 = _T_4019 & _GEN_539; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4013 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4015 = _T_4013 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3504; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_3504[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4016 = _T_4015 & _GEN_541; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4009 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4011 = _T_4009 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3500; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_3500[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4012 = _T_4011 & _GEN_543; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4005 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4007 = _T_4005 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3496; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_3496[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4008 = _T_4007 & _GEN_545; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [221:0] _T_4188 = {_T_4179,_T_4040,_T_4036,_T_4032,_T_4028,_T_4024,_T_4020,_T_4016,_T_4012,_T_4008}; // @[Cat.scala 29:58]
  wire  _T_4001 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4003 = _T_4001 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3492; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_3492[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4004 = _T_4003 & _GEN_547; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3997 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3999 = _T_3997 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3488; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_3488[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4000 = _T_3999 & _GEN_549; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3993 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3995 = _T_3993 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3484; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_3484[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3996 = _T_3995 & _GEN_551; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3989 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3991 = _T_3989 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3480; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_3480[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3992 = _T_3991 & _GEN_553; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3985 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3987 = _T_3985 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3476; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_3476[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3988 = _T_3987 & _GEN_555; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3981 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3983 = _T_3981 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3472; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_3472[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3984 = _T_3983 & _GEN_557; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3977 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3979 = _T_3977 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3468; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_3468[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3980 = _T_3979 & _GEN_559; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3973 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3975 = _T_3973 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3464; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_3464[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3976 = _T_3975 & _GEN_561; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3969 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3971 = _T_3969 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3460; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_3460[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3972 = _T_3971 & _GEN_563; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [275:0] _T_4197 = {_T_4188,_T_4004,_T_4000,_T_3996,_T_3992,_T_3988,_T_3984,_T_3980,_T_3976,_T_3972}; // @[Cat.scala 29:58]
  wire  _T_3965 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3967 = _T_3965 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3456; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_3456[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3968 = _T_3967 & _GEN_565; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3961 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3963 = _T_3961 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3452; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_3452[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3964 = _T_3963 & _GEN_567; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3957 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3959 = _T_3957 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3448; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_3448[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3960 = _T_3959 & _GEN_569; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3953 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3955 = _T_3953 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3444; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_3444[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3956 = _T_3955 & _GEN_571; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3949 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3951 = _T_3949 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3440; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_3440[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3952 = _T_3951 & _GEN_573; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3945 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3947 = _T_3945 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3436; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_3436[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3948 = _T_3947 & _GEN_575; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3941 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3943 = _T_3941 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3432; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_3432[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3944 = _T_3943 & _GEN_577; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3937 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3939 = _T_3937 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3428; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_3428[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3940 = _T_3939 & _GEN_579; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3933 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3935 = _T_3933 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3424; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_3424[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3936 = _T_3935 & _GEN_581; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [329:0] _T_4206 = {_T_4197,_T_3968,_T_3964,_T_3960,_T_3956,_T_3952,_T_3948,_T_3944,_T_3940,_T_3936}; // @[Cat.scala 29:58]
  wire  _T_3929 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3931 = _T_3929 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3420; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_3420[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3932 = _T_3931 & _GEN_583; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3925 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3927 = _T_3925 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3416; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_3416[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3928 = _T_3927 & _GEN_585; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3921 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3923 = _T_3921 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3412; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_3412[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3924 = _T_3923 & _GEN_587; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3917 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3919 = _T_3917 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3408; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_3408[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3920 = _T_3919 & _GEN_589; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3913 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3915 = _T_3913 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3404; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_3404[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3916 = _T_3915 & _GEN_591; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3909 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3911 = _T_3909 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3400; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_3400[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3912 = _T_3911 & _GEN_593; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3905 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3907 = _T_3905 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3396; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_3396[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3908 = _T_3907 & _GEN_595; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3901 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3903 = _T_3901 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3392; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_3392[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3904 = _T_3903 & _GEN_597; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3897 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3899 = _T_3897 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3388; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_3388[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3900 = _T_3899 & _GEN_599; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [383:0] _T_4215 = {_T_4206,_T_3932,_T_3928,_T_3924,_T_3920,_T_3916,_T_3912,_T_3908,_T_3904,_T_3900}; // @[Cat.scala 29:58]
  wire  _T_3893 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3895 = _T_3893 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3384; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_3384[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3896 = _T_3895 & _GEN_600; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3889 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3891 = _T_3889 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3380; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_3380[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3892 = _T_3891 & _GEN_601; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3885 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3887 = _T_3885 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3376; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_3376[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3888 = _T_3887 & _GEN_602; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3881 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3883 = _T_3881 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3372; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_3372[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3884 = _T_3883 & _GEN_603; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3877 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3879 = _T_3877 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3368; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_3368[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3880 = _T_3879 & _GEN_604; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3873 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3875 = _T_3873 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3364; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_3364[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3876 = _T_3875 & _GEN_605; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3869 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3871 = _T_3869 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3360; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_3360[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3872 = _T_3871 & _GEN_606; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3865 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3867 = _T_3865 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3356; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_3356[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3868 = _T_3867 & _GEN_607; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3861 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3863 = _T_3861 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3352; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_3352[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3864 = _T_3863 & _GEN_608; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [437:0] _T_4224 = {_T_4215,_T_3896,_T_3892,_T_3888,_T_3884,_T_3880,_T_3876,_T_3872,_T_3868,_T_3864}; // @[Cat.scala 29:58]
  wire  _T_3857 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3859 = _T_3857 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3348; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_3348[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3860 = _T_3859 & _GEN_609; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3853 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3855 = _T_3853 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3344; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_3344[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3856 = _T_3855 & _GEN_610; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3849 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3851 = _T_3849 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3340; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_3340[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3852 = _T_3851 & _GEN_611; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3845 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3847 = _T_3845 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3336; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_3336[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3848 = _T_3847 & _GEN_612; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3841 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3843 = _T_3841 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3332; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_3332[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3844 = _T_3843 & _GEN_613; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3837 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3839 = _T_3837 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3328; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_3328[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3840 = _T_3839 & _GEN_614; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3833 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3835 = _T_3833 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3324; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_3324[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3836 = _T_3835 & _GEN_615; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3829 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3831 = _T_3829 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3320; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_3320[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3832 = _T_3831 & _GEN_616; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3825 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3827 = _T_3825 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3316; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_3316[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3828 = _T_3827 & _GEN_617; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [491:0] _T_4233 = {_T_4224,_T_3860,_T_3856,_T_3852,_T_3848,_T_3844,_T_3840,_T_3836,_T_3832,_T_3828}; // @[Cat.scala 29:58]
  wire  _T_3821 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3823 = _T_3821 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3312; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_3312[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3824 = _T_3823 & _GEN_618; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3817 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3819 = _T_3817 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3308; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_3308[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3820 = _T_3819 & _GEN_619; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3813 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3815 = _T_3813 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3304; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_3304[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3816 = _T_3815 & _GEN_620; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3809 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3811 = _T_3809 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3300; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_3300[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3812 = _T_3811 & _GEN_621; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3805 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3807 = _T_3805 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3296; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_3296[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3808 = _T_3807 & _GEN_622; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3801 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3803 = _T_3801 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3292; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_3292[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3804 = _T_3803 & _GEN_623; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3797 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3799 = _T_3797 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3288; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_3288[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3800 = _T_3799 & _GEN_624; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3793 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3795 = _T_3793 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3284; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_3284[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3796 = _T_3795 & _GEN_625; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3789 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3791 = _T_3789 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3280; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_3280[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3792 = _T_3791 & _GEN_626; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [545:0] _T_4242 = {_T_4233,_T_3824,_T_3820,_T_3816,_T_3812,_T_3808,_T_3804,_T_3800,_T_3796,_T_3792}; // @[Cat.scala 29:58]
  wire  _T_3785 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3787 = _T_3785 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3276; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_3276[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3788 = _T_3787 & _GEN_627; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3781 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3783 = _T_3781 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3272; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_3272[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3784 = _T_3783 & _GEN_628; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3777 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3779 = _T_3777 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3268; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_3268[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3780 = _T_3779 & _GEN_629; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3773 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3775 = _T_3773 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3264; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_3264[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3776 = _T_3775 & _GEN_630; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3769 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3771 = _T_3769 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3260; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_3260[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3772 = _T_3771 & _GEN_631; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3765 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3767 = _T_3765 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3256; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_3256[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3768 = _T_3767 & _GEN_632; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3761 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3763 = _T_3761 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3252; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_3252[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3764 = _T_3763 & _GEN_633; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3757 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3759 = _T_3757 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3248; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_3248[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3760 = _T_3759 & _GEN_634; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3753 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3755 = _T_3753 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3244; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_3244[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3756 = _T_3755 & _GEN_635; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [599:0] _T_4251 = {_T_4242,_T_3788,_T_3784,_T_3780,_T_3776,_T_3772,_T_3768,_T_3764,_T_3760,_T_3756}; // @[Cat.scala 29:58]
  wire  _T_3749 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3751 = _T_3749 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3240; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_3240[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3752 = _T_3751 & _GEN_636; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3745 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3747 = _T_3745 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3236; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_3236[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3748 = _T_3747 & _GEN_637; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3741 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3743 = _T_3741 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3232; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_3232[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3744 = _T_3743 & _GEN_638; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3737 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3739 = _T_3737 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3228; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_3228[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3740 = _T_3739 & _GEN_639; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3733 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3735 = _T_3733 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3224; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_3224[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3736 = _T_3735 & _GEN_640; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3729 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3731 = _T_3729 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3220; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_3220[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3732 = _T_3731 & _GEN_641; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3725 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3727 = _T_3725 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3216; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_3216[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3728 = _T_3727 & _GEN_642; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3721 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3723 = _T_3721 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3212; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_3212[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3724 = _T_3723 & _GEN_643; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3717 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3719 = _T_3717 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3208; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_3208[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3720 = _T_3719 & _GEN_644; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [653:0] _T_4260 = {_T_4251,_T_3752,_T_3748,_T_3744,_T_3740,_T_3736,_T_3732,_T_3728,_T_3724,_T_3720}; // @[Cat.scala 29:58]
  wire  _T_3713 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3715 = _T_3713 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3204; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_3204[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3716 = _T_3715 & _GEN_645; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3709 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3711 = _T_3709 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3200; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_3200[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3712 = _T_3711 & _GEN_646; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3705 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3707 = _T_3705 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3196; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_3196[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3708 = _T_3707 & _GEN_647; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3701 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3703 = _T_3701 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3192; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_3192[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3704 = _T_3703 & _GEN_648; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3697 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3699 = _T_3697 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3188; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_3188[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3700 = _T_3699 & _GEN_649; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3693 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3695 = _T_3693 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3184; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_3184[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3696 = _T_3695 & _GEN_650; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3689 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3691 = _T_3689 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3180; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_3180[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3692 = _T_3691 & _GEN_651; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3685 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3687 = _T_3685 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3176; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_3176[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3688 = _T_3687 & _GEN_652; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3681 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3683 = _T_3681 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3172; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_3172[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3684 = _T_3683 & _GEN_653; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [707:0] _T_4269 = {_T_4260,_T_3716,_T_3712,_T_3708,_T_3704,_T_3700,_T_3696,_T_3692,_T_3688,_T_3684}; // @[Cat.scala 29:58]
  wire  _T_3677 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3679 = _T_3677 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3168; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3168[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3680 = _T_3679 & _GEN_654; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3673 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3675 = _T_3673 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3164; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3164[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3676 = _T_3675 & _GEN_655; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3669 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3671 = _T_3669 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3160; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3160[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3672 = _T_3671 & _GEN_656; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3665 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3667 = _T_3665 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3156; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3156[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3668 = _T_3667 & _GEN_657; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3661 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3663 = _T_3661 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3152; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3152[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3664 = _T_3663 & _GEN_658; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3657 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3659 = _T_3657 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3148; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3148[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3660 = _T_3659 & _GEN_659; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3653 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3655 = _T_3653 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3144; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3144[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3656 = _T_3655 & _GEN_660; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3649 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3651 = _T_3649 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3140; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3140[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3652 = _T_3651 & _GEN_661; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3645 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3647 = _T_3645 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3136; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3136[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3648 = _T_3647 & _GEN_662; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [761:0] _T_4278 = {_T_4269,_T_3680,_T_3676,_T_3672,_T_3668,_T_3664,_T_3660,_T_3656,_T_3652,_T_3648}; // @[Cat.scala 29:58]
  wire  _T_3641 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3643 = _T_3641 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3132; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3132[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3644 = _T_3643 & _GEN_663; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [767:0] _T_4279 = {_T_4278,_T_3644}; // @[Cat.scala 29:58]
  wire  way_status = _T_4279[0]; // @[el2_ifu_mem_ctl.scala 732:16]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 263:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 265:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 272:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 277:59]
  wire  _T_214 = _T_212 | _T_1391; // @[el2_ifu_mem_ctl.scala 277:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 277:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 283:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 283:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 283:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 290:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 290:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 290:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 291:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 291:32]
  wire  _T_274 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 294:75]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 294:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_1780 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 630:48]
  wire  _T_1781 = _T_1780 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 630:52]
  wire  bus_ifu_wr_data_error_ff = _T_1781 & miss_pending; // @[el2_ifu_mem_ctl.scala 630:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 376:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 375:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 294:145]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 294:143]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 297:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 298:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 317:30]
  wire  _T_9229 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 785:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 318:24]
  wire  _T_9231 = _T_9229 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 785:51]
  wire  _T_9233 = _T_9231 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 785:67]
  wire  _T_9235 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 785:86]
  wire  replace_way_mb_any_0 = _T_9233 | _T_9235; // @[el2_ifu_mem_ctl.scala 785:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9238 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:50]
  wire  _T_9240 = _T_9238 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:66]
  wire  _T_9242 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:85]
  wire  _T_9244 = _T_9242 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:100]
  wire  replace_way_mb_any_1 = _T_9240 | _T_9244; // @[el2_ifu_mem_ctl.scala 786:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 302:110]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 306:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 306:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 307:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 306:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 308:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 316:23]
  wire  _T_313 = _T_1406 & flush_final_f; // @[el2_ifu_mem_ctl.scala 320:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 320:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 320:53]
  wire  _T_1398 = ~_T_1393; // @[el2_ifu_mem_ctl.scala 467:46]
  wire  _T_1399 = _T_1391 & _T_1398; // @[el2_ifu_mem_ctl.scala 467:44]
  wire  stream_miss_f = _T_1399 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 467:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 320:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 320:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 326:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_1391; // @[el2_ifu_mem_ctl.scala 328:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 328:82]
  wire  _T_1412 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 472:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_1412}; // @[Cat.scala 29:58]
  wire  _T_1413 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1437 = _T_1413 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1416 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1438 = _T_1416 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1437 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1419 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1439 = _T_1419 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1422 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1440 = _T_1422 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1425 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1441 = _T_1425 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1428 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1442 = _T_1428 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1431 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1443 = _T_1431 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1450 = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1434 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1444 = _T_1434 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_1450 | _T_1444; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 474:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 332:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 332:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 627:61]
  wire  _T_1774 = ic_act_miss_f_delayed & _T_1407; // @[el2_ifu_mem_ctl.scala 628:53]
  wire  reset_tag_valid_for_miss = _T_1774 & _T_17; // @[el2_ifu_mem_ctl.scala 628:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 332:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 334:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 336:84]
  wire  _T_1768 = ~_T_1780; // @[el2_ifu_mem_ctl.scala 625:84]
  wire  _T_1769 = _T_100 & _T_1768; // @[el2_ifu_mem_ctl.scala 625:82]
  wire  bus_ifu_wr_en_ff_q = _T_1769 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 625:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 336:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 337:31]
  wire [6:0] ic_wr_ecc = m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 346:13]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] ic_miss_buff_ecc = m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 350:20]
  wire [3:0] _T_1453 = {ifu_bus_rid_ff[2:1],_T_1412,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1454 = _T_1453 == 4'h0; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_1501 = _T_1454 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1457 = _T_1453 == 4'h1; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_1502 = _T_1457 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1517 = _T_1501 | _T_1502; // @[Mux.scala 27:72]
  wire  _T_1460 = _T_1453 == 4'h2; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_1503 = _T_1460 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1518 = _T_1517 | _T_1503; // @[Mux.scala 27:72]
  wire  _T_1463 = _T_1453 == 4'h3; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_1504 = _T_1463 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1519 = _T_1518 | _T_1504; // @[Mux.scala 27:72]
  wire  _T_1466 = _T_1453 == 4'h4; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_1505 = _T_1466 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1520 = _T_1519 | _T_1505; // @[Mux.scala 27:72]
  wire  _T_1469 = _T_1453 == 4'h5; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_1506 = _T_1469 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1521 = _T_1520 | _T_1506; // @[Mux.scala 27:72]
  wire  _T_1472 = _T_1453 == 4'h6; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_1507 = _T_1472 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1522 = _T_1521 | _T_1507; // @[Mux.scala 27:72]
  wire  _T_1475 = _T_1453 == 4'h7; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_1508 = _T_1475 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1523 = _T_1522 | _T_1508; // @[Mux.scala 27:72]
  wire  _T_1478 = _T_1453 == 4'h8; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_1509 = _T_1478 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1524 = _T_1523 | _T_1509; // @[Mux.scala 27:72]
  wire  _T_1481 = _T_1453 == 4'h9; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_1510 = _T_1481 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1525 = _T_1524 | _T_1510; // @[Mux.scala 27:72]
  wire  _T_1484 = _T_1453 == 4'ha; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_1511 = _T_1484 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1526 = _T_1525 | _T_1511; // @[Mux.scala 27:72]
  wire  _T_1487 = _T_1453 == 4'hb; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_1512 = _T_1487 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1527 = _T_1526 | _T_1512; // @[Mux.scala 27:72]
  wire  _T_1490 = _T_1453 == 4'hc; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_1513 = _T_1490 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1528 = _T_1527 | _T_1513; // @[Mux.scala 27:72]
  wire  _T_1493 = _T_1453 == 4'hd; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_1514 = _T_1493 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1529 = _T_1528 | _T_1514; // @[Mux.scala 27:72]
  wire  _T_1496 = _T_1453 == 4'he; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_1515 = _T_1496 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1530 = _T_1529 | _T_1515; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1453 == 4'hf; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_1516 = _T_1499 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1531 = _T_1530 | _T_1516; // @[Mux.scala 27:72]
  wire [3:0] _T_1533 = {ifu_bus_rid_ff[2:1],_T_1412,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1534 = _T_1533 == 4'h0; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1557 = _T_1534 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1537 = _T_1533 == 4'h1; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1558 = _T_1537 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1565 = _T_1557 | _T_1558; // @[Mux.scala 27:72]
  wire  _T_1540 = _T_1533 == 4'h2; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1559 = _T_1540 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1566 = _T_1565 | _T_1559; // @[Mux.scala 27:72]
  wire  _T_1543 = _T_1533 == 4'h3; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1560 = _T_1543 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1567 = _T_1566 | _T_1560; // @[Mux.scala 27:72]
  wire  _T_1546 = _T_1533 == 4'h4; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1561 = _T_1546 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1568 = _T_1567 | _T_1561; // @[Mux.scala 27:72]
  wire  _T_1549 = _T_1533 == 4'h5; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1562 = _T_1549 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1569 = _T_1568 | _T_1562; // @[Mux.scala 27:72]
  wire  _T_1552 = _T_1533 == 4'h6; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1563 = _T_1552 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1570 = _T_1569 | _T_1563; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1533 == 4'h7; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1564 = _T_1555 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1571 = _T_1570 | _T_1564; // @[Mux.scala 27:72]
  wire [141:0] _T_392 = {ic_wr_ecc,ifu_bus_rdata_ff,ic_miss_buff_ecc,_T_1531,_T_1571}; // @[Cat.scala 29:58]
  wire [141:0] _T_395 = {ic_miss_buff_ecc,_T_1531,_T_1571,ic_wr_ecc,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_392 : _T_395; // @[el2_ifu_mem_ctl.scala 366:28]
  wire  _T_352 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 356:56]
  wire  _T_353 = _T_352 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 356:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 422:28]
  wire  _T_571 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 623:35]
  wire  _T_440 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_440; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_497 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 413:118]
  wire  _T_498 = ic_miss_buff_data_valid[0] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_498; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_594 = _T_571 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_574 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_441 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_441; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_501 = ic_miss_buff_data_valid[1] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_501; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_595 = _T_574 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_602 = _T_594 | _T_595; // @[Mux.scala 27:72]
  wire  _T_577 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_442 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_442; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_504 = ic_miss_buff_data_valid[2] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_504; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_596 = _T_577 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_603 = _T_602 | _T_596; // @[Mux.scala 27:72]
  wire  _T_580 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_443 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_443; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_507 = ic_miss_buff_data_valid[3] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_507; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_597 = _T_580 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_604 = _T_603 | _T_597; // @[Mux.scala 27:72]
  wire  _T_583 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_444 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_444; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_510 = ic_miss_buff_data_valid[4] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_510; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_598 = _T_583 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_605 = _T_604 | _T_598; // @[Mux.scala 27:72]
  wire  _T_586 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_445 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_445; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_513 = ic_miss_buff_data_valid[5] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_513; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_599 = _T_586 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_606 = _T_605 | _T_599; // @[Mux.scala 27:72]
  wire  _T_589 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_446 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_446; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_516 = ic_miss_buff_data_valid[6] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_516; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_600 = _T_589 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_607 = _T_606 | _T_600; // @[Mux.scala 27:72]
  wire  _T_592 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_447 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_447; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_519 = ic_miss_buff_data_valid[7] & _T_497; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_519; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_601 = _T_592 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_607 | _T_601; // @[Mux.scala 27:72]
  wire  _T_610 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 425:58]
  wire  _T_611 = bypass_valid_value_check & _T_610; // @[el2_ifu_mem_ctl.scala 425:56]
  wire  _T_613 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 425:77]
  wire  _T_614 = _T_611 & _T_613; // @[el2_ifu_mem_ctl.scala 425:75]
  wire  _T_619 = _T_611 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 426:75]
  wire  _T_620 = _T_614 | _T_619; // @[el2_ifu_mem_ctl.scala 425:95]
  wire  _T_622 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 427:56]
  wire  _T_625 = _T_622 & _T_613; // @[el2_ifu_mem_ctl.scala 427:74]
  wire  _T_626 = _T_620 | _T_625; // @[el2_ifu_mem_ctl.scala 426:94]
  wire  _T_630 = _T_622 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 428:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 423:70]
  wire  _T_631 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_647 = _T_631 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_633 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_648 = _T_633 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_655 = _T_647 | _T_648; // @[Mux.scala 27:72]
  wire  _T_635 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_649 = _T_635 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_656 = _T_655 | _T_649; // @[Mux.scala 27:72]
  wire  _T_637 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_650 = _T_637 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_657 = _T_656 | _T_650; // @[Mux.scala 27:72]
  wire  _T_639 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_651 = _T_639 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_658 = _T_657 | _T_651; // @[Mux.scala 27:72]
  wire  _T_641 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_652 = _T_641 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_659 = _T_658 | _T_652; // @[Mux.scala 27:72]
  wire  _T_643 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_653 = _T_643 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_660 = _T_659 | _T_653; // @[Mux.scala 27:72]
  wire  _T_645 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_654 = _T_645 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_661 = _T_660 | _T_654; // @[Mux.scala 27:72]
  wire  _T_663 = _T_630 & _T_661; // @[el2_ifu_mem_ctl.scala 428:69]
  wire  _T_664 = _T_626 | _T_663; // @[el2_ifu_mem_ctl.scala 427:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 429:95]
  wire  _T_667 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 429:95]
  wire  _T_668 = bypass_valid_value_check & _T_667; // @[el2_ifu_mem_ctl.scala 429:56]
  wire  bypass_data_ready_in = _T_664 | _T_668; // @[el2_ifu_mem_ctl.scala 428:181]
  wire  _T_669 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 433:53]
  wire  _T_670 = _T_669 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 433:73]
  wire  _T_672 = _T_670 & _T_317; // @[el2_ifu_mem_ctl.scala 433:96]
  wire  _T_674 = _T_672 & _T_58; // @[el2_ifu_mem_ctl.scala 433:118]
  wire  _T_676 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 434:73]
  wire  _T_678 = _T_676 & _T_317; // @[el2_ifu_mem_ctl.scala 434:96]
  wire  _T_680 = _T_678 & _T_58; // @[el2_ifu_mem_ctl.scala 434:118]
  wire  _T_681 = _T_674 | _T_680; // @[el2_ifu_mem_ctl.scala 433:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 436:58]
  wire  _T_682 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 435:54]
  wire  _T_683 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 435:76]
  wire  _T_684 = _T_682 & _T_683; // @[el2_ifu_mem_ctl.scala 435:74]
  wire  _T_686 = _T_684 & _T_317; // @[el2_ifu_mem_ctl.scala 435:96]
  wire  ic_crit_wd_rdy_new_in = _T_681 | _T_686; // @[el2_ifu_mem_ctl.scala 434:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 633:43]
  wire  _T_407 = ic_crit_wd_rdy | _T_1391; // @[el2_ifu_mem_ctl.scala 380:38]
  wire  _T_409 = _T_407 | _T_1407; // @[el2_ifu_mem_ctl.scala 380:64]
  wire  _T_410 = ~_T_409; // @[el2_ifu_mem_ctl.scala 380:21]
  wire  _T_411 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 380:98]
  wire  sel_ic_data = _T_410 & _T_411; // @[el2_ifu_mem_ctl.scala 380:96]
  wire  _T_1574 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 478:44]
  wire  _T_780 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 447:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 419:60]
  wire  _T_724 = _T_571 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_725 = _T_574 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_732 = _T_724 | _T_725; // @[Mux.scala 27:72]
  wire  _T_726 = _T_577 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_733 = _T_732 | _T_726; // @[Mux.scala 27:72]
  wire  _T_727 = _T_580 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_734 = _T_733 | _T_727; // @[Mux.scala 27:72]
  wire  _T_728 = _T_583 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_735 = _T_734 | _T_728; // @[Mux.scala 27:72]
  wire  _T_729 = _T_586 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_736 = _T_735 | _T_729; // @[Mux.scala 27:72]
  wire  _T_730 = _T_589 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_737 = _T_736 | _T_730; // @[Mux.scala 27:72]
  wire  _T_731 = _T_592 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_737 | _T_731; // @[Mux.scala 27:72]
  wire  _T_763 = _T_1324 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_764 = _T_1327 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_771 = _T_763 | _T_764; // @[Mux.scala 27:72]
  wire  _T_765 = _T_1330 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_772 = _T_771 | _T_765; // @[Mux.scala 27:72]
  wire  _T_766 = _T_1333 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_773 = _T_772 | _T_766; // @[Mux.scala 27:72]
  wire  _T_767 = _T_1336 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_774 = _T_773 | _T_767; // @[Mux.scala 27:72]
  wire  _T_768 = _T_1339 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_775 = _T_774 | _T_768; // @[Mux.scala 27:72]
  wire  _T_769 = _T_1342 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_776 = _T_775 | _T_769; // @[Mux.scala 27:72]
  wire  _T_770 = _T_1345 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_776 | _T_770; // @[Mux.scala 27:72]
  wire  _T_781 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 449:70]
  wire  ifu_byp_data_err_new = _T_780 ? ic_miss_buff_data_error_bypass : _T_781; // @[el2_ifu_mem_ctl.scala 447:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 391:42]
  wire  _T_1575 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 478:91]
  wire  _T_1576 = ~_T_1575; // @[el2_ifu_mem_ctl.scala 478:60]
  wire  ic_rd_parity_final_err = _T_1574 & _T_1576; // @[el2_ifu_mem_ctl.scala 478:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_8847 = _T_3641 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 760:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_8849 = _T_3645 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9102 = _T_8847 | _T_8849; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_8851 = _T_3649 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9103 = _T_9102 | _T_8851; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_8853 = _T_3653 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9104 = _T_9103 | _T_8853; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_8855 = _T_3657 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9105 = _T_9104 | _T_8855; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_8857 = _T_3661 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9106 = _T_9105 | _T_8857; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_8859 = _T_3665 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9107 = _T_9106 | _T_8859; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_8861 = _T_3669 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9108 = _T_9107 | _T_8861; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_8863 = _T_3673 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9109 = _T_9108 | _T_8863; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_8865 = _T_3677 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9110 = _T_9109 | _T_8865; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_8867 = _T_3681 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9111 = _T_9110 | _T_8867; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_8869 = _T_3685 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9112 = _T_9111 | _T_8869; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_8871 = _T_3689 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9113 = _T_9112 | _T_8871; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_8873 = _T_3693 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9114 = _T_9113 | _T_8873; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_8875 = _T_3697 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9115 = _T_9114 | _T_8875; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_8877 = _T_3701 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9116 = _T_9115 | _T_8877; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_8879 = _T_3705 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9117 = _T_9116 | _T_8879; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_8881 = _T_3709 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9118 = _T_9117 | _T_8881; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_8883 = _T_3713 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9119 = _T_9118 | _T_8883; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_8885 = _T_3717 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9120 = _T_9119 | _T_8885; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_8887 = _T_3721 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9121 = _T_9120 | _T_8887; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_8889 = _T_3725 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9122 = _T_9121 | _T_8889; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_8891 = _T_3729 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9123 = _T_9122 | _T_8891; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_8893 = _T_3733 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9124 = _T_9123 | _T_8893; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_8895 = _T_3737 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9125 = _T_9124 | _T_8895; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_8897 = _T_3741 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9126 = _T_9125 | _T_8897; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_8899 = _T_3745 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9127 = _T_9126 | _T_8899; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_8901 = _T_3749 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9128 = _T_9127 | _T_8901; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_8903 = _T_3753 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9129 = _T_9128 | _T_8903; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_8905 = _T_3757 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9130 = _T_9129 | _T_8905; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_8907 = _T_3761 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9131 = _T_9130 | _T_8907; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_8909 = _T_3765 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9132 = _T_9131 | _T_8909; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_8911 = _T_3769 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9133 = _T_9132 | _T_8911; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_8913 = _T_3773 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9134 = _T_9133 | _T_8913; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_8915 = _T_3777 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9135 = _T_9134 | _T_8915; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_8917 = _T_3781 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9136 = _T_9135 | _T_8917; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_8919 = _T_3785 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9137 = _T_9136 | _T_8919; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_8921 = _T_3789 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9138 = _T_9137 | _T_8921; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_8923 = _T_3793 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9139 = _T_9138 | _T_8923; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_8925 = _T_3797 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9140 = _T_9139 | _T_8925; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_8927 = _T_3801 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9141 = _T_9140 | _T_8927; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_8929 = _T_3805 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9142 = _T_9141 | _T_8929; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_8931 = _T_3809 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9143 = _T_9142 | _T_8931; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_8933 = _T_3813 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9144 = _T_9143 | _T_8933; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_8935 = _T_3817 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9145 = _T_9144 | _T_8935; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_8937 = _T_3821 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9146 = _T_9145 | _T_8937; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_8939 = _T_3825 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9147 = _T_9146 | _T_8939; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_8941 = _T_3829 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9148 = _T_9147 | _T_8941; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_8943 = _T_3833 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9149 = _T_9148 | _T_8943; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_8945 = _T_3837 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9150 = _T_9149 | _T_8945; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_8947 = _T_3841 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9151 = _T_9150 | _T_8947; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_8949 = _T_3845 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9152 = _T_9151 | _T_8949; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_8951 = _T_3849 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9153 = _T_9152 | _T_8951; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_8953 = _T_3853 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9154 = _T_9153 | _T_8953; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_8955 = _T_3857 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9155 = _T_9154 | _T_8955; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_8957 = _T_3861 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9156 = _T_9155 | _T_8957; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_8959 = _T_3865 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9157 = _T_9156 | _T_8959; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_8961 = _T_3869 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9158 = _T_9157 | _T_8961; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_8963 = _T_3873 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9159 = _T_9158 | _T_8963; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_8965 = _T_3877 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9160 = _T_9159 | _T_8965; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_8967 = _T_3881 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9161 = _T_9160 | _T_8967; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_8969 = _T_3885 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9162 = _T_9161 | _T_8969; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_8971 = _T_3889 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9163 = _T_9162 | _T_8971; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_8973 = _T_3893 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9164 = _T_9163 | _T_8973; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_8975 = _T_3897 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9165 = _T_9164 | _T_8975; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_8977 = _T_3901 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9166 = _T_9165 | _T_8977; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_8979 = _T_3905 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9167 = _T_9166 | _T_8979; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_8981 = _T_3909 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9168 = _T_9167 | _T_8981; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_8983 = _T_3913 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9169 = _T_9168 | _T_8983; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_8985 = _T_3917 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9170 = _T_9169 | _T_8985; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_8987 = _T_3921 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9171 = _T_9170 | _T_8987; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_8989 = _T_3925 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9172 = _T_9171 | _T_8989; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_8991 = _T_3929 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9173 = _T_9172 | _T_8991; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_8993 = _T_3933 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9174 = _T_9173 | _T_8993; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_8995 = _T_3937 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9175 = _T_9174 | _T_8995; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_8997 = _T_3941 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9176 = _T_9175 | _T_8997; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_8999 = _T_3945 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9177 = _T_9176 | _T_8999; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9001 = _T_3949 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9178 = _T_9177 | _T_9001; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9003 = _T_3953 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9179 = _T_9178 | _T_9003; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9005 = _T_3957 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9180 = _T_9179 | _T_9005; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9007 = _T_3961 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9181 = _T_9180 | _T_9007; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9009 = _T_3965 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9182 = _T_9181 | _T_9009; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9011 = _T_3969 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9183 = _T_9182 | _T_9011; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9013 = _T_3973 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9184 = _T_9183 | _T_9013; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9015 = _T_3977 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9185 = _T_9184 | _T_9015; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9017 = _T_3981 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9186 = _T_9185 | _T_9017; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9019 = _T_3985 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9187 = _T_9186 | _T_9019; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9021 = _T_3989 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9188 = _T_9187 | _T_9021; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9023 = _T_3993 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9189 = _T_9188 | _T_9023; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9025 = _T_3997 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9190 = _T_9189 | _T_9025; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9027 = _T_4001 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9191 = _T_9190 | _T_9027; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9029 = _T_4005 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9192 = _T_9191 | _T_9029; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9031 = _T_4009 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9193 = _T_9192 | _T_9031; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9033 = _T_4013 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9194 = _T_9193 | _T_9033; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9035 = _T_4017 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9195 = _T_9194 | _T_9035; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9037 = _T_4021 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9196 = _T_9195 | _T_9037; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9039 = _T_4025 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9197 = _T_9196 | _T_9039; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9041 = _T_4029 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9198 = _T_9197 | _T_9041; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9043 = _T_4033 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9199 = _T_9198 | _T_9043; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9045 = _T_4037 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9200 = _T_9199 | _T_9045; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9047 = _T_4041 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9201 = _T_9200 | _T_9047; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9049 = _T_4045 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9202 = _T_9201 | _T_9049; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9051 = _T_4049 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9203 = _T_9202 | _T_9051; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9053 = _T_4053 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9204 = _T_9203 | _T_9053; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9055 = _T_4057 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9205 = _T_9204 | _T_9055; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9057 = _T_4061 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9206 = _T_9205 | _T_9057; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9059 = _T_4065 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9207 = _T_9206 | _T_9059; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9061 = _T_4069 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9208 = _T_9207 | _T_9061; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9063 = _T_4073 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9209 = _T_9208 | _T_9063; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9065 = _T_4077 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9210 = _T_9209 | _T_9065; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9067 = _T_4081 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9211 = _T_9210 | _T_9067; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9069 = _T_4085 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9212 = _T_9211 | _T_9069; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9071 = _T_4089 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9213 = _T_9212 | _T_9071; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9073 = _T_4093 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9214 = _T_9213 | _T_9073; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9075 = _T_4097 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9215 = _T_9214 | _T_9075; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9077 = _T_4101 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9216 = _T_9215 | _T_9077; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9079 = _T_4105 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9217 = _T_9216 | _T_9079; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9081 = _T_4109 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9218 = _T_9217 | _T_9081; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9083 = _T_4113 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9219 = _T_9218 | _T_9083; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9085 = _T_4117 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9220 = _T_9219 | _T_9085; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9087 = _T_4121 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9221 = _T_9220 | _T_9087; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9089 = _T_4125 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9222 = _T_9221 | _T_9089; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9091 = _T_4129 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9223 = _T_9222 | _T_9091; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9093 = _T_4133 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9224 = _T_9223 | _T_9093; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9095 = _T_4137 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9225 = _T_9224 | _T_9095; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9097 = _T_4141 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9226 = _T_9225 | _T_9097; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9099 = _T_4145 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9227 = _T_9226 | _T_9099; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9101 = _T_4149 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9228 = _T_9227 | _T_9101; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8464 = _T_3641 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 760:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8466 = _T_3645 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8719 = _T_8464 | _T_8466; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8468 = _T_3649 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8720 = _T_8719 | _T_8468; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8470 = _T_3653 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8721 = _T_8720 | _T_8470; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8472 = _T_3657 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8722 = _T_8721 | _T_8472; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8474 = _T_3661 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8723 = _T_8722 | _T_8474; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8476 = _T_3665 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8724 = _T_8723 | _T_8476; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8478 = _T_3669 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8725 = _T_8724 | _T_8478; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8480 = _T_3673 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8726 = _T_8725 | _T_8480; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8482 = _T_3677 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8727 = _T_8726 | _T_8482; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8484 = _T_3681 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8728 = _T_8727 | _T_8484; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8486 = _T_3685 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8729 = _T_8728 | _T_8486; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8488 = _T_3689 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8730 = _T_8729 | _T_8488; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8490 = _T_3693 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8731 = _T_8730 | _T_8490; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8492 = _T_3697 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8732 = _T_8731 | _T_8492; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8494 = _T_3701 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8733 = _T_8732 | _T_8494; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8496 = _T_3705 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8734 = _T_8733 | _T_8496; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8498 = _T_3709 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8735 = _T_8734 | _T_8498; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8500 = _T_3713 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8736 = _T_8735 | _T_8500; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8502 = _T_3717 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8737 = _T_8736 | _T_8502; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8504 = _T_3721 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8738 = _T_8737 | _T_8504; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8506 = _T_3725 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8739 = _T_8738 | _T_8506; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8508 = _T_3729 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8740 = _T_8739 | _T_8508; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8510 = _T_3733 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8741 = _T_8740 | _T_8510; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8512 = _T_3737 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8742 = _T_8741 | _T_8512; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8514 = _T_3741 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8743 = _T_8742 | _T_8514; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8516 = _T_3745 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8744 = _T_8743 | _T_8516; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8518 = _T_3749 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8745 = _T_8744 | _T_8518; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8520 = _T_3753 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8746 = _T_8745 | _T_8520; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8522 = _T_3757 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8747 = _T_8746 | _T_8522; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_8524 = _T_3761 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8748 = _T_8747 | _T_8524; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_8526 = _T_3765 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8749 = _T_8748 | _T_8526; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_8528 = _T_3769 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8750 = _T_8749 | _T_8528; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_8530 = _T_3773 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8751 = _T_8750 | _T_8530; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_8532 = _T_3777 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8752 = _T_8751 | _T_8532; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_8534 = _T_3781 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8753 = _T_8752 | _T_8534; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_8536 = _T_3785 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8754 = _T_8753 | _T_8536; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_8538 = _T_3789 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8755 = _T_8754 | _T_8538; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_8540 = _T_3793 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8756 = _T_8755 | _T_8540; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_8542 = _T_3797 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8757 = _T_8756 | _T_8542; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_8544 = _T_3801 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8758 = _T_8757 | _T_8544; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_8546 = _T_3805 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8759 = _T_8758 | _T_8546; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_8548 = _T_3809 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8760 = _T_8759 | _T_8548; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_8550 = _T_3813 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8761 = _T_8760 | _T_8550; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_8552 = _T_3817 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8762 = _T_8761 | _T_8552; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_8554 = _T_3821 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8763 = _T_8762 | _T_8554; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_8556 = _T_3825 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8764 = _T_8763 | _T_8556; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_8558 = _T_3829 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8765 = _T_8764 | _T_8558; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_8560 = _T_3833 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8766 = _T_8765 | _T_8560; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_8562 = _T_3837 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8767 = _T_8766 | _T_8562; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_8564 = _T_3841 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8768 = _T_8767 | _T_8564; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_8566 = _T_3845 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8769 = _T_8768 | _T_8566; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_8568 = _T_3849 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8770 = _T_8769 | _T_8568; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_8570 = _T_3853 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8771 = _T_8770 | _T_8570; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_8572 = _T_3857 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8772 = _T_8771 | _T_8572; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_8574 = _T_3861 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8773 = _T_8772 | _T_8574; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_8576 = _T_3865 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8774 = _T_8773 | _T_8576; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_8578 = _T_3869 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8775 = _T_8774 | _T_8578; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_8580 = _T_3873 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8776 = _T_8775 | _T_8580; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_8582 = _T_3877 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8777 = _T_8776 | _T_8582; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_8584 = _T_3881 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8778 = _T_8777 | _T_8584; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_8586 = _T_3885 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8779 = _T_8778 | _T_8586; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_8588 = _T_3889 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8780 = _T_8779 | _T_8588; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_8590 = _T_3893 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8781 = _T_8780 | _T_8590; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_8592 = _T_3897 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8782 = _T_8781 | _T_8592; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_8594 = _T_3901 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8783 = _T_8782 | _T_8594; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_8596 = _T_3905 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8784 = _T_8783 | _T_8596; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_8598 = _T_3909 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8785 = _T_8784 | _T_8598; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_8600 = _T_3913 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8786 = _T_8785 | _T_8600; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_8602 = _T_3917 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8787 = _T_8786 | _T_8602; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_8604 = _T_3921 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8788 = _T_8787 | _T_8604; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_8606 = _T_3925 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8789 = _T_8788 | _T_8606; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_8608 = _T_3929 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8790 = _T_8789 | _T_8608; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_8610 = _T_3933 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8791 = _T_8790 | _T_8610; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_8612 = _T_3937 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8792 = _T_8791 | _T_8612; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_8614 = _T_3941 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8793 = _T_8792 | _T_8614; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_8616 = _T_3945 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8794 = _T_8793 | _T_8616; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_8618 = _T_3949 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8795 = _T_8794 | _T_8618; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_8620 = _T_3953 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8796 = _T_8795 | _T_8620; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_8622 = _T_3957 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8797 = _T_8796 | _T_8622; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_8624 = _T_3961 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8798 = _T_8797 | _T_8624; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_8626 = _T_3965 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8799 = _T_8798 | _T_8626; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_8628 = _T_3969 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8800 = _T_8799 | _T_8628; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_8630 = _T_3973 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8801 = _T_8800 | _T_8630; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_8632 = _T_3977 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8802 = _T_8801 | _T_8632; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_8634 = _T_3981 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8803 = _T_8802 | _T_8634; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_8636 = _T_3985 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8804 = _T_8803 | _T_8636; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_8638 = _T_3989 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8805 = _T_8804 | _T_8638; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_8640 = _T_3993 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8806 = _T_8805 | _T_8640; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_8642 = _T_3997 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8807 = _T_8806 | _T_8642; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_8644 = _T_4001 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8808 = _T_8807 | _T_8644; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_8646 = _T_4005 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8809 = _T_8808 | _T_8646; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_8648 = _T_4009 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8810 = _T_8809 | _T_8648; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_8650 = _T_4013 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8811 = _T_8810 | _T_8650; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_8652 = _T_4017 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8812 = _T_8811 | _T_8652; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_8654 = _T_4021 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8813 = _T_8812 | _T_8654; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_8656 = _T_4025 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8814 = _T_8813 | _T_8656; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_8658 = _T_4029 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8815 = _T_8814 | _T_8658; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_8660 = _T_4033 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8816 = _T_8815 | _T_8660; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_8662 = _T_4037 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8817 = _T_8816 | _T_8662; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_8664 = _T_4041 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8818 = _T_8817 | _T_8664; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_8666 = _T_4045 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8819 = _T_8818 | _T_8666; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_8668 = _T_4049 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8820 = _T_8819 | _T_8668; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_8670 = _T_4053 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8821 = _T_8820 | _T_8670; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_8672 = _T_4057 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8822 = _T_8821 | _T_8672; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_8674 = _T_4061 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8823 = _T_8822 | _T_8674; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_8676 = _T_4065 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8824 = _T_8823 | _T_8676; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_8678 = _T_4069 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8825 = _T_8824 | _T_8678; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_8680 = _T_4073 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8826 = _T_8825 | _T_8680; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_8682 = _T_4077 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8827 = _T_8826 | _T_8682; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_8684 = _T_4081 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8828 = _T_8827 | _T_8684; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_8686 = _T_4085 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8829 = _T_8828 | _T_8686; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_8688 = _T_4089 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8830 = _T_8829 | _T_8688; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_8690 = _T_4093 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8831 = _T_8830 | _T_8690; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_8692 = _T_4097 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8832 = _T_8831 | _T_8692; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_8694 = _T_4101 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8833 = _T_8832 | _T_8694; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_8696 = _T_4105 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8834 = _T_8833 | _T_8696; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_8698 = _T_4109 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8835 = _T_8834 | _T_8698; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_8700 = _T_4113 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8836 = _T_8835 | _T_8700; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_8702 = _T_4117 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8837 = _T_8836 | _T_8702; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_8704 = _T_4121 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8838 = _T_8837 | _T_8704; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_8706 = _T_4125 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8839 = _T_8838 | _T_8706; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_8708 = _T_4129 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8840 = _T_8839 | _T_8708; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_8710 = _T_4133 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8841 = _T_8840 | _T_8710; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_8712 = _T_4137 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8842 = _T_8841 | _T_8712; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_8714 = _T_4141 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8843 = _T_8842 | _T_8714; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_8716 = _T_4145 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8844 = _T_8843 | _T_8716; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_8718 = _T_4149 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8845 = _T_8844 | _T_8718; // @[el2_ifu_mem_ctl.scala 760:91]
  wire [1:0] ic_tag_valid_unq = {_T_9228,_T_8845}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 833:54]
  wire [1:0] _T_9267 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9268 = ic_debug_way_ff & _T_9267; // @[el2_ifu_mem_ctl.scala 814:67]
  wire [1:0] _T_9269 = ic_tag_valid_unq & _T_9268; // @[el2_ifu_mem_ctl.scala 814:48]
  wire  ic_debug_tag_val_rd_out = |_T_9269; // @[el2_ifu_mem_ctl.scala 814:115]
  wire [65:0] _T_364 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_365; // @[el2_ifu_mem_ctl.scala 362:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_1709; // @[el2_ifu_mem_ctl.scala 374:80]
  wire  _T_405 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 379:98]
  wire  sel_byp_data = _T_409 & _T_405; // @[el2_ifu_mem_ctl.scala 379:96]
  wire [63:0] _T_416 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_417 = _T_416 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 386:64]
  wire [63:0] _T_419 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_1271 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 455:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_785 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_833 = _T_785 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_788 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_834 = _T_788 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_849 = _T_833 | _T_834; // @[Mux.scala 27:72]
  wire  _T_791 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_835 = _T_791 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_850 = _T_849 | _T_835; // @[Mux.scala 27:72]
  wire  _T_794 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_836 = _T_794 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_851 = _T_850 | _T_836; // @[Mux.scala 27:72]
  wire  _T_797 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_837 = _T_797 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_852 = _T_851 | _T_837; // @[Mux.scala 27:72]
  wire  _T_800 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_838 = _T_800 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_853 = _T_852 | _T_838; // @[Mux.scala 27:72]
  wire  _T_803 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_839 = _T_803 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_854 = _T_853 | _T_839; // @[Mux.scala 27:72]
  wire  _T_806 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_840 = _T_806 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_855 = _T_854 | _T_840; // @[Mux.scala 27:72]
  wire  _T_809 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_841 = _T_809 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_856 = _T_855 | _T_841; // @[Mux.scala 27:72]
  wire  _T_812 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_842 = _T_812 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_857 = _T_856 | _T_842; // @[Mux.scala 27:72]
  wire  _T_815 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_843 = _T_815 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_858 = _T_857 | _T_843; // @[Mux.scala 27:72]
  wire  _T_818 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_844 = _T_818 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_859 = _T_858 | _T_844; // @[Mux.scala 27:72]
  wire  _T_821 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_845 = _T_821 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_860 = _T_859 | _T_845; // @[Mux.scala 27:72]
  wire  _T_824 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_846 = _T_824 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_861 = _T_860 | _T_846; // @[Mux.scala 27:72]
  wire  _T_827 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_847 = _T_827 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_862 = _T_861 | _T_847; // @[Mux.scala 27:72]
  wire  _T_830 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_848 = _T_830 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_863 = _T_862 | _T_848; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_865 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_913 = _T_865 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_868 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_914 = _T_868 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_929 = _T_913 | _T_914; // @[Mux.scala 27:72]
  wire  _T_871 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_915 = _T_871 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_930 = _T_929 | _T_915; // @[Mux.scala 27:72]
  wire  _T_874 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_916 = _T_874 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_931 = _T_930 | _T_916; // @[Mux.scala 27:72]
  wire  _T_877 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_917 = _T_877 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_932 = _T_931 | _T_917; // @[Mux.scala 27:72]
  wire  _T_880 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_918 = _T_880 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_933 = _T_932 | _T_918; // @[Mux.scala 27:72]
  wire  _T_883 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_919 = _T_883 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_934 = _T_933 | _T_919; // @[Mux.scala 27:72]
  wire  _T_886 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_920 = _T_886 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_935 = _T_934 | _T_920; // @[Mux.scala 27:72]
  wire  _T_889 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_921 = _T_889 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_936 = _T_935 | _T_921; // @[Mux.scala 27:72]
  wire  _T_892 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_922 = _T_892 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_937 = _T_936 | _T_922; // @[Mux.scala 27:72]
  wire  _T_895 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_923 = _T_895 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_938 = _T_937 | _T_923; // @[Mux.scala 27:72]
  wire  _T_898 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_924 = _T_898 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_939 = _T_938 | _T_924; // @[Mux.scala 27:72]
  wire  _T_901 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_925 = _T_901 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_940 = _T_939 | _T_925; // @[Mux.scala 27:72]
  wire  _T_904 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_926 = _T_904 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_941 = _T_940 | _T_926; // @[Mux.scala 27:72]
  wire  _T_907 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_927 = _T_907 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_942 = _T_941 | _T_927; // @[Mux.scala 27:72]
  wire  _T_910 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_928 = _T_910 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_943 = _T_942 | _T_928; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_945 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_993 = _T_945 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_948 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_994 = _T_948 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1009 = _T_993 | _T_994; // @[Mux.scala 27:72]
  wire  _T_951 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_995 = _T_951 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1010 = _T_1009 | _T_995; // @[Mux.scala 27:72]
  wire  _T_954 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_996 = _T_954 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1011 = _T_1010 | _T_996; // @[Mux.scala 27:72]
  wire  _T_957 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_997 = _T_957 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1012 = _T_1011 | _T_997; // @[Mux.scala 27:72]
  wire  _T_960 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_998 = _T_960 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1013 = _T_1012 | _T_998; // @[Mux.scala 27:72]
  wire  _T_963 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_999 = _T_963 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1014 = _T_1013 | _T_999; // @[Mux.scala 27:72]
  wire  _T_966 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1000 = _T_966 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1015 = _T_1014 | _T_1000; // @[Mux.scala 27:72]
  wire  _T_969 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1001 = _T_969 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1016 = _T_1015 | _T_1001; // @[Mux.scala 27:72]
  wire  _T_972 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1002 = _T_972 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1017 = _T_1016 | _T_1002; // @[Mux.scala 27:72]
  wire  _T_975 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1003 = _T_975 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1018 = _T_1017 | _T_1003; // @[Mux.scala 27:72]
  wire  _T_978 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1004 = _T_978 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1019 = _T_1018 | _T_1004; // @[Mux.scala 27:72]
  wire  _T_981 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1005 = _T_981 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1020 = _T_1019 | _T_1005; // @[Mux.scala 27:72]
  wire  _T_984 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1006 = _T_984 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1021 = _T_1020 | _T_1006; // @[Mux.scala 27:72]
  wire  _T_987 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1007 = _T_987 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1022 = _T_1021 | _T_1007; // @[Mux.scala 27:72]
  wire  _T_990 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1008 = _T_990 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1023 = _T_1022 | _T_1008; // @[Mux.scala 27:72]
  wire [79:0] _T_1026 = {_T_863,_T_943,_T_1023}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1027 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1075 = _T_1027 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1030 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1076 = _T_1030 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1091 = _T_1075 | _T_1076; // @[Mux.scala 27:72]
  wire  _T_1033 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1077 = _T_1033 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1092 = _T_1091 | _T_1077; // @[Mux.scala 27:72]
  wire  _T_1036 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1078 = _T_1036 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1093 = _T_1092 | _T_1078; // @[Mux.scala 27:72]
  wire  _T_1039 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1079 = _T_1039 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1094 = _T_1093 | _T_1079; // @[Mux.scala 27:72]
  wire  _T_1042 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1080 = _T_1042 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1095 = _T_1094 | _T_1080; // @[Mux.scala 27:72]
  wire  _T_1045 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1081 = _T_1045 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1096 = _T_1095 | _T_1081; // @[Mux.scala 27:72]
  wire  _T_1048 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1082 = _T_1048 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1097 = _T_1096 | _T_1082; // @[Mux.scala 27:72]
  wire  _T_1051 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1083 = _T_1051 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1098 = _T_1097 | _T_1083; // @[Mux.scala 27:72]
  wire  _T_1054 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1084 = _T_1054 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1099 = _T_1098 | _T_1084; // @[Mux.scala 27:72]
  wire  _T_1057 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1085 = _T_1057 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1100 = _T_1099 | _T_1085; // @[Mux.scala 27:72]
  wire  _T_1060 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1086 = _T_1060 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1101 = _T_1100 | _T_1086; // @[Mux.scala 27:72]
  wire  _T_1063 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1087 = _T_1063 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1102 = _T_1101 | _T_1087; // @[Mux.scala 27:72]
  wire  _T_1066 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1088 = _T_1066 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1103 = _T_1102 | _T_1088; // @[Mux.scala 27:72]
  wire  _T_1069 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1089 = _T_1069 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1104 = _T_1103 | _T_1089; // @[Mux.scala 27:72]
  wire  _T_1072 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1090 = _T_1072 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1105 = _T_1104 | _T_1090; // @[Mux.scala 27:72]
  wire [31:0] _T_1155 = _T_785 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1156 = _T_788 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1171 = _T_1155 | _T_1156; // @[Mux.scala 27:72]
  wire [31:0] _T_1157 = _T_791 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1172 = _T_1171 | _T_1157; // @[Mux.scala 27:72]
  wire [31:0] _T_1158 = _T_794 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1173 = _T_1172 | _T_1158; // @[Mux.scala 27:72]
  wire [31:0] _T_1159 = _T_797 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1174 = _T_1173 | _T_1159; // @[Mux.scala 27:72]
  wire [31:0] _T_1160 = _T_800 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1175 = _T_1174 | _T_1160; // @[Mux.scala 27:72]
  wire [31:0] _T_1161 = _T_803 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1176 = _T_1175 | _T_1161; // @[Mux.scala 27:72]
  wire [31:0] _T_1162 = _T_806 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1177 = _T_1176 | _T_1162; // @[Mux.scala 27:72]
  wire [31:0] _T_1163 = _T_809 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1178 = _T_1177 | _T_1163; // @[Mux.scala 27:72]
  wire [31:0] _T_1164 = _T_812 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1179 = _T_1178 | _T_1164; // @[Mux.scala 27:72]
  wire [31:0] _T_1165 = _T_815 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1180 = _T_1179 | _T_1165; // @[Mux.scala 27:72]
  wire [31:0] _T_1166 = _T_818 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1181 = _T_1180 | _T_1166; // @[Mux.scala 27:72]
  wire [31:0] _T_1167 = _T_821 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1182 = _T_1181 | _T_1167; // @[Mux.scala 27:72]
  wire [31:0] _T_1168 = _T_824 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1183 = _T_1182 | _T_1168; // @[Mux.scala 27:72]
  wire [31:0] _T_1169 = _T_827 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1184 = _T_1183 | _T_1169; // @[Mux.scala 27:72]
  wire [31:0] _T_1170 = _T_830 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1185 = _T_1184 | _T_1170; // @[Mux.scala 27:72]
  wire [79:0] _T_1268 = {_T_1105,_T_1185,_T_943}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1271 ? _T_1026 : _T_1268; // @[el2_ifu_mem_ctl.scala 451:37]
  wire [79:0] _T_1273 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_1271 ? ic_byp_data_only_pre_new : _T_1273; // @[el2_ifu_mem_ctl.scala 455:30]
  wire [79:0] _GEN_793 = {{16'd0}, _T_419}; // @[el2_ifu_mem_ctl.scala 386:109]
  wire [79:0] _T_420 = _GEN_793 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 386:109]
  wire [79:0] _GEN_794 = {{16'd0}, _T_417}; // @[el2_ifu_mem_ctl.scala 386:83]
  wire [79:0] ic_premux_data = _GEN_794 | _T_420; // @[el2_ifu_mem_ctl.scala 386:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 393:38]
  wire [1:0] _T_429 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 397:8]
  wire [7:0] _T_526 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_531 = ic_miss_buff_data_error[0] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  _T_1777 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 629:47]
  wire  _T_1778 = _T_1777 & _T_13; // @[el2_ifu_mem_ctl.scala 629:50]
  wire  bus_ifu_wr_data_error = _T_1778 & miss_pending; // @[el2_ifu_mem_ctl.scala 629:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_531; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_535 = ic_miss_buff_data_error[1] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_535; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_539 = ic_miss_buff_data_error[2] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_539; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_543 = ic_miss_buff_data_error[3] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_543; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_547 = ic_miss_buff_data_error[4] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_547; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_551 = ic_miss_buff_data_error[5] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_551; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_555 = ic_miss_buff_data_error[6] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_555; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_559 = ic_miss_buff_data_error[7] & _T_497; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_559; // @[el2_ifu_mem_ctl.scala 417:72]
  wire [7:0] _T_566 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_1583 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1591 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 498:65]
  wire  _T_1592 = _T_1591 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 498:88]
  wire  _T_1594 = _T_1592 & _T_1705; // @[el2_ifu_mem_ctl.scala 498:112]
  wire  _T_1595 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1596 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 503:50]
  wire  _T_1598 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1604 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1606 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_1604 | _T_1606; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_1598 ? _T_1596 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_1595 ? _T_1596 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_1583 ? _T_1594 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_1583 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_1597 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 504:56]
  wire  _GEN_43 = _T_1595 & _T_1597; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_1583 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 489:58]
  wire  _T_1580 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 488:49]
  wire  _T_1585 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 497:87]
  wire  _T_1599 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 507:54]
  wire  _T_1600 = _T_1599 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 507:84]
  wire  _T_1609 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 528:66]
  wire  _T_1610 = io_dec_tlu_flush_err_wb & _T_1609; // @[el2_ifu_mem_ctl.scala 528:52]
  wire  _T_1612 = _T_1610 & _T_1705; // @[el2_ifu_mem_ctl.scala 528:81]
  wire  _T_1614 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 531:59]
  wire  _T_1615 = _T_1614 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 531:86]
  wire  _T_1629 = _T_1614 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 534:81]
  wire  _T_1630 = _T_1629 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 534:103]
  wire  _T_1631 = _T_1630 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 534:126]
  wire  _T_1651 = _T_1629 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 541:103]
  wire  _T_1658 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 546:62]
  wire  _T_1659 = io_dec_tlu_flush_lower_wb & _T_1658; // @[el2_ifu_mem_ctl.scala 546:60]
  wire  _T_1660 = _T_1659 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 546:88]
  wire  _T_1661 = _T_1660 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 546:115]
  wire  _GEN_50 = _T_1657 & _T_1615; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_1640 ? _T_1651 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_1640 | _T_1657; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_1613 ? _T_1631 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_1613 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_1608 ? _T_1612 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_1673 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 563:64]
  wire  _T_1675 = _T_1673 & _T_1705; // @[el2_ifu_mem_ctl.scala 563:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_1677 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 563:133]
  wire  _T_1678 = _T_1677 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 563:164]
  wire  _T_1679 = _T_1678 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 563:184]
  wire  _T_1680 = _T_1679 & miss_pending; // @[el2_ifu_mem_ctl.scala 563:204]
  wire  _T_1681 = ~_T_1680; // @[el2_ifu_mem_ctl.scala 563:112]
  wire  ifc_bus_ic_req_ff_in = _T_1675 & _T_1681; // @[el2_ifu_mem_ctl.scala 563:110]
  wire  _T_1682 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 564:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 595:45]
  wire  _T_1699 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 598:35]
  wire  _T_1700 = _T_1699 & miss_pending; // @[el2_ifu_mem_ctl.scala 598:53]
  wire  bus_cmd_sent = _T_1700 & _T_1705; // @[el2_ifu_mem_ctl.scala 598:68]
  wire [2:0] _T_1690 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1692 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1694 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 596:51]
  wire  _T_1720 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 606:73]
  wire  _T_1721 = _T_1706 & _T_1720; // @[el2_ifu_mem_ctl.scala 606:71]
  wire  _T_1723 = last_data_recieved_ff & _T_497; // @[el2_ifu_mem_ctl.scala 606:114]
  wire  last_data_recieved_in = _T_1721 | _T_1723; // @[el2_ifu_mem_ctl.scala 606:89]
  wire [2:0] _T_1729 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 611:45]
  wire  _T_1732 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 612:81]
  wire  _T_1733 = _T_1732 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 612:97]
  wire  _T_1735 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 614:48]
  wire  _T_1736 = _T_1735 & miss_pending; // @[el2_ifu_mem_ctl.scala 614:68]
  wire  bus_inc_cmd_beat_cnt = _T_1736 & _T_1705; // @[el2_ifu_mem_ctl.scala 614:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 616:57]
  wire  _T_1740 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 617:31]
  wire  _T_1741 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 617:71]
  wire  _T_1742 = _T_1741 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 617:87]
  wire  _T_1743 = ~_T_1742; // @[el2_ifu_mem_ctl.scala 617:55]
  wire  bus_hold_cmd_beat_cnt = _T_1740 & _T_1743; // @[el2_ifu_mem_ctl.scala 617:53]
  wire  _T_1744 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 618:46]
  wire  bus_cmd_beat_en = _T_1744 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 618:62]
  wire [2:0] _T_1747 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 620:46]
  wire [2:0] _T_1749 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1750 = bus_inc_cmd_beat_cnt ? _T_1747 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1751 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1753 = _T_1749 | _T_1750; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_1753 | _T_1751; // @[Mux.scala 27:72]
  wire  _T_1757 = _T_1733 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 621:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 632:62]
  wire  _T_1785 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 637:50]
  wire  _T_1786 = io_ifc_dma_access_ok & _T_1785; // @[el2_ifu_mem_ctl.scala 637:47]
  wire  _T_1787 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 637:70]
  wire  ifc_dma_access_ok_d = _T_1786 & _T_1787; // @[el2_ifu_mem_ctl.scala 637:68]
  wire  _T_1791 = _T_1786 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 638:72]
  wire  _T_1792 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 638:111]
  wire  _T_1793 = _T_1791 & _T_1792; // @[el2_ifu_mem_ctl.scala 638:97]
  wire  ifc_dma_access_q_ok = _T_1793 & _T_1787; // @[el2_ifu_mem_ctl.scala 638:127]
  wire  _T_1796 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 641:40]
  wire  _T_1797 = _T_1796 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 641:58]
  wire  _T_1800 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 642:60]
  wire  _T_1801 = _T_1796 & _T_1800; // @[el2_ifu_mem_ctl.scala 642:58]
  wire  _T_1802 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 642:104]
  wire [2:0] _T_1807 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_1913 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_1922 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_1913}; // @[el2_lib.scala 268:22]
  wire  _T_1923 = ^_T_1922; // @[el2_lib.scala 268:29]
  wire [8:0] _T_1931 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_1940 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_1931}; // @[el2_lib.scala 268:39]
  wire  _T_1941 = ^_T_1940; // @[el2_lib.scala 268:46]
  wire [8:0] _T_1949 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_1958 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_1949}; // @[el2_lib.scala 268:56]
  wire  _T_1959 = ^_T_1958; // @[el2_lib.scala 268:63]
  wire [6:0] _T_1965 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_1973 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_1965}; // @[el2_lib.scala 268:73]
  wire  _T_1974 = ^_T_1973; // @[el2_lib.scala 268:80]
  wire [14:0] _T_1988 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_1965}; // @[el2_lib.scala 268:90]
  wire  _T_1989 = ^_T_1988; // @[el2_lib.scala 268:97]
  wire [5:0] _T_1994 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_1995 = ^_T_1994; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2000 = {_T_1923,_T_1941,_T_1959,_T_1974,_T_1989,_T_1995}; // @[Cat.scala 29:58]
  wire  _T_2001 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2002 = ^_T_2000; // @[el2_lib.scala 269:23]
  wire  _T_2003 = _T_2001 ^ _T_2002; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2109 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2118 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2109}; // @[el2_lib.scala 268:22]
  wire  _T_2119 = ^_T_2118; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2127 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2136 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2127}; // @[el2_lib.scala 268:39]
  wire  _T_2137 = ^_T_2136; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2145 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2154 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2145}; // @[el2_lib.scala 268:56]
  wire  _T_2155 = ^_T_2154; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2161 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2169 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2161}; // @[el2_lib.scala 268:73]
  wire  _T_2170 = ^_T_2169; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2184 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2161}; // @[el2_lib.scala 268:90]
  wire  _T_2185 = ^_T_2184; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2190 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_2191 = ^_T_2190; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2196 = {_T_2119,_T_2137,_T_2155,_T_2170,_T_2185,_T_2191}; // @[Cat.scala 29:58]
  wire  _T_2197 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_2198 = ^_T_2196; // @[el2_lib.scala 269:23]
  wire  _T_2199 = _T_2197 ^ _T_2198; // @[el2_lib.scala 269:18]
  wire [6:0] _T_2200 = {_T_2199,_T_2119,_T_2137,_T_2155,_T_2170,_T_2185,_T_2191}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2003,_T_1923,_T_1941,_T_1959,_T_1974,_T_1989,_T_1995,_T_2200}; // @[Cat.scala 29:58]
  wire  _T_2202 = ~_T_1796; // @[el2_ifu_mem_ctl.scala 647:45]
  wire  _T_2203 = iccm_correct_ecc & _T_2202; // @[el2_ifu_mem_ctl.scala 647:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_2204 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_2211 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 661:53]
  wire  _T_2543 = _T_2455[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2541 = _T_2455[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2539 = _T_2455[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2537 = _T_2455[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2535 = _T_2455[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2533 = _T_2455[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2531 = _T_2455[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2529 = _T_2455[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2527 = _T_2455[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2525 = _T_2455[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2601 = {_T_2543,_T_2541,_T_2539,_T_2537,_T_2535,_T_2533,_T_2531,_T_2529,_T_2527,_T_2525}; // @[el2_lib.scala 310:69]
  wire  _T_2523 = _T_2455[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2521 = _T_2455[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2519 = _T_2455[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2517 = _T_2455[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2515 = _T_2455[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2513 = _T_2455[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2511 = _T_2455[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2509 = _T_2455[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2507 = _T_2455[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2505 = _T_2455[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2592 = {_T_2523,_T_2521,_T_2519,_T_2517,_T_2515,_T_2513,_T_2511,_T_2509,_T_2507,_T_2505}; // @[el2_lib.scala 310:69]
  wire  _T_2503 = _T_2455[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2501 = _T_2455[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2499 = _T_2455[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2497 = _T_2455[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2495 = _T_2455[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2493 = _T_2455[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2491 = _T_2455[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2489 = _T_2455[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2487 = _T_2455[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2485 = _T_2455[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2582 = {_T_2503,_T_2501,_T_2499,_T_2497,_T_2495,_T_2493,_T_2491,_T_2489,_T_2487,_T_2485}; // @[el2_lib.scala 310:69]
  wire  _T_2483 = _T_2455[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2481 = _T_2455[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2479 = _T_2455[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2477 = _T_2455[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2475 = _T_2455[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2473 = _T_2455[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2471 = _T_2455[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2469 = _T_2455[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2467 = _T_2455[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_2583 = {_T_2582,_T_2483,_T_2481,_T_2479,_T_2477,_T_2475,_T_2473,_T_2471,_T_2469,_T_2467}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_2603 = {_T_2601,_T_2592,_T_2583}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2558 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2564 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_2558}; // @[Cat.scala 29:58]
  wire [38:0] _T_2604 = _T_2603 ^ _T_2564; // @[el2_lib.scala 310:76]
  wire [38:0] _T_2605 = _T_2459 ? _T_2604 : _T_2564; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_2605[37:32],_T_2605[30:16],_T_2605[14:8],_T_2605[6:4],_T_2605[2]}; // @[Cat.scala 29:58]
  wire  _T_2928 = _T_2840[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2926 = _T_2840[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2924 = _T_2840[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2922 = _T_2840[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2920 = _T_2840[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2918 = _T_2840[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2916 = _T_2840[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2914 = _T_2840[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2912 = _T_2840[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2910 = _T_2840[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2986 = {_T_2928,_T_2926,_T_2924,_T_2922,_T_2920,_T_2918,_T_2916,_T_2914,_T_2912,_T_2910}; // @[el2_lib.scala 310:69]
  wire  _T_2908 = _T_2840[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2906 = _T_2840[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2904 = _T_2840[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2902 = _T_2840[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2900 = _T_2840[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2898 = _T_2840[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2896 = _T_2840[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2894 = _T_2840[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2892 = _T_2840[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2890 = _T_2840[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2977 = {_T_2908,_T_2906,_T_2904,_T_2902,_T_2900,_T_2898,_T_2896,_T_2894,_T_2892,_T_2890}; // @[el2_lib.scala 310:69]
  wire  _T_2888 = _T_2840[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2886 = _T_2840[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2884 = _T_2840[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2882 = _T_2840[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2880 = _T_2840[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2878 = _T_2840[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2876 = _T_2840[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2874 = _T_2840[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2872 = _T_2840[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2870 = _T_2840[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2967 = {_T_2888,_T_2886,_T_2884,_T_2882,_T_2880,_T_2878,_T_2876,_T_2874,_T_2872,_T_2870}; // @[el2_lib.scala 310:69]
  wire  _T_2868 = _T_2840[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2866 = _T_2840[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2864 = _T_2840[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2862 = _T_2840[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2860 = _T_2840[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2858 = _T_2840[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2856 = _T_2840[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2854 = _T_2840[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2852 = _T_2840[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_2968 = {_T_2967,_T_2868,_T_2866,_T_2864,_T_2862,_T_2860,_T_2858,_T_2856,_T_2854,_T_2852}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_2988 = {_T_2986,_T_2977,_T_2968}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2943 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2949 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_2943}; // @[Cat.scala 29:58]
  wire [38:0] _T_2989 = _T_2988 ^ _T_2949; // @[el2_lib.scala 310:76]
  wire [38:0] _T_2990 = _T_2844 ? _T_2989 : _T_2949; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_2990[37:32],_T_2990[30:16],_T_2990[14:8],_T_2990[6:4],_T_2990[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 653:35]
  wire  _T_2463 = ~_T_2455[6]; // @[el2_lib.scala 303:55]
  wire  _T_2464 = _T_2457 & _T_2463; // @[el2_lib.scala 303:53]
  wire  _T_2848 = ~_T_2840[6]; // @[el2_lib.scala 303:55]
  wire  _T_2849 = _T_2842 & _T_2848; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_2464,_T_2849}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 655:53]
  wire [63:0] _T_2215 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_2216 = {iccm_dma_rdata_1_muxed,_T_2605[37:32],_T_2605[30:16],_T_2605[14:8],_T_2605[6:4],_T_2605[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 657:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 658:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 663:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 667:70]
  wire  _T_2221 = _T_1796 & _T_1785; // @[el2_ifu_mem_ctl.scala 670:65]
  wire  _T_2224 = _T_2202 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 671:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_2225 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_2227 = _T_2224 ? {{1'd0}, _T_2225} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 671:8]
  wire [31:0] _T_2228 = _T_2221 ? io_dma_mem_addr : {{16'd0}, _T_2227}; // @[el2_ifu_mem_ctl.scala 670:25]
  wire  _T_2617 = _T_2455 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_2618 = _T_2605[38] ^ _T_2617; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_2618,_T_2605[31],_T_2605[15],_T_2605[7],_T_2605[3],_T_2605[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3002 = _T_2840 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3003 = _T_2990[38] ^ _T_3002; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3003,_T_2990[31],_T_2990[15],_T_2990[7],_T_2990[3],_T_2990[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3019 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 683:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 685:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 686:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 694:62]
  wire  _T_3027 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 688:76]
  wire  _T_3028 = io_iccm_rd_ecc_single_err & _T_3027; // @[el2_ifu_mem_ctl.scala 688:74]
  wire  _T_3030 = _T_3028 & _T_317; // @[el2_ifu_mem_ctl.scala 688:104]
  wire  iccm_ecc_write_status = _T_3030 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 688:127]
  wire  _T_3031 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 689:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3031 & _T_317; // @[el2_ifu_mem_ctl.scala 689:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 693:51]
  wire [13:0] _T_3036 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 692:102]
  wire [38:0] _T_3040 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3045 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 697:41]
  wire  _T_3046 = io_ifc_fetch_req_bf & _T_3045; // @[el2_ifu_mem_ctl.scala 697:39]
  wire  _T_3047 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 697:72]
  wire  _T_3048 = _T_3046 & _T_3047; // @[el2_ifu_mem_ctl.scala 697:70]
  wire  _T_3050 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 698:34]
  wire  _T_3051 = _T_1391 & _T_3050; // @[el2_ifu_mem_ctl.scala 698:32]
  wire  _T_3054 = _T_1407 & _T_3050; // @[el2_ifu_mem_ctl.scala 699:37]
  wire  _T_3055 = _T_3051 | _T_3054; // @[el2_ifu_mem_ctl.scala 698:88]
  wire  _T_3056 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 700:19]
  wire  _T_3058 = _T_3056 & _T_3050; // @[el2_ifu_mem_ctl.scala 700:41]
  wire  _T_3059 = _T_3055 | _T_3058; // @[el2_ifu_mem_ctl.scala 699:88]
  wire  _T_3060 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 701:19]
  wire  _T_3062 = _T_3060 & _T_3050; // @[el2_ifu_mem_ctl.scala 701:35]
  wire  _T_3063 = _T_3059 | _T_3062; // @[el2_ifu_mem_ctl.scala 700:88]
  wire  _T_3066 = _T_1406 & _T_3050; // @[el2_ifu_mem_ctl.scala 702:38]
  wire  _T_3067 = _T_3063 | _T_3066; // @[el2_ifu_mem_ctl.scala 701:88]
  wire  _T_3069 = _T_1407 & miss_state_en; // @[el2_ifu_mem_ctl.scala 703:37]
  wire  _T_3070 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 703:71]
  wire  _T_3071 = _T_3069 & _T_3070; // @[el2_ifu_mem_ctl.scala 703:54]
  wire  _T_3072 = _T_3067 | _T_3071; // @[el2_ifu_mem_ctl.scala 702:57]
  wire  _T_3073 = ~_T_3072; // @[el2_ifu_mem_ctl.scala 698:5]
  wire  _T_3074 = _T_3048 & _T_3073; // @[el2_ifu_mem_ctl.scala 697:96]
  wire  _T_3075 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 704:28]
  wire  _T_3077 = _T_3075 & _T_3045; // @[el2_ifu_mem_ctl.scala 704:50]
  wire  _T_3079 = _T_3077 & _T_3047; // @[el2_ifu_mem_ctl.scala 704:81]
  wire  _T_3088 = ~_T_108; // @[el2_ifu_mem_ctl.scala 707:106]
  wire  _T_3089 = _T_1391 & _T_3088; // @[el2_ifu_mem_ctl.scala 707:104]
  wire  _T_3090 = _T_1407 | _T_3089; // @[el2_ifu_mem_ctl.scala 707:77]
  wire  _T_3094 = ~_T_51; // @[el2_ifu_mem_ctl.scala 707:172]
  wire  _T_3095 = _T_3090 & _T_3094; // @[el2_ifu_mem_ctl.scala 707:170]
  wire  _T_3096 = ~_T_3095; // @[el2_ifu_mem_ctl.scala 707:44]
  wire  _T_3100 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 710:64]
  wire  _T_3101 = ~_T_3100; // @[el2_ifu_mem_ctl.scala 710:50]
  wire  _T_3102 = _T_276 & _T_3101; // @[el2_ifu_mem_ctl.scala 710:48]
  wire  _T_3103 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 710:81]
  wire  ic_valid = _T_3102 & _T_3103; // @[el2_ifu_mem_ctl.scala 710:79]
  wire  _T_3105 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 711:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 714:14]
  wire  _T_3108 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 717:74]
  wire  _T_9250 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 791:45]
  wire  way_status_wr_en = _T_9250 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 791:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3108; // @[el2_ifu_mem_ctl.scala 717:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 719:14]
  wire [2:0] _T_3112 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 723:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 787:41]
  wire  way_status_new = _T_9250 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 790:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 725:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  _T_3129 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3130 = _T_3129 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3131 = _T_3130 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3133 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3134 = _T_3133 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3135 = _T_3134 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3137 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3138 = _T_3137 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3139 = _T_3138 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3141 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3142 = _T_3141 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3143 = _T_3142 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3145 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3146 = _T_3145 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3147 = _T_3146 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3149 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3150 = _T_3149 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3151 = _T_3150 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3153 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3154 = _T_3153 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3155 = _T_3154 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3157 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3158 = _T_3157 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3159 = _T_3158 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3163 = _T_3130 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3167 = _T_3134 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3171 = _T_3138 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3175 = _T_3142 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3179 = _T_3146 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3183 = _T_3150 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3187 = _T_3154 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3191 = _T_3158 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3195 = _T_3130 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3199 = _T_3134 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3203 = _T_3138 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3207 = _T_3142 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3211 = _T_3146 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3215 = _T_3150 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3219 = _T_3154 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3223 = _T_3158 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3227 = _T_3130 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3231 = _T_3134 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3235 = _T_3138 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3239 = _T_3142 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3243 = _T_3146 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3247 = _T_3150 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3251 = _T_3154 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3255 = _T_3158 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3259 = _T_3130 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3263 = _T_3134 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3267 = _T_3138 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3271 = _T_3142 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3275 = _T_3146 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3279 = _T_3150 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3283 = _T_3154 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3287 = _T_3158 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3291 = _T_3130 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3295 = _T_3134 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3299 = _T_3138 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3303 = _T_3142 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3307 = _T_3146 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3311 = _T_3150 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3315 = _T_3154 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3319 = _T_3158 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3323 = _T_3130 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3327 = _T_3134 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3331 = _T_3138 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3335 = _T_3142 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3339 = _T_3146 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3343 = _T_3150 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3347 = _T_3154 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3351 = _T_3158 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3355 = _T_3130 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3359 = _T_3134 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3363 = _T_3138 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3367 = _T_3142 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3371 = _T_3146 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3375 = _T_3150 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3379 = _T_3154 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3383 = _T_3158 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3387 = _T_3130 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3391 = _T_3134 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3395 = _T_3138 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3399 = _T_3142 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3403 = _T_3146 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3407 = _T_3150 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3411 = _T_3154 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3415 = _T_3158 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3419 = _T_3130 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3423 = _T_3134 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3427 = _T_3138 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3431 = _T_3142 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3435 = _T_3146 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3439 = _T_3150 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3443 = _T_3154 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3447 = _T_3158 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3451 = _T_3130 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3455 = _T_3134 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3459 = _T_3138 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3463 = _T_3142 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3467 = _T_3146 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3471 = _T_3150 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3475 = _T_3154 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3479 = _T_3158 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3483 = _T_3130 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3487 = _T_3134 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3491 = _T_3138 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3495 = _T_3142 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3499 = _T_3146 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3503 = _T_3150 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3507 = _T_3154 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3511 = _T_3158 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3515 = _T_3130 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3519 = _T_3134 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3523 = _T_3138 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3527 = _T_3142 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3531 = _T_3146 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3535 = _T_3150 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3539 = _T_3154 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3543 = _T_3158 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3547 = _T_3130 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3551 = _T_3134 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3555 = _T_3138 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3559 = _T_3142 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3563 = _T_3146 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3567 = _T_3150 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3571 = _T_3154 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3575 = _T_3158 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3579 = _T_3130 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3583 = _T_3134 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3587 = _T_3138 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3591 = _T_3142 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3595 = _T_3146 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3599 = _T_3150 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3603 = _T_3154 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3607 = _T_3158 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3611 = _T_3130 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3615 = _T_3134 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3619 = _T_3138 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3623 = _T_3142 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3627 = _T_3146 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3631 = _T_3150 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3635 = _T_3154 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3639 = _T_3158 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_9256 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 794:84]
  wire  _T_9257 = _T_9256 & miss_pending; // @[el2_ifu_mem_ctl.scala 794:108]
  wire  bus_wren_last_1 = _T_9257 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 794:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_9259 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 796:73]
  wire  _T_9254 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 794:84]
  wire  _T_9255 = _T_9254 & miss_pending; // @[el2_ifu_mem_ctl.scala 794:108]
  wire  bus_wren_last_0 = _T_9255 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 794:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_9258 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 796:73]
  wire [1:0] ifu_tag_wren = {_T_9259,_T_9258}; // @[Cat.scala 29:58]
  wire [1:0] _T_9293 = _T_3108 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9293 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 829:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 740:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 742:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 746:14]
  wire  _T_4288 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4290 = _T_4288 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4292 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4294 = _T_4292 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4295 = _T_4290 | _T_4294; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4296 = _T_4295 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4300 = _T_4288 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4304 = _T_4292 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4305 = _T_4300 | _T_4304; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4306 = _T_4305 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_0 = {_T_4296,_T_4306}; // @[Cat.scala 29:58]
  wire  _T_4308 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4310 = _T_4308 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4312 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4314 = _T_4312 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4315 = _T_4310 | _T_4314; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4316 = _T_4315 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4320 = _T_4308 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4324 = _T_4312 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4325 = _T_4320 | _T_4324; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4326 = _T_4325 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_1 = {_T_4316,_T_4326}; // @[Cat.scala 29:58]
  wire  _T_4328 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4330 = _T_4328 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4332 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4334 = _T_4332 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4335 = _T_4330 | _T_4334; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4336 = _T_4335 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4340 = _T_4328 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4344 = _T_4332 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4345 = _T_4340 | _T_4344; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4346 = _T_4345 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_2 = {_T_4336,_T_4346}; // @[Cat.scala 29:58]
  wire  _T_4348 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4350 = _T_4348 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4352 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4354 = _T_4352 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4355 = _T_4350 | _T_4354; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4356 = _T_4355 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4360 = _T_4348 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4364 = _T_4352 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4365 = _T_4360 | _T_4364; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4366 = _T_4365 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_3 = {_T_4356,_T_4366}; // @[Cat.scala 29:58]
  wire  _T_4369 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 756:64]
  wire  _T_4370 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 756:91]
  wire  _T_4371 = _T_4369 & _T_4370; // @[el2_ifu_mem_ctl.scala 756:89]
  wire  _T_4374 = _T_3641 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4375 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4377 = _T_4375 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4379 = _T_4377 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4380 = _T_4374 | _T_4379; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4390 = _T_3645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4391 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4393 = _T_4391 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4395 = _T_4393 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4396 = _T_4390 | _T_4395; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4406 = _T_3649 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4407 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4409 = _T_4407 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4411 = _T_4409 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4412 = _T_4406 | _T_4411; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4422 = _T_3653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4423 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4425 = _T_4423 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4427 = _T_4425 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4428 = _T_4422 | _T_4427; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4438 = _T_3657 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4439 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4441 = _T_4439 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4443 = _T_4441 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4444 = _T_4438 | _T_4443; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4454 = _T_3661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4455 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4457 = _T_4455 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4459 = _T_4457 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4460 = _T_4454 | _T_4459; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4470 = _T_3665 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4471 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4473 = _T_4471 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4475 = _T_4473 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4476 = _T_4470 | _T_4475; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4486 = _T_3669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4487 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4489 = _T_4487 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4491 = _T_4489 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4492 = _T_4486 | _T_4491; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4502 = _T_3673 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4503 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4505 = _T_4503 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4507 = _T_4505 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4508 = _T_4502 | _T_4507; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4518 = _T_3677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4519 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4521 = _T_4519 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4523 = _T_4521 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4524 = _T_4518 | _T_4523; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4534 = _T_3681 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4535 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4537 = _T_4535 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4539 = _T_4537 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4540 = _T_4534 | _T_4539; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4550 = _T_3685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4551 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4553 = _T_4551 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4555 = _T_4553 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4556 = _T_4550 | _T_4555; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4566 = _T_3689 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4567 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4569 = _T_4567 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4571 = _T_4569 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4572 = _T_4566 | _T_4571; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4582 = _T_3693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4583 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4585 = _T_4583 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4587 = _T_4585 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4588 = _T_4582 | _T_4587; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4598 = _T_3697 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4599 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4601 = _T_4599 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4603 = _T_4601 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4604 = _T_4598 | _T_4603; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4614 = _T_3701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4615 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4617 = _T_4615 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4619 = _T_4617 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4620 = _T_4614 | _T_4619; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4630 = _T_3705 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4631 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4633 = _T_4631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4635 = _T_4633 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4636 = _T_4630 | _T_4635; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4646 = _T_3709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4647 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4649 = _T_4647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4651 = _T_4649 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4652 = _T_4646 | _T_4651; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4662 = _T_3713 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4663 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4665 = _T_4663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4667 = _T_4665 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4668 = _T_4662 | _T_4667; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4678 = _T_3717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4679 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4681 = _T_4679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4683 = _T_4681 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4684 = _T_4678 | _T_4683; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4694 = _T_3721 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4695 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4697 = _T_4695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4699 = _T_4697 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4700 = _T_4694 | _T_4699; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4710 = _T_3725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4711 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4713 = _T_4711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4715 = _T_4713 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4716 = _T_4710 | _T_4715; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4726 = _T_3729 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4727 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4729 = _T_4727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4731 = _T_4729 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4732 = _T_4726 | _T_4731; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4742 = _T_3733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4743 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4745 = _T_4743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4747 = _T_4745 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4748 = _T_4742 | _T_4747; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4758 = _T_3737 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4759 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4761 = _T_4759 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4763 = _T_4761 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4764 = _T_4758 | _T_4763; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4774 = _T_3741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4775 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4777 = _T_4775 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4779 = _T_4777 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4780 = _T_4774 | _T_4779; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4790 = _T_3745 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4791 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4793 = _T_4791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4795 = _T_4793 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4796 = _T_4790 | _T_4795; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4806 = _T_3749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4807 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4809 = _T_4807 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4811 = _T_4809 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4812 = _T_4806 | _T_4811; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4822 = _T_3753 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4823 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4825 = _T_4823 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4827 = _T_4825 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4828 = _T_4822 | _T_4827; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4838 = _T_3757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4839 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4841 = _T_4839 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4843 = _T_4841 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4844 = _T_4838 | _T_4843; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4854 = _T_3761 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4855 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4857 = _T_4855 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4859 = _T_4857 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4860 = _T_4854 | _T_4859; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4870 = _T_3765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4871 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4873 = _T_4871 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4875 = _T_4873 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4876 = _T_4870 | _T_4875; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4886 = _T_3641 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4889 = _T_4375 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4891 = _T_4889 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4892 = _T_4886 | _T_4891; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4902 = _T_3645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4905 = _T_4391 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4907 = _T_4905 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4908 = _T_4902 | _T_4907; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4918 = _T_3649 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4921 = _T_4407 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4923 = _T_4921 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4924 = _T_4918 | _T_4923; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4934 = _T_3653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4937 = _T_4423 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4939 = _T_4937 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4940 = _T_4934 | _T_4939; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4950 = _T_3657 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4953 = _T_4439 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4955 = _T_4953 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4956 = _T_4950 | _T_4955; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4966 = _T_3661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4969 = _T_4455 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4971 = _T_4969 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4972 = _T_4966 | _T_4971; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4982 = _T_3665 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4985 = _T_4471 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4987 = _T_4985 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4988 = _T_4982 | _T_4987; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4998 = _T_3669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5001 = _T_4487 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5003 = _T_5001 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5004 = _T_4998 | _T_5003; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5014 = _T_3673 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5017 = _T_4503 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5019 = _T_5017 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5020 = _T_5014 | _T_5019; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5030 = _T_3677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5033 = _T_4519 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5035 = _T_5033 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5036 = _T_5030 | _T_5035; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5046 = _T_3681 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5049 = _T_4535 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5051 = _T_5049 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5052 = _T_5046 | _T_5051; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5062 = _T_3685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5065 = _T_4551 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5067 = _T_5065 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5068 = _T_5062 | _T_5067; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5078 = _T_3689 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5081 = _T_4567 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5083 = _T_5081 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5084 = _T_5078 | _T_5083; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5094 = _T_3693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5097 = _T_4583 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5099 = _T_5097 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5100 = _T_5094 | _T_5099; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5110 = _T_3697 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5113 = _T_4599 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5115 = _T_5113 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5116 = _T_5110 | _T_5115; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5126 = _T_3701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5129 = _T_4615 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5131 = _T_5129 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5132 = _T_5126 | _T_5131; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5142 = _T_3705 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5145 = _T_4631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5147 = _T_5145 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5148 = _T_5142 | _T_5147; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5158 = _T_3709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5161 = _T_4647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5163 = _T_5161 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5164 = _T_5158 | _T_5163; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5174 = _T_3713 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5177 = _T_4663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5179 = _T_5177 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5180 = _T_5174 | _T_5179; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5190 = _T_3717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5193 = _T_4679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5195 = _T_5193 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5196 = _T_5190 | _T_5195; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5206 = _T_3721 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5209 = _T_4695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5211 = _T_5209 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5212 = _T_5206 | _T_5211; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5222 = _T_3725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5225 = _T_4711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5227 = _T_5225 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5228 = _T_5222 | _T_5227; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5238 = _T_3729 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5241 = _T_4727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5243 = _T_5241 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5244 = _T_5238 | _T_5243; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5254 = _T_3733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5257 = _T_4743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5259 = _T_5257 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5260 = _T_5254 | _T_5259; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5270 = _T_3737 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5273 = _T_4759 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5275 = _T_5273 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5276 = _T_5270 | _T_5275; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5286 = _T_3741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5289 = _T_4775 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5291 = _T_5289 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5292 = _T_5286 | _T_5291; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5302 = _T_3745 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5305 = _T_4791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5307 = _T_5305 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5308 = _T_5302 | _T_5307; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5318 = _T_3749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5321 = _T_4807 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5323 = _T_5321 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5324 = _T_5318 | _T_5323; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5334 = _T_3753 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5337 = _T_4823 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5339 = _T_5337 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5340 = _T_5334 | _T_5339; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5350 = _T_3757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5353 = _T_4839 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5355 = _T_5353 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5356 = _T_5350 | _T_5355; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5366 = _T_3761 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5369 = _T_4855 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5371 = _T_5369 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5372 = _T_5366 | _T_5371; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5382 = _T_3765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5385 = _T_4871 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5387 = _T_5385 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5388 = _T_5382 | _T_5387; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5398 = _T_3769 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5399 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5401 = _T_5399 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5403 = _T_5401 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5404 = _T_5398 | _T_5403; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5414 = _T_3773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5415 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5417 = _T_5415 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5419 = _T_5417 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5420 = _T_5414 | _T_5419; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5430 = _T_3777 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5431 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5433 = _T_5431 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5435 = _T_5433 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5436 = _T_5430 | _T_5435; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5446 = _T_3781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5447 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5449 = _T_5447 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5451 = _T_5449 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5452 = _T_5446 | _T_5451; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5462 = _T_3785 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5463 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5465 = _T_5463 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5467 = _T_5465 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5468 = _T_5462 | _T_5467; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5478 = _T_3789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5479 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5481 = _T_5479 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5483 = _T_5481 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5484 = _T_5478 | _T_5483; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5494 = _T_3793 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5495 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5497 = _T_5495 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5499 = _T_5497 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5500 = _T_5494 | _T_5499; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5510 = _T_3797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5511 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5513 = _T_5511 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5515 = _T_5513 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5516 = _T_5510 | _T_5515; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5526 = _T_3801 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5527 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5529 = _T_5527 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5531 = _T_5529 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5532 = _T_5526 | _T_5531; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5542 = _T_3805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5543 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5545 = _T_5543 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5547 = _T_5545 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5548 = _T_5542 | _T_5547; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5558 = _T_3809 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5559 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5561 = _T_5559 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5563 = _T_5561 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5564 = _T_5558 | _T_5563; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5574 = _T_3813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5575 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5577 = _T_5575 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5579 = _T_5577 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5580 = _T_5574 | _T_5579; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5590 = _T_3817 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5591 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5593 = _T_5591 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5595 = _T_5593 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5596 = _T_5590 | _T_5595; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5606 = _T_3821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5607 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5609 = _T_5607 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5611 = _T_5609 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5612 = _T_5606 | _T_5611; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5622 = _T_3825 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5623 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5625 = _T_5623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5627 = _T_5625 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5628 = _T_5622 | _T_5627; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5638 = _T_3829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5639 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5641 = _T_5639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5643 = _T_5641 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5644 = _T_5638 | _T_5643; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5654 = _T_3833 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5655 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5657 = _T_5655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5659 = _T_5657 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5660 = _T_5654 | _T_5659; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5670 = _T_3837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5671 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5673 = _T_5671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5675 = _T_5673 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5676 = _T_5670 | _T_5675; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5686 = _T_3841 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5687 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5689 = _T_5687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5691 = _T_5689 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5692 = _T_5686 | _T_5691; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5702 = _T_3845 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5703 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5705 = _T_5703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5707 = _T_5705 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5708 = _T_5702 | _T_5707; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5718 = _T_3849 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5719 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5721 = _T_5719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5723 = _T_5721 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5724 = _T_5718 | _T_5723; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5734 = _T_3853 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5735 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5737 = _T_5735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5739 = _T_5737 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5740 = _T_5734 | _T_5739; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5750 = _T_3857 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5751 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5753 = _T_5751 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5755 = _T_5753 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5756 = _T_5750 | _T_5755; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5766 = _T_3861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5767 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5769 = _T_5767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5771 = _T_5769 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5772 = _T_5766 | _T_5771; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5782 = _T_3865 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5783 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5785 = _T_5783 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5787 = _T_5785 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5788 = _T_5782 | _T_5787; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5798 = _T_3869 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5799 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5801 = _T_5799 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5803 = _T_5801 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5804 = _T_5798 | _T_5803; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5814 = _T_3873 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5815 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5817 = _T_5815 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5819 = _T_5817 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5820 = _T_5814 | _T_5819; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5830 = _T_3877 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5831 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5833 = _T_5831 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5835 = _T_5833 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5836 = _T_5830 | _T_5835; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5846 = _T_3881 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5847 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5849 = _T_5847 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5851 = _T_5849 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5852 = _T_5846 | _T_5851; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5862 = _T_3885 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5863 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5865 = _T_5863 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5867 = _T_5865 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5868 = _T_5862 | _T_5867; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5878 = _T_3889 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5879 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5881 = _T_5879 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5883 = _T_5881 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5884 = _T_5878 | _T_5883; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5894 = _T_3893 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5895 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5897 = _T_5895 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5899 = _T_5897 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5900 = _T_5894 | _T_5899; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5910 = _T_3769 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5913 = _T_5399 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5915 = _T_5913 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5916 = _T_5910 | _T_5915; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5926 = _T_3773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5929 = _T_5415 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5931 = _T_5929 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5932 = _T_5926 | _T_5931; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5942 = _T_3777 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5945 = _T_5431 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5947 = _T_5945 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5948 = _T_5942 | _T_5947; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5958 = _T_3781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5961 = _T_5447 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5963 = _T_5961 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5964 = _T_5958 | _T_5963; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5974 = _T_3785 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5977 = _T_5463 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5979 = _T_5977 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5980 = _T_5974 | _T_5979; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5990 = _T_3789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5993 = _T_5479 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5995 = _T_5993 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5996 = _T_5990 | _T_5995; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6006 = _T_3793 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6009 = _T_5495 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6011 = _T_6009 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6012 = _T_6006 | _T_6011; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6022 = _T_3797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6025 = _T_5511 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6027 = _T_6025 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6028 = _T_6022 | _T_6027; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6038 = _T_3801 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6041 = _T_5527 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6043 = _T_6041 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6044 = _T_6038 | _T_6043; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6054 = _T_3805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6057 = _T_5543 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6059 = _T_6057 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6060 = _T_6054 | _T_6059; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6070 = _T_3809 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6073 = _T_5559 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6075 = _T_6073 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6076 = _T_6070 | _T_6075; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6086 = _T_3813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6089 = _T_5575 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6091 = _T_6089 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6092 = _T_6086 | _T_6091; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6102 = _T_3817 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6105 = _T_5591 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6107 = _T_6105 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6108 = _T_6102 | _T_6107; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6118 = _T_3821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6121 = _T_5607 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6123 = _T_6121 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6124 = _T_6118 | _T_6123; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6134 = _T_3825 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6137 = _T_5623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6139 = _T_6137 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6140 = _T_6134 | _T_6139; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6150 = _T_3829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6153 = _T_5639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6155 = _T_6153 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6156 = _T_6150 | _T_6155; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6166 = _T_3833 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6169 = _T_5655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6171 = _T_6169 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6172 = _T_6166 | _T_6171; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6182 = _T_3837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6185 = _T_5671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6187 = _T_6185 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6188 = _T_6182 | _T_6187; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6198 = _T_3841 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6201 = _T_5687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6203 = _T_6201 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6204 = _T_6198 | _T_6203; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6214 = _T_3845 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6217 = _T_5703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6219 = _T_6217 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6220 = _T_6214 | _T_6219; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6230 = _T_3849 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6233 = _T_5719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6235 = _T_6233 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6236 = _T_6230 | _T_6235; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6246 = _T_3853 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6249 = _T_5735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6251 = _T_6249 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6252 = _T_6246 | _T_6251; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6262 = _T_3857 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6265 = _T_5751 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6267 = _T_6265 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6268 = _T_6262 | _T_6267; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6278 = _T_3861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6281 = _T_5767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6283 = _T_6281 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6284 = _T_6278 | _T_6283; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6294 = _T_3865 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6297 = _T_5783 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6299 = _T_6297 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6300 = _T_6294 | _T_6299; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6310 = _T_3869 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6313 = _T_5799 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6315 = _T_6313 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6316 = _T_6310 | _T_6315; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6326 = _T_3873 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6329 = _T_5815 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6331 = _T_6329 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6332 = _T_6326 | _T_6331; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6342 = _T_3877 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6345 = _T_5831 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6347 = _T_6345 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6348 = _T_6342 | _T_6347; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6358 = _T_3881 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6361 = _T_5847 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6363 = _T_6361 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6364 = _T_6358 | _T_6363; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6374 = _T_3885 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6377 = _T_5863 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6379 = _T_6377 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6380 = _T_6374 | _T_6379; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6390 = _T_3889 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6393 = _T_5879 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6395 = _T_6393 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6396 = _T_6390 | _T_6395; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6406 = _T_3893 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6409 = _T_5895 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6411 = _T_6409 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6412 = _T_6406 | _T_6411; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6422 = _T_3897 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6423 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6425 = _T_6423 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6427 = _T_6425 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6428 = _T_6422 | _T_6427; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6438 = _T_3901 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6439 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6441 = _T_6439 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6443 = _T_6441 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6444 = _T_6438 | _T_6443; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6454 = _T_3905 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6455 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6457 = _T_6455 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6459 = _T_6457 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6460 = _T_6454 | _T_6459; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6470 = _T_3909 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6471 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6473 = _T_6471 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6475 = _T_6473 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6476 = _T_6470 | _T_6475; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6486 = _T_3913 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6487 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6489 = _T_6487 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6491 = _T_6489 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6492 = _T_6486 | _T_6491; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6502 = _T_3917 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6503 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6505 = _T_6503 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6507 = _T_6505 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6508 = _T_6502 | _T_6507; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6518 = _T_3921 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6519 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6521 = _T_6519 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6523 = _T_6521 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6524 = _T_6518 | _T_6523; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6534 = _T_3925 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6535 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6537 = _T_6535 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6539 = _T_6537 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6540 = _T_6534 | _T_6539; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6550 = _T_3929 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6551 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6553 = _T_6551 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6555 = _T_6553 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6556 = _T_6550 | _T_6555; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6566 = _T_3933 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6567 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6569 = _T_6567 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6571 = _T_6569 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6572 = _T_6566 | _T_6571; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6582 = _T_3937 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6583 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6585 = _T_6583 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6587 = _T_6585 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6588 = _T_6582 | _T_6587; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6598 = _T_3941 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6599 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6601 = _T_6599 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6603 = _T_6601 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6604 = _T_6598 | _T_6603; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6614 = _T_3945 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6615 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6617 = _T_6615 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6619 = _T_6617 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6620 = _T_6614 | _T_6619; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6630 = _T_3949 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6631 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6633 = _T_6631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6635 = _T_6633 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6636 = _T_6630 | _T_6635; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6646 = _T_3953 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6647 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6649 = _T_6647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6651 = _T_6649 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6652 = _T_6646 | _T_6651; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6662 = _T_3957 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6663 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6665 = _T_6663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6667 = _T_6665 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6668 = _T_6662 | _T_6667; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6678 = _T_3961 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6679 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6681 = _T_6679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6683 = _T_6681 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6684 = _T_6678 | _T_6683; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6694 = _T_3965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6695 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6697 = _T_6695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6699 = _T_6697 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6700 = _T_6694 | _T_6699; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6710 = _T_3969 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6711 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6713 = _T_6711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6715 = _T_6713 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6716 = _T_6710 | _T_6715; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6726 = _T_3973 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6727 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6729 = _T_6727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6731 = _T_6729 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6732 = _T_6726 | _T_6731; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6742 = _T_3977 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6743 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6745 = _T_6743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6747 = _T_6745 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6748 = _T_6742 | _T_6747; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6758 = _T_3981 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6759 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6761 = _T_6759 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6763 = _T_6761 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6764 = _T_6758 | _T_6763; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6774 = _T_3985 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6775 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6777 = _T_6775 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6779 = _T_6777 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6780 = _T_6774 | _T_6779; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6790 = _T_3989 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6791 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6793 = _T_6791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6795 = _T_6793 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6796 = _T_6790 | _T_6795; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6806 = _T_3993 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6807 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6809 = _T_6807 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6811 = _T_6809 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6812 = _T_6806 | _T_6811; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6822 = _T_3997 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6823 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6825 = _T_6823 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6827 = _T_6825 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6828 = _T_6822 | _T_6827; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6838 = _T_4001 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6839 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6841 = _T_6839 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6843 = _T_6841 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6844 = _T_6838 | _T_6843; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6854 = _T_4005 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6855 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6857 = _T_6855 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6859 = _T_6857 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6860 = _T_6854 | _T_6859; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6870 = _T_4009 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6871 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6873 = _T_6871 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6875 = _T_6873 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6876 = _T_6870 | _T_6875; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6886 = _T_4013 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6887 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6889 = _T_6887 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6891 = _T_6889 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6892 = _T_6886 | _T_6891; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6902 = _T_4017 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6903 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6905 = _T_6903 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6907 = _T_6905 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6908 = _T_6902 | _T_6907; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6918 = _T_4021 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6919 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6921 = _T_6919 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6923 = _T_6921 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6924 = _T_6918 | _T_6923; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6934 = _T_3897 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6937 = _T_6423 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6939 = _T_6937 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6940 = _T_6934 | _T_6939; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6950 = _T_3901 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6953 = _T_6439 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6955 = _T_6953 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6956 = _T_6950 | _T_6955; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6966 = _T_3905 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6969 = _T_6455 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6971 = _T_6969 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6972 = _T_6966 | _T_6971; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6982 = _T_3909 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6985 = _T_6471 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6987 = _T_6985 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6988 = _T_6982 | _T_6987; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6998 = _T_3913 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7001 = _T_6487 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7003 = _T_7001 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7004 = _T_6998 | _T_7003; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7014 = _T_3917 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7017 = _T_6503 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7019 = _T_7017 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7020 = _T_7014 | _T_7019; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7030 = _T_3921 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7033 = _T_6519 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7035 = _T_7033 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7036 = _T_7030 | _T_7035; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7046 = _T_3925 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7049 = _T_6535 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7051 = _T_7049 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7052 = _T_7046 | _T_7051; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7062 = _T_3929 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7065 = _T_6551 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7067 = _T_7065 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7068 = _T_7062 | _T_7067; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7078 = _T_3933 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7081 = _T_6567 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7083 = _T_7081 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7084 = _T_7078 | _T_7083; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7094 = _T_3937 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7097 = _T_6583 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7099 = _T_7097 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7100 = _T_7094 | _T_7099; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7110 = _T_3941 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7113 = _T_6599 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7115 = _T_7113 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7116 = _T_7110 | _T_7115; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7126 = _T_3945 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7129 = _T_6615 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7131 = _T_7129 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7132 = _T_7126 | _T_7131; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7142 = _T_3949 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7145 = _T_6631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7147 = _T_7145 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7148 = _T_7142 | _T_7147; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7158 = _T_3953 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7161 = _T_6647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7163 = _T_7161 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7164 = _T_7158 | _T_7163; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7174 = _T_3957 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7177 = _T_6663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7179 = _T_7177 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7180 = _T_7174 | _T_7179; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7190 = _T_3961 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7193 = _T_6679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7195 = _T_7193 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7196 = _T_7190 | _T_7195; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7206 = _T_3965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7209 = _T_6695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7211 = _T_7209 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7212 = _T_7206 | _T_7211; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7222 = _T_3969 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7225 = _T_6711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7227 = _T_7225 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7228 = _T_7222 | _T_7227; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7238 = _T_3973 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7241 = _T_6727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7243 = _T_7241 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7244 = _T_7238 | _T_7243; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7254 = _T_3977 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7257 = _T_6743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7259 = _T_7257 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7260 = _T_7254 | _T_7259; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7270 = _T_3981 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7273 = _T_6759 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7275 = _T_7273 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7276 = _T_7270 | _T_7275; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7286 = _T_3985 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7289 = _T_6775 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7291 = _T_7289 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7292 = _T_7286 | _T_7291; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7302 = _T_3989 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7305 = _T_6791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7307 = _T_7305 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7308 = _T_7302 | _T_7307; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7318 = _T_3993 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7321 = _T_6807 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7323 = _T_7321 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7324 = _T_7318 | _T_7323; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7334 = _T_3997 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7337 = _T_6823 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7339 = _T_7337 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7340 = _T_7334 | _T_7339; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7350 = _T_4001 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7353 = _T_6839 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7355 = _T_7353 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7356 = _T_7350 | _T_7355; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7366 = _T_4005 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7369 = _T_6855 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7371 = _T_7369 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7372 = _T_7366 | _T_7371; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7382 = _T_4009 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7385 = _T_6871 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7387 = _T_7385 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7388 = _T_7382 | _T_7387; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7398 = _T_4013 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7401 = _T_6887 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7403 = _T_7401 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7404 = _T_7398 | _T_7403; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7414 = _T_4017 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7417 = _T_6903 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7419 = _T_7417 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7420 = _T_7414 | _T_7419; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7430 = _T_4021 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7433 = _T_6919 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7435 = _T_7433 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7436 = _T_7430 | _T_7435; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7446 = _T_4025 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7447 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7449 = _T_7447 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7451 = _T_7449 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7452 = _T_7446 | _T_7451; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7462 = _T_4029 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7463 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7465 = _T_7463 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7467 = _T_7465 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7468 = _T_7462 | _T_7467; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7478 = _T_4033 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7479 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7481 = _T_7479 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7483 = _T_7481 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7484 = _T_7478 | _T_7483; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7494 = _T_4037 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7495 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7497 = _T_7495 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7499 = _T_7497 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7500 = _T_7494 | _T_7499; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7510 = _T_4041 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7511 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7513 = _T_7511 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7515 = _T_7513 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7516 = _T_7510 | _T_7515; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7526 = _T_4045 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7527 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7529 = _T_7527 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7531 = _T_7529 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7532 = _T_7526 | _T_7531; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7542 = _T_4049 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7543 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7545 = _T_7543 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7547 = _T_7545 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7548 = _T_7542 | _T_7547; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7558 = _T_4053 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7559 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7561 = _T_7559 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7563 = _T_7561 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7564 = _T_7558 | _T_7563; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7574 = _T_4057 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7575 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7577 = _T_7575 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7579 = _T_7577 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7580 = _T_7574 | _T_7579; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7590 = _T_4061 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7591 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7593 = _T_7591 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7595 = _T_7593 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7596 = _T_7590 | _T_7595; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7606 = _T_4065 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7607 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7609 = _T_7607 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7611 = _T_7609 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7612 = _T_7606 | _T_7611; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7622 = _T_4069 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7623 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7625 = _T_7623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7627 = _T_7625 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7628 = _T_7622 | _T_7627; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7638 = _T_4073 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7639 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7641 = _T_7639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7643 = _T_7641 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7644 = _T_7638 | _T_7643; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7654 = _T_4077 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7655 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7657 = _T_7655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7659 = _T_7657 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7660 = _T_7654 | _T_7659; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7670 = _T_4081 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7671 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7673 = _T_7671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7675 = _T_7673 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7676 = _T_7670 | _T_7675; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7686 = _T_4085 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7687 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7689 = _T_7687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7691 = _T_7689 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7692 = _T_7686 | _T_7691; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7702 = _T_4089 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7703 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7705 = _T_7703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7707 = _T_7705 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7708 = _T_7702 | _T_7707; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7718 = _T_4093 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7719 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7721 = _T_7719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7723 = _T_7721 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7724 = _T_7718 | _T_7723; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7734 = _T_4097 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7735 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7737 = _T_7735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7739 = _T_7737 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7740 = _T_7734 | _T_7739; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7750 = _T_4101 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7751 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7753 = _T_7751 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7755 = _T_7753 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7756 = _T_7750 | _T_7755; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7766 = _T_4105 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7767 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7769 = _T_7767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7771 = _T_7769 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7772 = _T_7766 | _T_7771; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7782 = _T_4109 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7783 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7785 = _T_7783 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7787 = _T_7785 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7788 = _T_7782 | _T_7787; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7798 = _T_4113 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7799 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7801 = _T_7799 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7803 = _T_7801 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7804 = _T_7798 | _T_7803; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7814 = _T_4117 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7815 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7817 = _T_7815 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7819 = _T_7817 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7820 = _T_7814 | _T_7819; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7830 = _T_4121 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7831 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7833 = _T_7831 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7835 = _T_7833 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7836 = _T_7830 | _T_7835; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7846 = _T_4125 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7847 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7849 = _T_7847 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7851 = _T_7849 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7852 = _T_7846 | _T_7851; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7862 = _T_4129 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7863 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7865 = _T_7863 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7867 = _T_7865 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7868 = _T_7862 | _T_7867; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7878 = _T_4133 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7879 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7881 = _T_7879 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7883 = _T_7881 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7884 = _T_7878 | _T_7883; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7894 = _T_4137 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7895 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7897 = _T_7895 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7899 = _T_7897 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7900 = _T_7894 | _T_7899; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7910 = _T_4141 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7911 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7913 = _T_7911 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7915 = _T_7913 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7916 = _T_7910 | _T_7915; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7926 = _T_4145 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7927 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7929 = _T_7927 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7931 = _T_7929 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7932 = _T_7926 | _T_7931; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7942 = _T_4149 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7943 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7945 = _T_7943 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7947 = _T_7945 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7948 = _T_7942 | _T_7947; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7958 = _T_4025 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7961 = _T_7447 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7963 = _T_7961 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7964 = _T_7958 | _T_7963; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7974 = _T_4029 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7977 = _T_7463 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7979 = _T_7977 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7980 = _T_7974 | _T_7979; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7990 = _T_4033 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7993 = _T_7479 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7995 = _T_7993 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7996 = _T_7990 | _T_7995; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8006 = _T_4037 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8009 = _T_7495 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8011 = _T_8009 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8012 = _T_8006 | _T_8011; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8022 = _T_4041 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8025 = _T_7511 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8027 = _T_8025 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8028 = _T_8022 | _T_8027; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8038 = _T_4045 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8041 = _T_7527 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8043 = _T_8041 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8044 = _T_8038 | _T_8043; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8054 = _T_4049 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8057 = _T_7543 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8059 = _T_8057 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8060 = _T_8054 | _T_8059; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8070 = _T_4053 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8073 = _T_7559 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8075 = _T_8073 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8076 = _T_8070 | _T_8075; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8086 = _T_4057 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8089 = _T_7575 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8091 = _T_8089 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8092 = _T_8086 | _T_8091; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8102 = _T_4061 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8105 = _T_7591 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8107 = _T_8105 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8108 = _T_8102 | _T_8107; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8118 = _T_4065 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8121 = _T_7607 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8123 = _T_8121 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8124 = _T_8118 | _T_8123; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8134 = _T_4069 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8137 = _T_7623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8139 = _T_8137 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8140 = _T_8134 | _T_8139; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8150 = _T_4073 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8153 = _T_7639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8155 = _T_8153 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8156 = _T_8150 | _T_8155; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8166 = _T_4077 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8169 = _T_7655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8171 = _T_8169 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8172 = _T_8166 | _T_8171; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8182 = _T_4081 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8185 = _T_7671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8187 = _T_8185 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8188 = _T_8182 | _T_8187; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8198 = _T_4085 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8201 = _T_7687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8203 = _T_8201 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8204 = _T_8198 | _T_8203; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8214 = _T_4089 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8217 = _T_7703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8219 = _T_8217 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8220 = _T_8214 | _T_8219; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8230 = _T_4093 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8233 = _T_7719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8235 = _T_8233 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8236 = _T_8230 | _T_8235; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8246 = _T_4097 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8249 = _T_7735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8251 = _T_8249 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8252 = _T_8246 | _T_8251; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8262 = _T_4101 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8265 = _T_7751 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8267 = _T_8265 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8268 = _T_8262 | _T_8267; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8278 = _T_4105 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8281 = _T_7767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8283 = _T_8281 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8284 = _T_8278 | _T_8283; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8294 = _T_4109 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8297 = _T_7783 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8299 = _T_8297 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8300 = _T_8294 | _T_8299; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8310 = _T_4113 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8313 = _T_7799 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8315 = _T_8313 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8316 = _T_8310 | _T_8315; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8326 = _T_4117 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8329 = _T_7815 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8331 = _T_8329 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8332 = _T_8326 | _T_8331; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8342 = _T_4121 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8345 = _T_7831 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8347 = _T_8345 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8348 = _T_8342 | _T_8347; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8358 = _T_4125 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8361 = _T_7847 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8363 = _T_8361 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8364 = _T_8358 | _T_8363; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8374 = _T_4129 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8377 = _T_7863 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8379 = _T_8377 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8380 = _T_8374 | _T_8379; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8390 = _T_4133 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8393 = _T_7879 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8395 = _T_8393 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8396 = _T_8390 | _T_8395; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8406 = _T_4137 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8409 = _T_7895 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8411 = _T_8409 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8412 = _T_8406 | _T_8411; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8422 = _T_4141 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8425 = _T_7911 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8427 = _T_8425 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8428 = _T_8422 | _T_8427; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8438 = _T_4145 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8441 = _T_7927 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8443 = _T_8441 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8444 = _T_8438 | _T_8443; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8454 = _T_4149 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8457 = _T_7943 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8459 = _T_8457 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8460 = _T_8454 | _T_8459; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_9261 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 811:63]
  wire  _T_9262 = _T_9261 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 811:85]
  wire [1:0] _T_9264 = _T_9262 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9271; // @[el2_ifu_mem_ctl.scala 816:57]
  reg  _T_9272; // @[el2_ifu_mem_ctl.scala 817:56]
  reg  _T_9273; // @[el2_ifu_mem_ctl.scala 818:59]
  wire  _T_9274 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 819:80]
  wire  _T_9275 = ifu_bus_arvalid_ff & _T_9274; // @[el2_ifu_mem_ctl.scala 819:78]
  wire  _T_9276 = _T_9275 & miss_pending; // @[el2_ifu_mem_ctl.scala 819:100]
  reg  _T_9277; // @[el2_ifu_mem_ctl.scala 819:58]
  reg  _T_9278; // @[el2_ifu_mem_ctl.scala 820:58]
  wire  _T_9281 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 827:71]
  wire  _T_9283 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 827:124]
  wire  _T_9285 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 828:50]
  wire  _T_9287 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 828:103]
  wire [3:0] _T_9290 = {_T_9281,_T_9283,_T_9285,_T_9287}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 830:53]
  reg  _T_9301; // @[Reg.scala 27:20]
  rvecc_encode_64 m1 ( // @[el2_ifu_mem_ctl.scala 343:18]
    .io_din(m1_io_din),
    .io_ecc_out(m1_io_ecc_out)
  );
  rvecc_encode_64 m2 ( // @[el2_ifu_mem_ctl.scala 344:18]
    .io_din(m2_io_din),
    .io_ecc_out(m2_io_ecc_out)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 329:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 328:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 192:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3096; // @[el2_ifu_mem_ctl.scala 707:21]
  assign io_ifu_pmu_ic_miss = _T_9271; // @[el2_ifu_mem_ctl.scala 816:22]
  assign io_ifu_pmu_ic_hit = _T_9272; // @[el2_ifu_mem_ctl.scala 817:21]
  assign io_ifu_pmu_bus_error = _T_9273; // @[el2_ifu_mem_ctl.scala 818:24]
  assign io_ifu_pmu_bus_busy = _T_9277; // @[el2_ifu_mem_ctl.scala 819:23]
  assign io_ifu_pmu_bus_trxn = _T_9278; // @[el2_ifu_mem_ctl.scala 820:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 143:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 142:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 141:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 152:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 145:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 136:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 134:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 135:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 153:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 569:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_1690; // @[el2_ifu_mem_ctl.scala 570:19]
  assign io_ifu_axi_araddr = _T_1692 & _T_1694; // @[el2_ifu_mem_ctl.scala 571:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 574:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 149:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 572:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 575:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 573:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 151:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 146:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 576:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 666:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 664:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 668:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 659:20]
  assign io_iccm_ready = _T_1793 & _T_1787; // @[el2_ifu_mem_ctl.scala 639:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 338:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 706:15]
  assign io_ic_rd_en = _T_3074 | _T_3079; // @[el2_ifu_mem_ctl.scala 697:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 353:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 353:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 354:23]
  assign io_ifu_ic_debug_rd_data = _T_365; // @[el2_ifu_mem_ctl.scala 362:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 823:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 825:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 826:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 824:25]
  assign io_ic_debug_way = _T_9290[1:0]; // @[el2_ifu_mem_ctl.scala 827:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9264; // @[el2_ifu_mem_ctl.scala 811:19]
  assign io_iccm_rw_addr = _T_2228[14:0]; // @[el2_ifu_mem_ctl.scala 670:19]
  assign io_iccm_wren = _T_1797 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 641:16]
  assign io_iccm_rden = _T_1801 | _T_1802; // @[el2_ifu_mem_ctl.scala 642:16]
  assign io_iccm_wr_data = _T_2203 ? _T_2204 : _T_2211; // @[el2_ifu_mem_ctl.scala 647:19]
  assign io_iccm_wr_size = _T_1807 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 644:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 290:15]
  assign io_ic_access_fault_f = _T_1575 & _T_317; // @[el2_ifu_mem_ctl.scala 395:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_429; // @[el2_ifu_mem_ctl.scala 396:29]
  assign io_iccm_rd_ecc_single_err = _T_3019 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 683:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 684:29]
  assign io_ic_error_start = _T_353 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 356:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 190:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 400:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 392:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 389:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 390:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9301; // @[el2_ifu_mem_ctl.scala 834:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_1580; // @[el2_ifu_mem_ctl.scala 488:27]
  assign io_iccm_correction_state = _T_1608 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 523:28 el2_ifu_mem_ctl.scala 536:32 el2_ifu_mem_ctl.scala 543:32 el2_ifu_mem_ctl.scala 550:32]
  assign io_ic_miss_buff_ecc = m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 351:23]
  assign io_ic_wr_ecc = m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 347:16]
  assign m1_io_din = ifu_bus_rdata_ff; // @[el2_ifu_mem_ctl.scala 345:13]
  assign m2_io_din = {_T_1531,_T_1571}; // @[el2_ifu_mem_ctl.scala 349:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4284 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_3640 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_3636 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_3632 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_3628 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_3624 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_3620 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_3616 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_3612 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_3608 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_3604 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_3600 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_3596 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_3592 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_3588 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_3584 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_3580 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_3576 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_3572 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_3568 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_3564 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_3560 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_3556 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_3552 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_3548 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_3544 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_3540 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_3536 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_3532 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_3528 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_3524 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_3520 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_3516 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_3512 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_3508 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_3504 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_3500 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_3496 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_3492 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_3488 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_3484 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_3480 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_3476 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_3472 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_3468 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_3464 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_3460 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_3456 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_3452 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_3448 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_3444 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_3440 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_3436 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_3432 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_3428 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_3424 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_3420 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_3416 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_3412 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_3408 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_3404 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_3400 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_3396 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_3392 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_3388 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_3384 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_3380 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_3376 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_3372 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_3368 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_3364 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_3360 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_3356 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_3352 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_3348 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_3344 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_3340 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_3336 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_3332 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_3328 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_3324 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_3320 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_3316 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_3312 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_3308 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_3304 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_3300 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_3296 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_3292 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_3288 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_3284 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_3280 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_3276 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_3272 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_3268 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_3264 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_3260 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_3256 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_3252 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_3248 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_3244 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_3240 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_3236 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_3232 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_3228 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_3224 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_3220 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_3216 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_3212 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_3208 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_3204 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_3200 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_3196 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_3192 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3188 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3184 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3180 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3176 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3172 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3168 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3164 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3160 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3156 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3152 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3148 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3144 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3140 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3136 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3132 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_365 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_9271 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_9272 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_9273 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_9277 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9278 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9301 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_3640 <= 3'h0;
    end else if (_T_3639) begin
      _T_3640 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3636 <= 3'h0;
    end else if (_T_3635) begin
      _T_3636 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3632 <= 3'h0;
    end else if (_T_3631) begin
      _T_3632 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3628 <= 3'h0;
    end else if (_T_3627) begin
      _T_3628 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3624 <= 3'h0;
    end else if (_T_3623) begin
      _T_3624 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3620 <= 3'h0;
    end else if (_T_3619) begin
      _T_3620 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3616 <= 3'h0;
    end else if (_T_3615) begin
      _T_3616 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3612 <= 3'h0;
    end else if (_T_3611) begin
      _T_3612 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3608 <= 3'h0;
    end else if (_T_3607) begin
      _T_3608 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3604 <= 3'h0;
    end else if (_T_3603) begin
      _T_3604 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3600 <= 3'h0;
    end else if (_T_3599) begin
      _T_3600 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3596 <= 3'h0;
    end else if (_T_3595) begin
      _T_3596 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3592 <= 3'h0;
    end else if (_T_3591) begin
      _T_3592 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3588 <= 3'h0;
    end else if (_T_3587) begin
      _T_3588 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3584 <= 3'h0;
    end else if (_T_3583) begin
      _T_3584 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3580 <= 3'h0;
    end else if (_T_3579) begin
      _T_3580 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3576 <= 3'h0;
    end else if (_T_3575) begin
      _T_3576 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3572 <= 3'h0;
    end else if (_T_3571) begin
      _T_3572 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3568 <= 3'h0;
    end else if (_T_3567) begin
      _T_3568 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3564 <= 3'h0;
    end else if (_T_3563) begin
      _T_3564 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3560 <= 3'h0;
    end else if (_T_3559) begin
      _T_3560 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3556 <= 3'h0;
    end else if (_T_3555) begin
      _T_3556 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3552 <= 3'h0;
    end else if (_T_3551) begin
      _T_3552 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3548 <= 3'h0;
    end else if (_T_3547) begin
      _T_3548 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3544 <= 3'h0;
    end else if (_T_3543) begin
      _T_3544 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3540 <= 3'h0;
    end else if (_T_3539) begin
      _T_3540 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3536 <= 3'h0;
    end else if (_T_3535) begin
      _T_3536 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3532 <= 3'h0;
    end else if (_T_3531) begin
      _T_3532 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3528 <= 3'h0;
    end else if (_T_3527) begin
      _T_3528 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3524 <= 3'h0;
    end else if (_T_3523) begin
      _T_3524 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3520 <= 3'h0;
    end else if (_T_3519) begin
      _T_3520 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3516 <= 3'h0;
    end else if (_T_3515) begin
      _T_3516 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3512 <= 3'h0;
    end else if (_T_3511) begin
      _T_3512 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3508 <= 3'h0;
    end else if (_T_3507) begin
      _T_3508 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3504 <= 3'h0;
    end else if (_T_3503) begin
      _T_3504 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3500 <= 3'h0;
    end else if (_T_3499) begin
      _T_3500 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3496 <= 3'h0;
    end else if (_T_3495) begin
      _T_3496 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3492 <= 3'h0;
    end else if (_T_3491) begin
      _T_3492 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3488 <= 3'h0;
    end else if (_T_3487) begin
      _T_3488 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3484 <= 3'h0;
    end else if (_T_3483) begin
      _T_3484 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3480 <= 3'h0;
    end else if (_T_3479) begin
      _T_3480 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3476 <= 3'h0;
    end else if (_T_3475) begin
      _T_3476 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3472 <= 3'h0;
    end else if (_T_3471) begin
      _T_3472 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3468 <= 3'h0;
    end else if (_T_3467) begin
      _T_3468 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3464 <= 3'h0;
    end else if (_T_3463) begin
      _T_3464 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3460 <= 3'h0;
    end else if (_T_3459) begin
      _T_3460 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3456 <= 3'h0;
    end else if (_T_3455) begin
      _T_3456 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3452 <= 3'h0;
    end else if (_T_3451) begin
      _T_3452 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3448 <= 3'h0;
    end else if (_T_3447) begin
      _T_3448 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3444 <= 3'h0;
    end else if (_T_3443) begin
      _T_3444 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3440 <= 3'h0;
    end else if (_T_3439) begin
      _T_3440 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3436 <= 3'h0;
    end else if (_T_3435) begin
      _T_3436 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3432 <= 3'h0;
    end else if (_T_3431) begin
      _T_3432 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3428 <= 3'h0;
    end else if (_T_3427) begin
      _T_3428 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3424 <= 3'h0;
    end else if (_T_3423) begin
      _T_3424 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3420 <= 3'h0;
    end else if (_T_3419) begin
      _T_3420 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3416 <= 3'h0;
    end else if (_T_3415) begin
      _T_3416 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3412 <= 3'h0;
    end else if (_T_3411) begin
      _T_3412 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3408 <= 3'h0;
    end else if (_T_3407) begin
      _T_3408 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3404 <= 3'h0;
    end else if (_T_3403) begin
      _T_3404 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3400 <= 3'h0;
    end else if (_T_3399) begin
      _T_3400 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3396 <= 3'h0;
    end else if (_T_3395) begin
      _T_3396 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3392 <= 3'h0;
    end else if (_T_3391) begin
      _T_3392 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3388 <= 3'h0;
    end else if (_T_3387) begin
      _T_3388 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3384 <= 3'h0;
    end else if (_T_3383) begin
      _T_3384 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3380 <= 3'h0;
    end else if (_T_3379) begin
      _T_3380 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3376 <= 3'h0;
    end else if (_T_3375) begin
      _T_3376 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3372 <= 3'h0;
    end else if (_T_3371) begin
      _T_3372 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3368 <= 3'h0;
    end else if (_T_3367) begin
      _T_3368 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3364 <= 3'h0;
    end else if (_T_3363) begin
      _T_3364 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3360 <= 3'h0;
    end else if (_T_3359) begin
      _T_3360 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3356 <= 3'h0;
    end else if (_T_3355) begin
      _T_3356 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3352 <= 3'h0;
    end else if (_T_3351) begin
      _T_3352 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3348 <= 3'h0;
    end else if (_T_3347) begin
      _T_3348 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3344 <= 3'h0;
    end else if (_T_3343) begin
      _T_3344 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3340 <= 3'h0;
    end else if (_T_3339) begin
      _T_3340 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3336 <= 3'h0;
    end else if (_T_3335) begin
      _T_3336 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3332 <= 3'h0;
    end else if (_T_3331) begin
      _T_3332 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3328 <= 3'h0;
    end else if (_T_3327) begin
      _T_3328 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3324 <= 3'h0;
    end else if (_T_3323) begin
      _T_3324 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3320 <= 3'h0;
    end else if (_T_3319) begin
      _T_3320 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3316 <= 3'h0;
    end else if (_T_3315) begin
      _T_3316 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3312 <= 3'h0;
    end else if (_T_3311) begin
      _T_3312 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3308 <= 3'h0;
    end else if (_T_3307) begin
      _T_3308 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3304 <= 3'h0;
    end else if (_T_3303) begin
      _T_3304 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3300 <= 3'h0;
    end else if (_T_3299) begin
      _T_3300 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3296 <= 3'h0;
    end else if (_T_3295) begin
      _T_3296 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3292 <= 3'h0;
    end else if (_T_3291) begin
      _T_3292 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3288 <= 3'h0;
    end else if (_T_3287) begin
      _T_3288 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3284 <= 3'h0;
    end else if (_T_3283) begin
      _T_3284 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3280 <= 3'h0;
    end else if (_T_3279) begin
      _T_3280 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3276 <= 3'h0;
    end else if (_T_3275) begin
      _T_3276 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3272 <= 3'h0;
    end else if (_T_3271) begin
      _T_3272 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3268 <= 3'h0;
    end else if (_T_3267) begin
      _T_3268 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3264 <= 3'h0;
    end else if (_T_3263) begin
      _T_3264 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3260 <= 3'h0;
    end else if (_T_3259) begin
      _T_3260 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3256 <= 3'h0;
    end else if (_T_3255) begin
      _T_3256 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3252 <= 3'h0;
    end else if (_T_3251) begin
      _T_3252 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3248 <= 3'h0;
    end else if (_T_3247) begin
      _T_3248 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3244 <= 3'h0;
    end else if (_T_3243) begin
      _T_3244 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3240 <= 3'h0;
    end else if (_T_3239) begin
      _T_3240 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3236 <= 3'h0;
    end else if (_T_3235) begin
      _T_3236 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3232 <= 3'h0;
    end else if (_T_3231) begin
      _T_3232 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3228 <= 3'h0;
    end else if (_T_3227) begin
      _T_3228 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3224 <= 3'h0;
    end else if (_T_3223) begin
      _T_3224 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3220 <= 3'h0;
    end else if (_T_3219) begin
      _T_3220 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3216 <= 3'h0;
    end else if (_T_3215) begin
      _T_3216 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3212 <= 3'h0;
    end else if (_T_3211) begin
      _T_3212 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3208 <= 3'h0;
    end else if (_T_3207) begin
      _T_3208 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3204 <= 3'h0;
    end else if (_T_3203) begin
      _T_3204 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3200 <= 3'h0;
    end else if (_T_3199) begin
      _T_3200 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3196 <= 3'h0;
    end else if (_T_3195) begin
      _T_3196 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3192 <= 3'h0;
    end else if (_T_3191) begin
      _T_3192 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3188 <= 3'h0;
    end else if (_T_3187) begin
      _T_3188 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3184 <= 3'h0;
    end else if (_T_3183) begin
      _T_3184 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3180 <= 3'h0;
    end else if (_T_3179) begin
      _T_3180 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3176 <= 3'h0;
    end else if (_T_3175) begin
      _T_3176 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3172 <= 3'h0;
    end else if (_T_3171) begin
      _T_3172 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3168 <= 3'h0;
    end else if (_T_3167) begin
      _T_3168 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3164 <= 3'h0;
    end else if (_T_3163) begin
      _T_3164 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3160 <= 3'h0;
    end else if (_T_3159) begin
      _T_3160 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3156 <= 3'h0;
    end else if (_T_3155) begin
      _T_3156 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3152 <= 3'h0;
    end else if (_T_3151) begin
      _T_3152 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3148 <= 3'h0;
    end else if (_T_3147) begin
      _T_3148 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3144 <= 3'h0;
    end else if (_T_3143) begin
      _T_3144 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3140 <= 3'h0;
    end else if (_T_3139) begin
      _T_3140 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3136 <= 3'h0;
    end else if (_T_3135) begin
      _T_3136 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3132 <= 3'h0;
    end else if (_T_3131) begin
      _T_3132 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_289;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_1733) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_1729;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_4892) begin
      ic_tag_valid_out_1_0 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_4908) begin
      ic_tag_valid_out_1_1 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_4924) begin
      ic_tag_valid_out_1_2 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_4940) begin
      ic_tag_valid_out_1_3 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_4956) begin
      ic_tag_valid_out_1_4 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_4972) begin
      ic_tag_valid_out_1_5 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_4988) begin
      ic_tag_valid_out_1_6 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5004) begin
      ic_tag_valid_out_1_7 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5020) begin
      ic_tag_valid_out_1_8 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5036) begin
      ic_tag_valid_out_1_9 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5052) begin
      ic_tag_valid_out_1_10 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5068) begin
      ic_tag_valid_out_1_11 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5084) begin
      ic_tag_valid_out_1_12 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5100) begin
      ic_tag_valid_out_1_13 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5116) begin
      ic_tag_valid_out_1_14 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5132) begin
      ic_tag_valid_out_1_15 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5148) begin
      ic_tag_valid_out_1_16 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5164) begin
      ic_tag_valid_out_1_17 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5180) begin
      ic_tag_valid_out_1_18 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5196) begin
      ic_tag_valid_out_1_19 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5212) begin
      ic_tag_valid_out_1_20 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5228) begin
      ic_tag_valid_out_1_21 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5244) begin
      ic_tag_valid_out_1_22 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5260) begin
      ic_tag_valid_out_1_23 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5276) begin
      ic_tag_valid_out_1_24 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5292) begin
      ic_tag_valid_out_1_25 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5308) begin
      ic_tag_valid_out_1_26 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5324) begin
      ic_tag_valid_out_1_27 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_5340) begin
      ic_tag_valid_out_1_28 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_5356) begin
      ic_tag_valid_out_1_29 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_5372) begin
      ic_tag_valid_out_1_30 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_5388) begin
      ic_tag_valid_out_1_31 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_5916) begin
      ic_tag_valid_out_1_32 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_5932) begin
      ic_tag_valid_out_1_33 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_5948) begin
      ic_tag_valid_out_1_34 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_5964) begin
      ic_tag_valid_out_1_35 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_5980) begin
      ic_tag_valid_out_1_36 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_5996) begin
      ic_tag_valid_out_1_37 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6012) begin
      ic_tag_valid_out_1_38 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6028) begin
      ic_tag_valid_out_1_39 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6044) begin
      ic_tag_valid_out_1_40 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6060) begin
      ic_tag_valid_out_1_41 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6076) begin
      ic_tag_valid_out_1_42 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6092) begin
      ic_tag_valid_out_1_43 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6108) begin
      ic_tag_valid_out_1_44 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6124) begin
      ic_tag_valid_out_1_45 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6140) begin
      ic_tag_valid_out_1_46 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6156) begin
      ic_tag_valid_out_1_47 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6172) begin
      ic_tag_valid_out_1_48 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6188) begin
      ic_tag_valid_out_1_49 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6204) begin
      ic_tag_valid_out_1_50 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6220) begin
      ic_tag_valid_out_1_51 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6236) begin
      ic_tag_valid_out_1_52 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6252) begin
      ic_tag_valid_out_1_53 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6268) begin
      ic_tag_valid_out_1_54 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6284) begin
      ic_tag_valid_out_1_55 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6300) begin
      ic_tag_valid_out_1_56 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6316) begin
      ic_tag_valid_out_1_57 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6332) begin
      ic_tag_valid_out_1_58 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6348) begin
      ic_tag_valid_out_1_59 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6364) begin
      ic_tag_valid_out_1_60 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6380) begin
      ic_tag_valid_out_1_61 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_6396) begin
      ic_tag_valid_out_1_62 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_6412) begin
      ic_tag_valid_out_1_63 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_6940) begin
      ic_tag_valid_out_1_64 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_6956) begin
      ic_tag_valid_out_1_65 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_6972) begin
      ic_tag_valid_out_1_66 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_6988) begin
      ic_tag_valid_out_1_67 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7004) begin
      ic_tag_valid_out_1_68 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7020) begin
      ic_tag_valid_out_1_69 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7036) begin
      ic_tag_valid_out_1_70 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7052) begin
      ic_tag_valid_out_1_71 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7068) begin
      ic_tag_valid_out_1_72 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7084) begin
      ic_tag_valid_out_1_73 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7100) begin
      ic_tag_valid_out_1_74 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7116) begin
      ic_tag_valid_out_1_75 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7132) begin
      ic_tag_valid_out_1_76 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7148) begin
      ic_tag_valid_out_1_77 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7164) begin
      ic_tag_valid_out_1_78 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7180) begin
      ic_tag_valid_out_1_79 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7196) begin
      ic_tag_valid_out_1_80 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7212) begin
      ic_tag_valid_out_1_81 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7228) begin
      ic_tag_valid_out_1_82 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7244) begin
      ic_tag_valid_out_1_83 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7260) begin
      ic_tag_valid_out_1_84 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7276) begin
      ic_tag_valid_out_1_85 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7292) begin
      ic_tag_valid_out_1_86 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7308) begin
      ic_tag_valid_out_1_87 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7324) begin
      ic_tag_valid_out_1_88 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7340) begin
      ic_tag_valid_out_1_89 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7356) begin
      ic_tag_valid_out_1_90 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7372) begin
      ic_tag_valid_out_1_91 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7388) begin
      ic_tag_valid_out_1_92 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7404) begin
      ic_tag_valid_out_1_93 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7420) begin
      ic_tag_valid_out_1_94 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7436) begin
      ic_tag_valid_out_1_95 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_7964) begin
      ic_tag_valid_out_1_96 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_7980) begin
      ic_tag_valid_out_1_97 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_7996) begin
      ic_tag_valid_out_1_98 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8012) begin
      ic_tag_valid_out_1_99 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8028) begin
      ic_tag_valid_out_1_100 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8044) begin
      ic_tag_valid_out_1_101 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8060) begin
      ic_tag_valid_out_1_102 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8076) begin
      ic_tag_valid_out_1_103 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8092) begin
      ic_tag_valid_out_1_104 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8108) begin
      ic_tag_valid_out_1_105 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8124) begin
      ic_tag_valid_out_1_106 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8140) begin
      ic_tag_valid_out_1_107 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8156) begin
      ic_tag_valid_out_1_108 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8172) begin
      ic_tag_valid_out_1_109 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8188) begin
      ic_tag_valid_out_1_110 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8204) begin
      ic_tag_valid_out_1_111 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8220) begin
      ic_tag_valid_out_1_112 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8236) begin
      ic_tag_valid_out_1_113 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8252) begin
      ic_tag_valid_out_1_114 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8268) begin
      ic_tag_valid_out_1_115 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8284) begin
      ic_tag_valid_out_1_116 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8300) begin
      ic_tag_valid_out_1_117 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8316) begin
      ic_tag_valid_out_1_118 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8332) begin
      ic_tag_valid_out_1_119 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8348) begin
      ic_tag_valid_out_1_120 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8364) begin
      ic_tag_valid_out_1_121 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8380) begin
      ic_tag_valid_out_1_122 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8396) begin
      ic_tag_valid_out_1_123 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8412) begin
      ic_tag_valid_out_1_124 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8428) begin
      ic_tag_valid_out_1_125 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8444) begin
      ic_tag_valid_out_1_126 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8460) begin
      ic_tag_valid_out_1_127 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_4380) begin
      ic_tag_valid_out_0_0 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_4396) begin
      ic_tag_valid_out_0_1 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_4412) begin
      ic_tag_valid_out_0_2 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_4428) begin
      ic_tag_valid_out_0_3 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_4444) begin
      ic_tag_valid_out_0_4 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_4460) begin
      ic_tag_valid_out_0_5 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_4476) begin
      ic_tag_valid_out_0_6 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_4492) begin
      ic_tag_valid_out_0_7 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_4508) begin
      ic_tag_valid_out_0_8 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_4524) begin
      ic_tag_valid_out_0_9 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_4540) begin
      ic_tag_valid_out_0_10 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_4556) begin
      ic_tag_valid_out_0_11 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_4572) begin
      ic_tag_valid_out_0_12 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_4588) begin
      ic_tag_valid_out_0_13 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_4604) begin
      ic_tag_valid_out_0_14 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_4620) begin
      ic_tag_valid_out_0_15 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_4636) begin
      ic_tag_valid_out_0_16 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_4652) begin
      ic_tag_valid_out_0_17 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_4668) begin
      ic_tag_valid_out_0_18 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_4684) begin
      ic_tag_valid_out_0_19 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_4700) begin
      ic_tag_valid_out_0_20 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_4716) begin
      ic_tag_valid_out_0_21 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_4732) begin
      ic_tag_valid_out_0_22 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_4748) begin
      ic_tag_valid_out_0_23 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_4764) begin
      ic_tag_valid_out_0_24 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_4780) begin
      ic_tag_valid_out_0_25 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_4796) begin
      ic_tag_valid_out_0_26 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_4812) begin
      ic_tag_valid_out_0_27 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_4828) begin
      ic_tag_valid_out_0_28 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_4844) begin
      ic_tag_valid_out_0_29 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_4860) begin
      ic_tag_valid_out_0_30 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_4876) begin
      ic_tag_valid_out_0_31 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_5404) begin
      ic_tag_valid_out_0_32 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_5420) begin
      ic_tag_valid_out_0_33 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_5436) begin
      ic_tag_valid_out_0_34 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_5452) begin
      ic_tag_valid_out_0_35 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_5468) begin
      ic_tag_valid_out_0_36 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_5484) begin
      ic_tag_valid_out_0_37 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_5500) begin
      ic_tag_valid_out_0_38 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_5516) begin
      ic_tag_valid_out_0_39 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_5532) begin
      ic_tag_valid_out_0_40 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_5548) begin
      ic_tag_valid_out_0_41 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_5564) begin
      ic_tag_valid_out_0_42 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_5580) begin
      ic_tag_valid_out_0_43 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_5596) begin
      ic_tag_valid_out_0_44 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_5612) begin
      ic_tag_valid_out_0_45 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_5628) begin
      ic_tag_valid_out_0_46 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_5644) begin
      ic_tag_valid_out_0_47 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_5660) begin
      ic_tag_valid_out_0_48 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_5676) begin
      ic_tag_valid_out_0_49 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_5692) begin
      ic_tag_valid_out_0_50 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_5708) begin
      ic_tag_valid_out_0_51 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_5724) begin
      ic_tag_valid_out_0_52 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_5740) begin
      ic_tag_valid_out_0_53 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_5756) begin
      ic_tag_valid_out_0_54 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_5772) begin
      ic_tag_valid_out_0_55 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_5788) begin
      ic_tag_valid_out_0_56 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_5804) begin
      ic_tag_valid_out_0_57 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_5820) begin
      ic_tag_valid_out_0_58 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_5836) begin
      ic_tag_valid_out_0_59 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_5852) begin
      ic_tag_valid_out_0_60 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_5868) begin
      ic_tag_valid_out_0_61 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_5884) begin
      ic_tag_valid_out_0_62 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_5900) begin
      ic_tag_valid_out_0_63 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_6428) begin
      ic_tag_valid_out_0_64 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_6444) begin
      ic_tag_valid_out_0_65 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_6460) begin
      ic_tag_valid_out_0_66 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_6476) begin
      ic_tag_valid_out_0_67 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_6492) begin
      ic_tag_valid_out_0_68 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_6508) begin
      ic_tag_valid_out_0_69 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_6524) begin
      ic_tag_valid_out_0_70 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_6540) begin
      ic_tag_valid_out_0_71 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_6556) begin
      ic_tag_valid_out_0_72 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_6572) begin
      ic_tag_valid_out_0_73 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_6588) begin
      ic_tag_valid_out_0_74 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_6604) begin
      ic_tag_valid_out_0_75 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_6620) begin
      ic_tag_valid_out_0_76 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_6636) begin
      ic_tag_valid_out_0_77 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_6652) begin
      ic_tag_valid_out_0_78 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_6668) begin
      ic_tag_valid_out_0_79 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_6684) begin
      ic_tag_valid_out_0_80 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_6700) begin
      ic_tag_valid_out_0_81 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_6716) begin
      ic_tag_valid_out_0_82 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_6732) begin
      ic_tag_valid_out_0_83 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_6748) begin
      ic_tag_valid_out_0_84 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_6764) begin
      ic_tag_valid_out_0_85 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_6780) begin
      ic_tag_valid_out_0_86 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_6796) begin
      ic_tag_valid_out_0_87 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_6812) begin
      ic_tag_valid_out_0_88 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_6828) begin
      ic_tag_valid_out_0_89 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_6844) begin
      ic_tag_valid_out_0_90 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_6860) begin
      ic_tag_valid_out_0_91 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_6876) begin
      ic_tag_valid_out_0_92 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_6892) begin
      ic_tag_valid_out_0_93 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_6908) begin
      ic_tag_valid_out_0_94 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_6924) begin
      ic_tag_valid_out_0_95 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7452) begin
      ic_tag_valid_out_0_96 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_7468) begin
      ic_tag_valid_out_0_97 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_7484) begin
      ic_tag_valid_out_0_98 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_7500) begin
      ic_tag_valid_out_0_99 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_7516) begin
      ic_tag_valid_out_0_100 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_7532) begin
      ic_tag_valid_out_0_101 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_7548) begin
      ic_tag_valid_out_0_102 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_7564) begin
      ic_tag_valid_out_0_103 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_7580) begin
      ic_tag_valid_out_0_104 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_7596) begin
      ic_tag_valid_out_0_105 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_7612) begin
      ic_tag_valid_out_0_106 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_7628) begin
      ic_tag_valid_out_0_107 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_7644) begin
      ic_tag_valid_out_0_108 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_7660) begin
      ic_tag_valid_out_0_109 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_7676) begin
      ic_tag_valid_out_0_110 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_7692) begin
      ic_tag_valid_out_0_111 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_7708) begin
      ic_tag_valid_out_0_112 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_7724) begin
      ic_tag_valid_out_0_113 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_7740) begin
      ic_tag_valid_out_0_114 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_7756) begin
      ic_tag_valid_out_0_115 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_7772) begin
      ic_tag_valid_out_0_116 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_7788) begin
      ic_tag_valid_out_0_117 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_7804) begin
      ic_tag_valid_out_0_118 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_7820) begin
      ic_tag_valid_out_0_119 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_7836) begin
      ic_tag_valid_out_0_120 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_7852) begin
      ic_tag_valid_out_0_121 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_7868) begin
      ic_tag_valid_out_0_122 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_7884) begin
      ic_tag_valid_out_0_123 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_7900) begin
      ic_tag_valid_out_0_124 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_7916) begin
      ic_tag_valid_out_0_125 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_7932) begin
      ic_tag_valid_out_0_126 <= _T_4371;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_7948) begin
      ic_tag_valid_out_0_127 <= _T_4371;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_365 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_365 <= {{5'd0}, _T_364};
    end else begin
      _T_365 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_1682) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_1757) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_1801;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_1583) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_1585) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_1595) begin
        perr_state <= 3'h0;
      end else if (_T_1598) begin
        if (_T_1600) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_1604) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_1608) begin
        err_stop_state <= 2'h1;
      end else if (_T_1613) begin
        if (_T_1615) begin
          err_stop_state <= 2'h0;
        end else if (_T_1636) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_1640) begin
        if (_T_1615) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_1657) begin
        if (_T_1661) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_526;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_4284 <= 7'h0;
    end else if (_T_3105) begin
      _T_4284 <= io_ic_debug_addr[9:3];
    end else begin
      _T_4284 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_566;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3040;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_2215;
    end else begin
      iccm_dma_rdata <= _T_2216;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3036;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3105) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3108) begin
      way_status_new_ff <= _T_3112;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3108) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_9301 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9301 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_9271 <= 1'h0;
    end else begin
      _T_9271 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_9272 <= 1'h0;
    end else begin
      _T_9272 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_9273 <= 1'h0;
    end else begin
      _T_9273 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_9277 <= 1'h0;
    end else begin
      _T_9277 <= _T_9276;
    end
    if (reset) begin
      _T_9278 <= 1'h0;
    end else begin
      _T_9278 <= bus_cmd_sent;
    end
  end
endmodule
