module el2_ifu_compress_ctl(
  input         clock,
  input         reset,
  input  [15:0] io_din,
  output [31:0] io_dout,
  output [31:0] io_l1,
  output [31:0] io_l2,
  output [31:0] io_l3,
  output        io_legal,
  output [31:0] io_o
);
  wire  _T_2 = ~io_din[14]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_4 = ~io_din[13]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_7 = ~io_din[6]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_9 = ~io_din[5]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_11 = io_din[15] & _T_2; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_12 = _T_11 & _T_4; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_13 = _T_12 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_14 = _T_13 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_15 = _T_14 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_16 = _T_15 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_23 = ~io_din[11]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_28 = _T_12 & _T_23; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_29 = _T_28 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_30 = _T_29 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  out_30 = _T_16 | _T_30; // @[el2_ifu_compress_ctl.scala 23:53]
  wire  _T_38 = ~io_din[10]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_40 = ~io_din[9]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_42 = ~io_din[8]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_44 = ~io_din[7]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_50 = ~io_din[4]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_52 = ~io_din[3]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_54 = ~io_din[2]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_56 = _T_2 & io_din[12]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_57 = _T_56 & _T_23; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_58 = _T_57 & _T_38; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_59 = _T_58 & _T_40; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_60 = _T_59 & _T_42; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_61 = _T_60 & _T_44; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_62 = _T_61 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_63 = _T_62 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_64 = _T_63 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_65 = _T_64 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_66 = _T_65 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  out_20 = _T_66 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_79 = _T_28 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_90 = _T_12 & _T_38; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_91 = _T_90 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_92 = _T_79 | _T_91; // @[el2_ifu_compress_ctl.scala 25:46]
  wire  _T_102 = _T_12 & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_103 = _T_102 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_104 = _T_92 | _T_103; // @[el2_ifu_compress_ctl.scala 25:80]
  wire  _T_114 = _T_12 & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_115 = _T_114 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  out_14 = _T_104 | _T_115; // @[el2_ifu_compress_ctl.scala 25:113]
  wire  _T_128 = _T_12 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_129 = _T_128 & _T_38; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_130 = _T_129 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_142 = _T_128 & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_143 = _T_142 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_144 = _T_130 | _T_143; // @[el2_ifu_compress_ctl.scala 27:50]
  wire  _T_147 = ~io_din[0]; // @[el2_ifu_compress_ctl.scala 27:101]
  wire  _T_148 = io_din[14] & _T_147; // @[el2_ifu_compress_ctl.scala 27:99]
  wire  out_13 = _T_144 | _T_148; // @[el2_ifu_compress_ctl.scala 27:86]
  wire  _T_161 = _T_102 & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_162 = _T_161 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_175 = _T_162 | _T_79; // @[el2_ifu_compress_ctl.scala 28:47]
  wire  _T_188 = _T_175 | _T_91; // @[el2_ifu_compress_ctl.scala 28:81]
  wire  _T_190 = ~io_din[15]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_194 = _T_190 & _T_2; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_195 = _T_194 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_196 = _T_188 | _T_195; // @[el2_ifu_compress_ctl.scala 28:115]
  wire  _T_200 = io_din[15] & io_din[14]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_201 = _T_200 & io_din[13]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  out_12 = _T_196 | _T_201; // @[el2_ifu_compress_ctl.scala 29:26]
  wire  _T_217 = _T_11 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_218 = _T_217 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_219 = _T_218 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_220 = _T_219 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_221 = _T_220 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_224 = _T_221 & _T_147; // @[el2_ifu_compress_ctl.scala 30:53]
  wire  _T_228 = _T_2 & io_din[13]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_229 = _T_224 | _T_228; // @[el2_ifu_compress_ctl.scala 30:67]
  wire  _T_234 = _T_200 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  out_6 = _T_229 | _T_234; // @[el2_ifu_compress_ctl.scala 30:88]
  wire  _T_239 = io_din[15] & _T_147; // @[el2_ifu_compress_ctl.scala 32:24]
  wire  _T_243 = io_din[15] & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_244 = _T_243 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_245 = _T_239 | _T_244; // @[el2_ifu_compress_ctl.scala 32:39]
  wire  _T_249 = io_din[13] & _T_42; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_250 = _T_245 | _T_249; // @[el2_ifu_compress_ctl.scala 32:63]
  wire  _T_253 = io_din[13] & io_din[7]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_254 = _T_250 | _T_253; // @[el2_ifu_compress_ctl.scala 32:83]
  wire  _T_257 = io_din[13] & io_din[9]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_258 = _T_254 | _T_257; // @[el2_ifu_compress_ctl.scala 32:102]
  wire  _T_261 = io_din[13] & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_262 = _T_258 | _T_261; // @[el2_ifu_compress_ctl.scala 33:22]
  wire  _T_265 = io_din[13] & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_266 = _T_262 | _T_265; // @[el2_ifu_compress_ctl.scala 33:42]
  wire  _T_271 = _T_266 | _T_228; // @[el2_ifu_compress_ctl.scala 33:62]
  wire  out_5 = _T_271 | _T_200; // @[el2_ifu_compress_ctl.scala 33:83]
  wire  _T_288 = _T_2 & _T_23; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_289 = _T_288 & _T_38; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_290 = _T_289 & _T_40; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_291 = _T_290 & _T_42; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_292 = _T_291 & _T_44; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_295 = _T_292 & _T_147; // @[el2_ifu_compress_ctl.scala 36:50]
  wire  _T_303 = _T_194 & _T_147; // @[el2_ifu_compress_ctl.scala 36:87]
  wire  _T_304 = _T_295 | _T_303; // @[el2_ifu_compress_ctl.scala 36:65]
  wire  _T_308 = _T_2 & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_311 = _T_308 & _T_147; // @[el2_ifu_compress_ctl.scala 37:23]
  wire  _T_312 = _T_304 | _T_311; // @[el2_ifu_compress_ctl.scala 36:102]
  wire  _T_317 = _T_190 & io_din[14]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_318 = _T_317 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_319 = _T_312 | _T_318; // @[el2_ifu_compress_ctl.scala 37:38]
  wire  _T_323 = _T_2 & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_326 = _T_323 & _T_147; // @[el2_ifu_compress_ctl.scala 37:82]
  wire  _T_327 = _T_319 | _T_326; // @[el2_ifu_compress_ctl.scala 37:62]
  wire  _T_331 = _T_2 & io_din[4]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_334 = _T_331 & _T_147; // @[el2_ifu_compress_ctl.scala 38:23]
  wire  _T_335 = _T_327 | _T_334; // @[el2_ifu_compress_ctl.scala 37:97]
  wire  _T_339 = _T_2 & io_din[3]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_342 = _T_339 & _T_147; // @[el2_ifu_compress_ctl.scala 38:58]
  wire  _T_343 = _T_335 | _T_342; // @[el2_ifu_compress_ctl.scala 38:38]
  wire  _T_347 = _T_2 & io_din[2]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_350 = _T_347 & _T_147; // @[el2_ifu_compress_ctl.scala 38:93]
  wire  _T_351 = _T_343 | _T_350; // @[el2_ifu_compress_ctl.scala 38:73]
  wire  _T_357 = _T_2 & _T_4; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_358 = _T_357 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  out_4 = _T_351 | _T_358; // @[el2_ifu_compress_ctl.scala 38:108]
  wire  _T_380 = _T_56 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_381 = _T_380 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_382 = _T_381 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_383 = _T_382 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_384 = _T_383 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_385 = _T_384 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_386 = _T_385 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_403 = _T_56 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_404 = _T_403 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_405 = _T_404 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_406 = _T_405 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_407 = _T_406 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_408 = _T_407 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_409 = _T_408 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_410 = _T_386 | _T_409; // @[el2_ifu_compress_ctl.scala 45:59]
  wire  _T_427 = _T_56 & io_din[9]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_428 = _T_427 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_429 = _T_428 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_430 = _T_429 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_431 = _T_430 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_432 = _T_431 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_433 = _T_432 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_434 = _T_410 | _T_433; // @[el2_ifu_compress_ctl.scala 46:59]
  wire  _T_451 = _T_56 & io_din[8]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_452 = _T_451 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_453 = _T_452 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_454 = _T_453 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_455 = _T_454 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_456 = _T_455 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_457 = _T_456 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_458 = _T_434 | _T_457; // @[el2_ifu_compress_ctl.scala 47:58]
  wire  _T_475 = _T_56 & io_din[7]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_476 = _T_475 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_477 = _T_476 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_478 = _T_477 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_479 = _T_478 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_480 = _T_479 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_481 = _T_480 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_482 = _T_458 | _T_481; // @[el2_ifu_compress_ctl.scala 48:55]
  wire  _T_487 = ~io_din[12]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_499 = _T_11 & _T_487; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_500 = _T_499 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_501 = _T_500 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_502 = _T_501 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_503 = _T_502 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_504 = _T_503 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_507 = _T_504 & _T_147; // @[el2_ifu_compress_ctl.scala 50:56]
  wire  _T_508 = _T_482 | _T_507; // @[el2_ifu_compress_ctl.scala 49:57]
  wire  _T_514 = _T_190 & io_din[13]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_515 = _T_514 & _T_42; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_516 = _T_508 | _T_515; // @[el2_ifu_compress_ctl.scala 50:71]
  wire  _T_522 = _T_514 & io_din[7]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_523 = _T_516 | _T_522; // @[el2_ifu_compress_ctl.scala 51:34]
  wire  _T_529 = _T_514 & io_din[9]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_530 = _T_523 | _T_529; // @[el2_ifu_compress_ctl.scala 52:33]
  wire  _T_536 = _T_514 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_537 = _T_530 | _T_536; // @[el2_ifu_compress_ctl.scala 53:33]
  wire  _T_543 = _T_514 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_544 = _T_537 | _T_543; // @[el2_ifu_compress_ctl.scala 54:34]
  wire  out_2 = _T_544 | _T_228; // @[el2_ifu_compress_ctl.scala 55:34]
  wire [4:0] rs2d = io_din[6:2]; // @[el2_ifu_compress_ctl.scala 64:20]
  wire [4:0] rdd = io_din[11:7]; // @[el2_ifu_compress_ctl.scala 65:19]
  wire [4:0] rdpd = {2'h1,io_din[9:7]}; // @[Cat.scala 29:58]
  wire [4:0] rs2pd = {2'h1,io_din[4:2]}; // @[Cat.scala 29:58]
  wire  _T_557 = _T_308 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_564 = _T_317 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_565 = _T_564 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_566 = _T_557 | _T_565; // @[el2_ifu_compress_ctl.scala 69:33]
  wire  _T_572 = _T_323 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_573 = _T_566 | _T_572; // @[el2_ifu_compress_ctl.scala 69:58]
  wire  _T_580 = _T_317 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_581 = _T_580 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_582 = _T_573 | _T_581; // @[el2_ifu_compress_ctl.scala 69:79]
  wire  _T_588 = _T_331 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_589 = _T_582 | _T_588; // @[el2_ifu_compress_ctl.scala 69:104]
  wire  _T_596 = _T_317 & io_din[9]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_597 = _T_596 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_598 = _T_589 | _T_597; // @[el2_ifu_compress_ctl.scala 70:24]
  wire  _T_604 = _T_339 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_605 = _T_598 | _T_604; // @[el2_ifu_compress_ctl.scala 70:48]
  wire  _T_613 = _T_317 & _T_42; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_614 = _T_613 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_615 = _T_605 | _T_614; // @[el2_ifu_compress_ctl.scala 70:69]
  wire  _T_621 = _T_347 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_622 = _T_615 | _T_621; // @[el2_ifu_compress_ctl.scala 70:94]
  wire  _T_629 = _T_317 & io_din[7]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_630 = _T_629 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_631 = _T_622 | _T_630; // @[el2_ifu_compress_ctl.scala 71:22]
  wire  _T_635 = _T_190 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_636 = _T_631 | _T_635; // @[el2_ifu_compress_ctl.scala 71:46]
  wire  _T_642 = _T_190 & _T_4; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_643 = _T_642 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  rdrd = _T_636 | _T_643; // @[el2_ifu_compress_ctl.scala 71:65]
  wire  _T_651 = _T_380 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_659 = _T_403 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_660 = _T_651 | _T_659; // @[el2_ifu_compress_ctl.scala 73:38]
  wire  _T_668 = _T_427 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_669 = _T_660 | _T_668; // @[el2_ifu_compress_ctl.scala 73:63]
  wire  _T_677 = _T_451 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_678 = _T_669 | _T_677; // @[el2_ifu_compress_ctl.scala 73:87]
  wire  _T_686 = _T_475 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_687 = _T_678 | _T_686; // @[el2_ifu_compress_ctl.scala 73:111]
  wire  _T_703 = _T_2 & _T_487; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_704 = _T_703 & _T_7; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_705 = _T_704 & _T_9; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_706 = _T_705 & _T_50; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_707 = _T_706 & _T_52; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_708 = _T_707 & _T_54; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_709 = _T_708 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_710 = _T_687 | _T_709; // @[el2_ifu_compress_ctl.scala 74:27]
  wire  _T_717 = _T_56 & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_718 = _T_717 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_719 = _T_710 | _T_718; // @[el2_ifu_compress_ctl.scala 74:65]
  wire  _T_726 = _T_56 & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_727 = _T_726 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_728 = _T_719 | _T_727; // @[el2_ifu_compress_ctl.scala 74:89]
  wire  _T_735 = _T_56 & io_din[4]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_736 = _T_735 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_737 = _T_728 | _T_736; // @[el2_ifu_compress_ctl.scala 74:113]
  wire  _T_744 = _T_56 & io_din[3]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_745 = _T_744 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_746 = _T_737 | _T_745; // @[el2_ifu_compress_ctl.scala 75:27]
  wire  _T_753 = _T_56 & io_din[2]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_754 = _T_753 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_755 = _T_746 | _T_754; // @[el2_ifu_compress_ctl.scala 75:51]
  wire  _T_764 = _T_194 & _T_4; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_765 = _T_764 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  rdrs1 = _T_755 | _T_765; // @[el2_ifu_compress_ctl.scala 75:75]
  wire  _T_769 = io_din[15] & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_770 = _T_769 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_774 = io_din[15] & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_775 = _T_774 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_776 = _T_770 | _T_775; // @[el2_ifu_compress_ctl.scala 77:34]
  wire  _T_780 = io_din[15] & io_din[4]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_781 = _T_780 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_782 = _T_776 | _T_781; // @[el2_ifu_compress_ctl.scala 77:54]
  wire  _T_786 = io_din[15] & io_din[3]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_787 = _T_786 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_788 = _T_782 | _T_787; // @[el2_ifu_compress_ctl.scala 77:74]
  wire  _T_792 = io_din[15] & io_din[2]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_793 = _T_792 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_794 = _T_788 | _T_793; // @[el2_ifu_compress_ctl.scala 77:94]
  wire  _T_799 = _T_200 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  rs2rs2 = _T_794 | _T_799; // @[el2_ifu_compress_ctl.scala 77:114]
  wire  rdprd = _T_12 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_812 = io_din[15] & _T_4; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_813 = _T_812 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_819 = _T_813 | _T_234; // @[el2_ifu_compress_ctl.scala 81:36]
  wire  _T_822 = ~io_din[1]; // @[el2_ifu_compress_ctl.scala 20:83]
  wire  _T_823 = io_din[14] & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_826 = _T_823 & _T_147; // @[el2_ifu_compress_ctl.scala 81:76]
  wire  rdprs1 = _T_819 | _T_826; // @[el2_ifu_compress_ctl.scala 81:57]
  wire  _T_838 = _T_128 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_839 = _T_838 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_843 = io_din[15] & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_846 = _T_843 & _T_147; // @[el2_ifu_compress_ctl.scala 83:66]
  wire  rs2prs2 = _T_839 | _T_846; // @[el2_ifu_compress_ctl.scala 83:47]
  wire  _T_851 = _T_190 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  rs2prd = _T_851 & _T_147; // @[el2_ifu_compress_ctl.scala 84:33]
  wire  _T_858 = _T_2 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  uimm9_2 = _T_858 & _T_147; // @[el2_ifu_compress_ctl.scala 85:34]
  wire  _T_867 = _T_317 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  ulwimm6_2 = _T_867 & _T_147; // @[el2_ifu_compress_ctl.scala 86:39]
  wire  ulwspimm7_2 = _T_317 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_889 = _T_317 & io_din[13]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_890 = _T_889 & _T_23; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_891 = _T_890 & _T_38; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_892 = _T_891 & _T_40; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_893 = _T_892 & io_din[8]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  rdeq2 = _T_893 & _T_44; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1019 = _T_194 & io_din[13]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  rdeq1 = _T_482 | _T_1019; // @[el2_ifu_compress_ctl.scala 91:42]
  wire  _T_1042 = io_din[14] & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1043 = rdeq2 | _T_1042; // @[el2_ifu_compress_ctl.scala 92:53]
  wire  rs1eq2 = _T_1043 | uimm9_2; // @[el2_ifu_compress_ctl.scala 92:71]
  wire  _T_1084 = _T_357 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1085 = _T_1084 & _T_38; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1086 = _T_1085 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  simm5_0 = _T_1086 | _T_643; // @[el2_ifu_compress_ctl.scala 95:45]
  wire  _T_1104 = _T_889 & io_din[7]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1113 = _T_889 & _T_42; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1114 = _T_1104 | _T_1113; // @[el2_ifu_compress_ctl.scala 97:44]
  wire  _T_1122 = _T_889 & io_din[9]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1123 = _T_1114 | _T_1122; // @[el2_ifu_compress_ctl.scala 97:70]
  wire  _T_1131 = _T_889 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1132 = _T_1123 | _T_1131; // @[el2_ifu_compress_ctl.scala 97:95]
  wire  _T_1140 = _T_889 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  sluimm17_12 = _T_1132 | _T_1140; // @[el2_ifu_compress_ctl.scala 98:29]
  wire  uimm5_0 = _T_79 | _T_195; // @[el2_ifu_compress_ctl.scala 99:45]
  wire [6:0] l1_6 = {out_6,out_5,out_4,_T_228,out_2,1'h1,1'h1}; // @[Cat.scala 29:58]
  wire [4:0] _T_1184 = rdrd ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1185 = rdprd ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1186 = rs2prd ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1187 = rdeq1 ? 5'h1 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1188 = rdeq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1189 = _T_1184 | _T_1185; // @[Mux.scala 27:72]
  wire [4:0] _T_1190 = _T_1189 | _T_1186; // @[Mux.scala 27:72]
  wire [4:0] _T_1191 = _T_1190 | _T_1187; // @[Mux.scala 27:72]
  wire [4:0] l1_11 = _T_1191 | _T_1188; // @[Mux.scala 27:72]
  wire [4:0] _T_1202 = rdrs1 ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1203 = rdprs1 ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1204 = rs1eq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1205 = _T_1202 | _T_1203; // @[Mux.scala 27:72]
  wire [4:0] l1_19 = _T_1205 | _T_1204; // @[Mux.scala 27:72]
  wire [4:0] _T_1211 = {3'h0,1'h0,out_20}; // @[Cat.scala 29:58]
  wire [4:0] _T_1214 = rs2rs2 ? rs2d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1215 = rs2prs2 ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1216 = _T_1214 | _T_1215; // @[Mux.scala 27:72]
  wire [4:0] l1_24 = _T_1211 | _T_1216; // @[el2_ifu_compress_ctl.scala 110:67]
  wire [14:0] _T_1224 = {out_14,out_13,out_12,l1_11,l1_6}; // @[Cat.scala 29:58]
  wire [16:0] _T_1226 = {1'h0,out_30,2'h0,3'h0,l1_24,l1_19}; // @[Cat.scala 29:58]
  wire [31:0] l1 = {1'h0,out_30,2'h0,3'h0,l1_24,l1_19,_T_1224}; // @[Cat.scala 29:58]
  wire [5:0] simm5d = {io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [5:0] simm9d = {io_din[12],io_din[4:3],io_din[5],io_din[2],io_din[6]}; // @[Cat.scala 29:58]
  wire [8:0] sjald_12 = io_din[12] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [19:0] sjald = {sjald_12,io_din[12],io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:4],io_din[3]}; // @[Cat.scala 29:58]
  wire [14:0] _T_1273 = io_din[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [19:0] sluimmd = {_T_1273,rs2d}; // @[Cat.scala 29:58]
  wire [6:0] _T_1279 = simm5d[5] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_1281 = {_T_1279,simm5d[4:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1284 = {2'h0,io_din[10:7],io_din[12:11],io_din[5],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [2:0] _T_1288 = simm9d[5] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_1291 = {_T_1288,simm9d[4:0],4'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1294 = {5'h0,io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1297 = {4'h0,io_din[3:2],io_din[12],io_din[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1299 = {6'h0,io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1304 = {sjald[19],sjald[9:0],sjald[10]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1306 = simm5_0 ? _T_1281 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1307 = uimm9_2 ? _T_1284 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1308 = rdeq2 ? _T_1291 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1309 = ulwimm6_2 ? _T_1294 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1310 = ulwspimm7_2 ? _T_1297 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1311 = uimm5_0 ? _T_1299 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1312 = _T_228 ? _T_1304 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1313 = sluimm17_12 ? sluimmd[19:8] : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1314 = _T_1306 | _T_1307; // @[Mux.scala 27:72]
  wire [11:0] _T_1315 = _T_1314 | _T_1308; // @[Mux.scala 27:72]
  wire [11:0] _T_1316 = _T_1315 | _T_1309; // @[Mux.scala 27:72]
  wire [11:0] _T_1317 = _T_1316 | _T_1310; // @[Mux.scala 27:72]
  wire [11:0] _T_1318 = _T_1317 | _T_1311; // @[Mux.scala 27:72]
  wire [11:0] _T_1319 = _T_1318 | _T_1312; // @[Mux.scala 27:72]
  wire [11:0] _T_1320 = _T_1319 | _T_1313; // @[Mux.scala 27:72]
  wire [11:0] l2_31 = l1[31:20] | _T_1320; // @[el2_ifu_compress_ctl.scala 126:25]
  wire [8:0] _T_1327 = _T_228 ? sjald[19:11] : 9'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1328 = sluimm17_12 ? sluimmd[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [8:0] _GEN_0 = {{1'd0}, _T_1328}; // @[Mux.scala 27:72]
  wire [8:0] _T_1329 = _T_1327 | _GEN_0; // @[Mux.scala 27:72]
  wire [8:0] _GEN_1 = {{1'd0}, l1[19:12]}; // @[el2_ifu_compress_ctl.scala 136:25]
  wire [8:0] l2_19 = _GEN_1 | _T_1329; // @[el2_ifu_compress_ctl.scala 136:25]
  wire [32:0] l2 = {l2_31,l2_19,l1[11:0]}; // @[Cat.scala 29:58]
  wire [8:0] sbr8d = {io_din[12],io_din[6],io_din[5],io_din[2],io_din[11],io_din[10],io_din[4],io_din[3],1'h0}; // @[Cat.scala 29:58]
  wire [6:0] uswimm6d = {io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [7:0] uswspimm7d = {io_din[8:7],io_din[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_1360 = sbr8d[8] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _T_1362 = {_T_1360,sbr8d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1365 = {5'h0,uswimm6d[6:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1368 = {4'h0,uswspimm7d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1369 = _T_234 ? _T_1362 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1370 = _T_846 ? _T_1365 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1371 = _T_799 ? _T_1368 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1372 = _T_1369 | _T_1370; // @[Mux.scala 27:72]
  wire [6:0] _T_1373 = _T_1372 | _T_1371; // @[Mux.scala 27:72]
  wire [6:0] l3_31 = l2[31:25] | _T_1373; // @[el2_ifu_compress_ctl.scala 142:25]
  wire [12:0] l3_24 = l2[24:12]; // @[el2_ifu_compress_ctl.scala 145:17]
  wire [4:0] _T_1379 = {sbr8d[4:1],sbr8d[8]}; // @[Cat.scala 29:58]
  wire [4:0] _T_1384 = _T_234 ? _T_1379 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1385 = _T_846 ? uswimm6d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1386 = _T_799 ? uswspimm7d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1387 = _T_1384 | _T_1385; // @[Mux.scala 27:72]
  wire [4:0] _T_1388 = _T_1387 | _T_1386; // @[Mux.scala 27:72]
  wire [4:0] l3_11 = l2[11:7] | _T_1388; // @[el2_ifu_compress_ctl.scala 146:24]
  wire [11:0] _T_1391 = {l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire [19:0] _T_1392 = {l3_31,l3_24}; // @[Cat.scala 29:58]
  wire [31:0] l3 = {l3_31,l3_24,l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire  _T_1399 = _T_4 & _T_487; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1400 = _T_1399 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1401 = _T_1400 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1404 = _T_1401 & _T_147; // @[el2_ifu_compress_ctl.scala 151:39]
  wire  _T_1412 = _T_1399 & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1413 = _T_1412 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1416 = _T_1413 & _T_147; // @[el2_ifu_compress_ctl.scala 151:79]
  wire  _T_1417 = _T_1404 | _T_1416; // @[el2_ifu_compress_ctl.scala 151:54]
  wire  _T_1426 = _T_642 & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1427 = _T_1426 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1428 = _T_1417 | _T_1427; // @[el2_ifu_compress_ctl.scala 151:94]
  wire  _T_1436 = _T_1399 & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1437 = _T_1436 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1440 = _T_1437 & _T_147; // @[el2_ifu_compress_ctl.scala 152:55]
  wire  _T_1441 = _T_1428 | _T_1440; // @[el2_ifu_compress_ctl.scala 152:30]
  wire  _T_1449 = _T_1399 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1450 = _T_1449 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1453 = _T_1450 & _T_147; // @[el2_ifu_compress_ctl.scala 152:96]
  wire  _T_1454 = _T_1441 | _T_1453; // @[el2_ifu_compress_ctl.scala 152:70]
  wire  _T_1463 = _T_642 & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1464 = _T_1463 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1465 = _T_1454 | _T_1464; // @[el2_ifu_compress_ctl.scala 152:111]
  wire  _T_1472 = io_din[15] & _T_487; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1473 = _T_1472 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1474 = _T_1473 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1475 = _T_1465 | _T_1474; // @[el2_ifu_compress_ctl.scala 153:29]
  wire  _T_1483 = _T_1399 & io_din[9]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1484 = _T_1483 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1487 = _T_1484 & _T_147; // @[el2_ifu_compress_ctl.scala 153:79]
  wire  _T_1488 = _T_1475 | _T_1487; // @[el2_ifu_compress_ctl.scala 153:54]
  wire  _T_1495 = _T_487 & io_din[6]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1496 = _T_1495 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1497 = _T_1496 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1498 = _T_1488 | _T_1497; // @[el2_ifu_compress_ctl.scala 153:94]
  wire  _T_1507 = _T_642 & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1508 = _T_1507 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1509 = _T_1498 | _T_1508; // @[el2_ifu_compress_ctl.scala 153:118]
  wire  _T_1517 = _T_1399 & io_din[8]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1518 = _T_1517 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1521 = _T_1518 & _T_147; // @[el2_ifu_compress_ctl.scala 154:28]
  wire  _T_1522 = _T_1509 | _T_1521; // @[el2_ifu_compress_ctl.scala 153:144]
  wire  _T_1529 = _T_487 & io_din[5]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1530 = _T_1529 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1531 = _T_1530 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1532 = _T_1522 | _T_1531; // @[el2_ifu_compress_ctl.scala 154:43]
  wire  _T_1541 = _T_642 & io_din[10]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1542 = _T_1541 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1543 = _T_1532 | _T_1542; // @[el2_ifu_compress_ctl.scala 154:67]
  wire  _T_1551 = _T_1399 & io_din[7]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1552 = _T_1551 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1555 = _T_1552 & _T_147; // @[el2_ifu_compress_ctl.scala 155:28]
  wire  _T_1556 = _T_1543 | _T_1555; // @[el2_ifu_compress_ctl.scala 154:94]
  wire  _T_1564 = io_din[12] & io_din[11]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1565 = _T_1564 & _T_38; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1566 = _T_1565 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1567 = _T_1566 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1568 = _T_1556 | _T_1567; // @[el2_ifu_compress_ctl.scala 155:43]
  wire  _T_1577 = _T_642 & io_din[9]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1578 = _T_1577 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1579 = _T_1568 | _T_1578; // @[el2_ifu_compress_ctl.scala 155:71]
  wire  _T_1587 = _T_1399 & io_din[4]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1588 = _T_1587 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1591 = _T_1588 & _T_147; // @[el2_ifu_compress_ctl.scala 156:28]
  wire  _T_1592 = _T_1579 | _T_1591; // @[el2_ifu_compress_ctl.scala 155:97]
  wire  _T_1598 = io_din[13] & io_din[12]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1599 = _T_1598 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1600 = _T_1599 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1601 = _T_1592 | _T_1600; // @[el2_ifu_compress_ctl.scala 156:43]
  wire  _T_1610 = _T_642 & io_din[8]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1611 = _T_1610 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1612 = _T_1601 | _T_1611; // @[el2_ifu_compress_ctl.scala 156:67]
  wire  _T_1620 = _T_1399 & io_din[3]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1621 = _T_1620 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1624 = _T_1621 & _T_147; // @[el2_ifu_compress_ctl.scala 157:28]
  wire  _T_1625 = _T_1612 | _T_1624; // @[el2_ifu_compress_ctl.scala 156:93]
  wire  _T_1631 = io_din[13] & io_din[4]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1632 = _T_1631 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1633 = _T_1632 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1634 = _T_1625 | _T_1633; // @[el2_ifu_compress_ctl.scala 157:43]
  wire  _T_1642 = _T_1399 & io_din[2]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1643 = _T_1642 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1646 = _T_1643 & _T_147; // @[el2_ifu_compress_ctl.scala 157:91]
  wire  _T_1647 = _T_1634 | _T_1646; // @[el2_ifu_compress_ctl.scala 157:66]
  wire  _T_1656 = _T_642 & io_din[7]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1657 = _T_1656 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1658 = _T_1647 | _T_1657; // @[el2_ifu_compress_ctl.scala 157:106]
  wire  _T_1664 = io_din[13] & io_din[3]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1665 = _T_1664 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1666 = _T_1665 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1667 = _T_1658 | _T_1666; // @[el2_ifu_compress_ctl.scala 158:29]
  wire  _T_1673 = io_din[13] & io_din[2]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1674 = _T_1673 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1675 = _T_1674 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1676 = _T_1667 | _T_1675; // @[el2_ifu_compress_ctl.scala 158:52]
  wire  _T_1682 = io_din[14] & _T_4; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1683 = _T_1682 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1684 = _T_1676 | _T_1683; // @[el2_ifu_compress_ctl.scala 158:75]
  wire  _T_1693 = _T_703 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1694 = _T_1693 & io_din[0]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1695 = _T_1684 | _T_1694; // @[el2_ifu_compress_ctl.scala 158:98]
  wire  _T_1702 = _T_812 & io_din[12]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1703 = _T_1702 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1706 = _T_1703 & _T_147; // @[el2_ifu_compress_ctl.scala 159:54]
  wire  _T_1707 = _T_1695 | _T_1706; // @[el2_ifu_compress_ctl.scala 159:29]
  wire  _T_1716 = _T_642 & _T_487; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1717 = _T_1716 & io_din[1]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1720 = _T_1717 & _T_147; // @[el2_ifu_compress_ctl.scala 159:96]
  wire  _T_1721 = _T_1707 | _T_1720; // @[el2_ifu_compress_ctl.scala 159:69]
  wire  _T_1730 = _T_642 & io_din[12]; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1731 = _T_1730 & _T_822; // @[el2_ifu_compress_ctl.scala 20:110]
  wire  _T_1732 = _T_1721 | _T_1731; // @[el2_ifu_compress_ctl.scala 159:111]
  wire  _T_1739 = _T_1682 & _T_147; // @[el2_ifu_compress_ctl.scala 160:50]
  wire  legal = _T_1732 | _T_1739; // @[el2_ifu_compress_ctl.scala 160:30]
  wire [31:0] _T_1741 = legal ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [9:0] _T_1751 = {1'h0,out_30,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0}; // @[Cat.scala 29:58]
  wire [18:0] _T_1760 = {_T_1751,1'h0,out_20,1'h0,1'h0,1'h0,1'h0,1'h0,out_14,out_13}; // @[Cat.scala 29:58]
  wire [27:0] _T_1769 = {_T_1760,out_12,1'h0,1'h0,1'h0,1'h0,1'h0,out_6,out_5,out_4}; // @[Cat.scala 29:58]
  wire [30:0] _T_1772 = {_T_1769,_T_228,out_2,1'h1}; // @[Cat.scala 29:58]
  assign io_dout = l3 & _T_1741; // @[el2_ifu_compress_ctl.scala 162:10]
  assign io_l1 = {_T_1226,_T_1224}; // @[el2_ifu_compress_ctl.scala 163:9]
  assign io_l2 = l2[31:0]; // @[el2_ifu_compress_ctl.scala 164:9]
  assign io_l3 = {_T_1392,_T_1391}; // @[el2_ifu_compress_ctl.scala 165:9]
  assign io_legal = _T_1732 | _T_1739; // @[el2_ifu_compress_ctl.scala 166:12]
  assign io_o = {_T_1772,1'h1}; // @[el2_ifu_compress_ctl.scala 167:8]
endmodule
