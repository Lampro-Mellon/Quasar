module rvclkhdr(
  input   io_clk,
  input   io_en
);
  wire  clkhdr_Q; // @[lib.scala 334:26]
  wire  clkhdr_CK; // @[lib.scala 334:26]
  wire  clkhdr_EN; // @[lib.scala 334:26]
  wire  clkhdr_SE; // @[lib.scala 334:26]
  gated_latch clkhdr ( // @[lib.scala 334:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign clkhdr_CK = io_clk; // @[lib.scala 336:18]
  assign clkhdr_EN = io_en; // @[lib.scala 337:18]
  assign clkhdr_SE = 1'h0; // @[lib.scala 338:18]
endmodule
module ifu_bp_ctl(
  input         clock,
  input         reset,
  input         io_active_clk,
  input         io_ic_hit_f,
  input         io_exu_flush_final,
  input  [30:0] io_ifc_fetch_addr_f,
  input         io_ifc_fetch_req_f,
  input         io_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_dec_bp_dec_tlu_bpred_disable,
  input         io_dec_tlu_flush_lower_wb,
  input  [7:0]  io_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_bp_exu_i0_br_way_r,
  input         io_exu_bp_exu_mp_pkt_valid,
  input         io_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_bp_exu_mp_pkt_bits_br_error,
  input         io_exu_bp_exu_mp_pkt_bits_br_start_error,
  input         io_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_bp_exu_mp_pkt_bits_way,
  input         io_exu_bp_exu_mp_pkt_bits_pret,
  input  [30:0] io_exu_bp_exu_mp_pkt_bits_prett,
  input  [7:0]  io_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_bp_exu_mp_btag,
  input  [8:0]  io_dec_fa_error_index,
  output        io_ifu_bp_hit_taken_f,
  output [30:0] io_ifu_bp_btb_target_f,
  output        io_ifu_bp_inst_mask_f,
  output [7:0]  io_ifu_bp_fghr_f,
  output [1:0]  io_ifu_bp_way_f,
  output [1:0]  io_ifu_bp_ret_f,
  output [1:0]  io_ifu_bp_hist1_f,
  output [1:0]  io_ifu_bp_hist0_f,
  output [1:0]  io_ifu_bp_pc4_f,
  output [1:0]  io_ifu_bp_valid_f,
  output [11:0] io_ifu_bp_poffset_f,
  output [8:0]  io_ifu_bp_fa_index_f_0,
  output [8:0]  io_ifu_bp_fa_index_f_1,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [255:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_23_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_24_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_25_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_26_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_27_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_28_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_29_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_30_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_31_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_32_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_33_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_34_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_35_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_36_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_37_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_38_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_39_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_40_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_41_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_42_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_43_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_44_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_45_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_46_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_47_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_47_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_48_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_48_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_49_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_49_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_50_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_50_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_51_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_51_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_52_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_52_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_53_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_53_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_54_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_54_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_55_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_55_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_56_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_56_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_57_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_57_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_58_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_58_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_59_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_59_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_60_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_60_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_61_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_61_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_62_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_62_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_63_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_63_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_64_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_64_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_65_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_65_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_66_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_66_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_67_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_67_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_68_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_68_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_69_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_69_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_70_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_70_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_71_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_71_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_72_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_72_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_73_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_73_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_74_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_74_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_75_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_75_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_76_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_76_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_77_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_77_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_78_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_78_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_79_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_79_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_80_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_80_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_81_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_81_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_82_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_82_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_83_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_83_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_84_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_84_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_85_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_85_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_86_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_86_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_87_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_87_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_88_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_88_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_89_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_89_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_90_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_90_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_91_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_91_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_92_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_92_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_93_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_93_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_94_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_94_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_95_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_95_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_96_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_96_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_97_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_97_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_98_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_98_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_99_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_99_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_100_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_100_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_101_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_101_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_102_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_102_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_103_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_103_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_104_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_104_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_105_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_105_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_106_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_106_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_107_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_107_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_108_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_108_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_109_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_109_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_110_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_110_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_111_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_111_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_112_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_112_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_113_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_113_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_114_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_114_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_115_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_115_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_116_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_116_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_117_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_117_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_118_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_118_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_119_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_119_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_120_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_120_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_121_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_121_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_122_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_122_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_123_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_123_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_124_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_124_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_125_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_125_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_126_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_126_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_127_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_127_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_128_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_128_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_129_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_129_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_130_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_130_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_131_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_131_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_132_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_132_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_133_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_133_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_134_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_134_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_135_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_135_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_136_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_136_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_137_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_137_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_138_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_138_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_139_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_139_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_140_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_140_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_141_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_141_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_142_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_142_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_143_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_143_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_144_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_144_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_145_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_145_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_146_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_146_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_147_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_147_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_148_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_148_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_149_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_149_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_150_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_150_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_151_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_151_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_152_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_152_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_153_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_153_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_154_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_154_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_155_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_155_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_156_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_156_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_157_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_157_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_158_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_158_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_159_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_159_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_160_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_160_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_161_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_161_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_162_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_162_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_163_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_163_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_164_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_164_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_165_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_165_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_166_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_166_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_167_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_167_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_168_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_168_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_169_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_169_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_170_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_170_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_171_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_171_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_172_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_172_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_173_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_173_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_174_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_174_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_175_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_175_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_176_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_176_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_177_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_177_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_178_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_178_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_179_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_179_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_180_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_180_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_181_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_181_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_182_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_182_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_183_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_183_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_184_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_184_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_185_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_185_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_186_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_186_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_187_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_187_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_188_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_188_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_189_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_189_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_190_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_190_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_191_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_191_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_192_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_192_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_193_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_193_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_194_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_194_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_195_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_195_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_196_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_196_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_197_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_197_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_198_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_198_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_199_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_199_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_200_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_200_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_201_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_201_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_202_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_202_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_203_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_203_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_204_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_204_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_205_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_205_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_206_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_206_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_207_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_207_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_208_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_208_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_209_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_209_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_210_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_210_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_211_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_211_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_212_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_212_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_213_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_213_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_214_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_214_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_215_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_215_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_216_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_216_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_217_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_217_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_218_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_218_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_219_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_219_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_220_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_220_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_221_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_221_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_222_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_222_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_223_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_223_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_224_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_224_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_225_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_225_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_226_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_226_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_227_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_227_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_228_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_228_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_229_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_229_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_230_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_230_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_231_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_231_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_232_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_232_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_233_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_233_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_234_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_234_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_235_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_235_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_236_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_236_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_237_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_237_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_238_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_238_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_239_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_239_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_240_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_240_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_241_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_241_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_242_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_242_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_243_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_243_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_244_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_244_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_245_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_245_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_246_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_246_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_247_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_247_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_248_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_248_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_249_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_249_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_250_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_250_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_251_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_251_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_252_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_252_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_253_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_253_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_254_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_254_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_255_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_255_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_256_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_256_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_257_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_257_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_258_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_258_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_259_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_259_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_260_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_260_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_261_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_261_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_262_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_262_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_263_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_263_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_264_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_264_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_265_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_265_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_266_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_266_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_267_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_267_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_268_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_268_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_269_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_269_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_270_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_270_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_271_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_271_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_272_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_272_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_273_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_273_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_274_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_274_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_275_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_275_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_276_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_276_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_277_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_277_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_278_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_278_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_279_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_279_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_280_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_280_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_281_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_281_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_282_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_282_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_283_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_283_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_284_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_284_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_285_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_285_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_286_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_286_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_287_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_287_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_288_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_288_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_289_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_289_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_290_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_290_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_291_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_291_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_292_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_292_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_293_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_293_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_294_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_294_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_295_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_295_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_296_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_296_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_297_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_297_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_298_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_298_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_299_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_299_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_300_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_300_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_301_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_301_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_302_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_302_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_303_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_303_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_304_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_304_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_305_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_305_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_306_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_306_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_307_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_307_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_308_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_308_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_309_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_309_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_310_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_310_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_311_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_311_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_312_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_312_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_313_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_313_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_314_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_314_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_315_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_315_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_316_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_316_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_317_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_317_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_318_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_318_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_319_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_319_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_320_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_320_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_321_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_321_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_322_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_322_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_323_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_323_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_324_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_324_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_325_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_325_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_326_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_326_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_327_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_327_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_328_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_328_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_329_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_329_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_330_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_330_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_331_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_331_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_332_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_332_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_333_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_333_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_334_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_334_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_335_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_335_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_336_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_336_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_337_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_337_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_338_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_338_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_339_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_339_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_340_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_340_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_341_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_341_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_342_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_342_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_343_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_343_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_344_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_344_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_345_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_345_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_346_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_346_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_347_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_347_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_348_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_348_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_349_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_349_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_350_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_350_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_351_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_351_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_352_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_352_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_353_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_353_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_354_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_354_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_355_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_355_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_356_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_356_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_357_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_357_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_358_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_358_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_359_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_359_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_360_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_360_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_361_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_361_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_362_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_362_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_363_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_363_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_364_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_364_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_365_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_365_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_366_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_366_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_367_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_367_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_368_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_368_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_369_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_369_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_370_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_370_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_371_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_371_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_372_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_372_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_373_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_373_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_374_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_374_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_375_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_375_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_376_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_376_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_377_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_377_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_378_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_378_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_379_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_379_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_380_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_380_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_381_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_381_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_382_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_382_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_383_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_383_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_384_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_384_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_385_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_385_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_386_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_386_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_387_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_387_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_388_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_388_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_389_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_389_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_390_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_390_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_391_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_391_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_392_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_392_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_393_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_393_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_394_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_394_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_395_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_395_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_396_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_396_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_397_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_397_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_398_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_398_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_399_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_399_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_400_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_400_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_401_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_401_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_402_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_402_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_403_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_403_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_404_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_404_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_405_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_405_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_406_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_406_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_407_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_407_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_408_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_408_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_409_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_409_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_410_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_410_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_411_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_411_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_412_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_412_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_413_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_413_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_414_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_414_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_415_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_415_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_416_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_416_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_417_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_417_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_418_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_418_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_419_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_419_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_420_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_420_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_421_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_421_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_422_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_422_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_423_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_423_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_424_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_424_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_425_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_425_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_426_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_426_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_427_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_427_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_428_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_428_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_429_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_429_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_430_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_430_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_431_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_431_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_432_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_432_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_433_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_433_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_434_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_434_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_435_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_435_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_436_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_436_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_437_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_437_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_438_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_438_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_439_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_439_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_440_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_440_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_441_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_441_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_442_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_442_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_443_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_443_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_444_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_444_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_445_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_445_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_446_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_446_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_447_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_447_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_448_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_448_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_449_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_449_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_450_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_450_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_451_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_451_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_452_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_452_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_453_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_453_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_454_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_454_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_455_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_455_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_456_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_456_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_457_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_457_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_458_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_458_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_459_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_459_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_460_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_460_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_461_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_461_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_462_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_462_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_463_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_463_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_464_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_464_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_465_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_465_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_466_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_466_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_467_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_467_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_468_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_468_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_469_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_469_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_470_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_470_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_471_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_471_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_472_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_472_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_473_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_473_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_474_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_474_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_475_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_475_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_476_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_476_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_477_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_477_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_478_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_478_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_479_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_479_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_480_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_480_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_481_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_481_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_482_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_482_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_483_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_483_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_484_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_484_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_485_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_485_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_486_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_486_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_487_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_487_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_488_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_488_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_489_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_489_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_490_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_490_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_491_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_491_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_492_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_492_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_493_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_493_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_494_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_494_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_495_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_495_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_496_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_496_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_497_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_497_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_498_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_498_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_499_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_499_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_500_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_500_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_501_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_501_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_502_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_502_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_503_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_503_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_504_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_504_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_505_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_505_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_506_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_506_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_507_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_507_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_508_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_508_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_509_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_509_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_510_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_510_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_511_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_511_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_512_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_512_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_513_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_513_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_514_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_514_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_515_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_515_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_516_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_516_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_517_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_517_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_518_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_518_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_519_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_519_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_520_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_520_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_521_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_521_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_en; // @[lib.scala 343:22]
  wire  _T_21 = io_dec_bp_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 135:54]
  reg  leak_one_f_d1; // @[Reg.scala 27:20]
  wire  _T_22 = ~io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 135:102]
  wire  _T_23 = leak_one_f_d1 & _T_22; // @[ifu_bp_ctl.scala 135:100]
  wire  leak_one_f = _T_21 | _T_23; // @[ifu_bp_ctl.scala 135:83]
  wire  _T = ~leak_one_f; // @[ifu_bp_ctl.scala 82:58]
  wire  exu_mp_valid = io_exu_bp_exu_mp_pkt_bits_misp & _T; // @[ifu_bp_ctl.scala 82:56]
  wire  dec_tlu_error_wb = io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error | io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu_bp_ctl.scala 105:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[lib.scala 51:85]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_bp_ctl.scala 113:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[lib.scala 51:85]
  wire  _T_147 = ~io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 191:37]
  wire  _T_2149 = btb_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_2661 = _T_2149 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2151 = btb_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_2662 = _T_2151 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2917 = _T_2661 | _T_2662; // @[Mux.scala 27:72]
  wire  _T_2153 = btb_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_2663 = _T_2153 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2918 = _T_2917 | _T_2663; // @[Mux.scala 27:72]
  wire  _T_2155 = btb_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_2664 = _T_2155 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2919 = _T_2918 | _T_2664; // @[Mux.scala 27:72]
  wire  _T_2157 = btb_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_2665 = _T_2157 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2920 = _T_2919 | _T_2665; // @[Mux.scala 27:72]
  wire  _T_2159 = btb_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_2666 = _T_2159 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2921 = _T_2920 | _T_2666; // @[Mux.scala 27:72]
  wire  _T_2161 = btb_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_2667 = _T_2161 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2922 = _T_2921 | _T_2667; // @[Mux.scala 27:72]
  wire  _T_2163 = btb_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_2668 = _T_2163 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2923 = _T_2922 | _T_2668; // @[Mux.scala 27:72]
  wire  _T_2165 = btb_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_2669 = _T_2165 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2924 = _T_2923 | _T_2669; // @[Mux.scala 27:72]
  wire  _T_2167 = btb_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_2670 = _T_2167 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2925 = _T_2924 | _T_2670; // @[Mux.scala 27:72]
  wire  _T_2169 = btb_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_2671 = _T_2169 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2926 = _T_2925 | _T_2671; // @[Mux.scala 27:72]
  wire  _T_2171 = btb_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_2672 = _T_2171 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2927 = _T_2926 | _T_2672; // @[Mux.scala 27:72]
  wire  _T_2173 = btb_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_2673 = _T_2173 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2928 = _T_2927 | _T_2673; // @[Mux.scala 27:72]
  wire  _T_2175 = btb_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_2674 = _T_2175 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2929 = _T_2928 | _T_2674; // @[Mux.scala 27:72]
  wire  _T_2177 = btb_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_2675 = _T_2177 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2930 = _T_2929 | _T_2675; // @[Mux.scala 27:72]
  wire  _T_2179 = btb_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_2676 = _T_2179 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2931 = _T_2930 | _T_2676; // @[Mux.scala 27:72]
  wire  _T_2181 = btb_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_2677 = _T_2181 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2932 = _T_2931 | _T_2677; // @[Mux.scala 27:72]
  wire  _T_2183 = btb_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_2678 = _T_2183 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2933 = _T_2932 | _T_2678; // @[Mux.scala 27:72]
  wire  _T_2185 = btb_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_2679 = _T_2185 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2934 = _T_2933 | _T_2679; // @[Mux.scala 27:72]
  wire  _T_2187 = btb_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_2680 = _T_2187 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2935 = _T_2934 | _T_2680; // @[Mux.scala 27:72]
  wire  _T_2189 = btb_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_2681 = _T_2189 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2936 = _T_2935 | _T_2681; // @[Mux.scala 27:72]
  wire  _T_2191 = btb_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_2682 = _T_2191 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2937 = _T_2936 | _T_2682; // @[Mux.scala 27:72]
  wire  _T_2193 = btb_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_2683 = _T_2193 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2938 = _T_2937 | _T_2683; // @[Mux.scala 27:72]
  wire  _T_2195 = btb_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_2684 = _T_2195 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2939 = _T_2938 | _T_2684; // @[Mux.scala 27:72]
  wire  _T_2197 = btb_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_2685 = _T_2197 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2940 = _T_2939 | _T_2685; // @[Mux.scala 27:72]
  wire  _T_2199 = btb_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_2686 = _T_2199 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2941 = _T_2940 | _T_2686; // @[Mux.scala 27:72]
  wire  _T_2201 = btb_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_2687 = _T_2201 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2942 = _T_2941 | _T_2687; // @[Mux.scala 27:72]
  wire  _T_2203 = btb_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_2688 = _T_2203 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2943 = _T_2942 | _T_2688; // @[Mux.scala 27:72]
  wire  _T_2205 = btb_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_2689 = _T_2205 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2944 = _T_2943 | _T_2689; // @[Mux.scala 27:72]
  wire  _T_2207 = btb_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_2690 = _T_2207 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2945 = _T_2944 | _T_2690; // @[Mux.scala 27:72]
  wire  _T_2209 = btb_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_2691 = _T_2209 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2946 = _T_2945 | _T_2691; // @[Mux.scala 27:72]
  wire  _T_2211 = btb_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_2692 = _T_2211 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2947 = _T_2946 | _T_2692; // @[Mux.scala 27:72]
  wire  _T_2213 = btb_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_2693 = _T_2213 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2948 = _T_2947 | _T_2693; // @[Mux.scala 27:72]
  wire  _T_2215 = btb_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_2694 = _T_2215 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2949 = _T_2948 | _T_2694; // @[Mux.scala 27:72]
  wire  _T_2217 = btb_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_2695 = _T_2217 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2950 = _T_2949 | _T_2695; // @[Mux.scala 27:72]
  wire  _T_2219 = btb_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_2696 = _T_2219 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2951 = _T_2950 | _T_2696; // @[Mux.scala 27:72]
  wire  _T_2221 = btb_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_2697 = _T_2221 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2952 = _T_2951 | _T_2697; // @[Mux.scala 27:72]
  wire  _T_2223 = btb_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_2698 = _T_2223 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2953 = _T_2952 | _T_2698; // @[Mux.scala 27:72]
  wire  _T_2225 = btb_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_2699 = _T_2225 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2954 = _T_2953 | _T_2699; // @[Mux.scala 27:72]
  wire  _T_2227 = btb_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_2700 = _T_2227 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2955 = _T_2954 | _T_2700; // @[Mux.scala 27:72]
  wire  _T_2229 = btb_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_2701 = _T_2229 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2956 = _T_2955 | _T_2701; // @[Mux.scala 27:72]
  wire  _T_2231 = btb_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_2702 = _T_2231 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2957 = _T_2956 | _T_2702; // @[Mux.scala 27:72]
  wire  _T_2233 = btb_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_2703 = _T_2233 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2958 = _T_2957 | _T_2703; // @[Mux.scala 27:72]
  wire  _T_2235 = btb_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_2704 = _T_2235 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2959 = _T_2958 | _T_2704; // @[Mux.scala 27:72]
  wire  _T_2237 = btb_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_2705 = _T_2237 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2960 = _T_2959 | _T_2705; // @[Mux.scala 27:72]
  wire  _T_2239 = btb_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_2706 = _T_2239 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2961 = _T_2960 | _T_2706; // @[Mux.scala 27:72]
  wire  _T_2241 = btb_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_2707 = _T_2241 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2962 = _T_2961 | _T_2707; // @[Mux.scala 27:72]
  wire  _T_2243 = btb_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_2708 = _T_2243 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2963 = _T_2962 | _T_2708; // @[Mux.scala 27:72]
  wire  _T_2245 = btb_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_2709 = _T_2245 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2964 = _T_2963 | _T_2709; // @[Mux.scala 27:72]
  wire  _T_2247 = btb_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_2710 = _T_2247 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2965 = _T_2964 | _T_2710; // @[Mux.scala 27:72]
  wire  _T_2249 = btb_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_2711 = _T_2249 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2966 = _T_2965 | _T_2711; // @[Mux.scala 27:72]
  wire  _T_2251 = btb_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_2712 = _T_2251 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2967 = _T_2966 | _T_2712; // @[Mux.scala 27:72]
  wire  _T_2253 = btb_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_2713 = _T_2253 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2968 = _T_2967 | _T_2713; // @[Mux.scala 27:72]
  wire  _T_2255 = btb_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_2714 = _T_2255 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2969 = _T_2968 | _T_2714; // @[Mux.scala 27:72]
  wire  _T_2257 = btb_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_2715 = _T_2257 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2970 = _T_2969 | _T_2715; // @[Mux.scala 27:72]
  wire  _T_2259 = btb_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_2716 = _T_2259 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2971 = _T_2970 | _T_2716; // @[Mux.scala 27:72]
  wire  _T_2261 = btb_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_2717 = _T_2261 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2972 = _T_2971 | _T_2717; // @[Mux.scala 27:72]
  wire  _T_2263 = btb_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_2718 = _T_2263 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2973 = _T_2972 | _T_2718; // @[Mux.scala 27:72]
  wire  _T_2265 = btb_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_2719 = _T_2265 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2974 = _T_2973 | _T_2719; // @[Mux.scala 27:72]
  wire  _T_2267 = btb_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_2720 = _T_2267 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2975 = _T_2974 | _T_2720; // @[Mux.scala 27:72]
  wire  _T_2269 = btb_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_2721 = _T_2269 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2976 = _T_2975 | _T_2721; // @[Mux.scala 27:72]
  wire  _T_2271 = btb_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_2722 = _T_2271 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2977 = _T_2976 | _T_2722; // @[Mux.scala 27:72]
  wire  _T_2273 = btb_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_2723 = _T_2273 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2978 = _T_2977 | _T_2723; // @[Mux.scala 27:72]
  wire  _T_2275 = btb_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_2724 = _T_2275 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2979 = _T_2978 | _T_2724; // @[Mux.scala 27:72]
  wire  _T_2277 = btb_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_2725 = _T_2277 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2980 = _T_2979 | _T_2725; // @[Mux.scala 27:72]
  wire  _T_2279 = btb_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_2726 = _T_2279 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2981 = _T_2980 | _T_2726; // @[Mux.scala 27:72]
  wire  _T_2281 = btb_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_2727 = _T_2281 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2982 = _T_2981 | _T_2727; // @[Mux.scala 27:72]
  wire  _T_2283 = btb_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_2728 = _T_2283 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2983 = _T_2982 | _T_2728; // @[Mux.scala 27:72]
  wire  _T_2285 = btb_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_2729 = _T_2285 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2984 = _T_2983 | _T_2729; // @[Mux.scala 27:72]
  wire  _T_2287 = btb_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_2730 = _T_2287 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2985 = _T_2984 | _T_2730; // @[Mux.scala 27:72]
  wire  _T_2289 = btb_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_2731 = _T_2289 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2986 = _T_2985 | _T_2731; // @[Mux.scala 27:72]
  wire  _T_2291 = btb_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_2732 = _T_2291 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2987 = _T_2986 | _T_2732; // @[Mux.scala 27:72]
  wire  _T_2293 = btb_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_2733 = _T_2293 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2988 = _T_2987 | _T_2733; // @[Mux.scala 27:72]
  wire  _T_2295 = btb_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_2734 = _T_2295 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2989 = _T_2988 | _T_2734; // @[Mux.scala 27:72]
  wire  _T_2297 = btb_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_2735 = _T_2297 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2990 = _T_2989 | _T_2735; // @[Mux.scala 27:72]
  wire  _T_2299 = btb_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_2736 = _T_2299 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2991 = _T_2990 | _T_2736; // @[Mux.scala 27:72]
  wire  _T_2301 = btb_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_2737 = _T_2301 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2992 = _T_2991 | _T_2737; // @[Mux.scala 27:72]
  wire  _T_2303 = btb_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_2738 = _T_2303 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2993 = _T_2992 | _T_2738; // @[Mux.scala 27:72]
  wire  _T_2305 = btb_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_2739 = _T_2305 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2994 = _T_2993 | _T_2739; // @[Mux.scala 27:72]
  wire  _T_2307 = btb_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_2740 = _T_2307 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2995 = _T_2994 | _T_2740; // @[Mux.scala 27:72]
  wire  _T_2309 = btb_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_2741 = _T_2309 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2996 = _T_2995 | _T_2741; // @[Mux.scala 27:72]
  wire  _T_2311 = btb_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_2742 = _T_2311 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2997 = _T_2996 | _T_2742; // @[Mux.scala 27:72]
  wire  _T_2313 = btb_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_2743 = _T_2313 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2998 = _T_2997 | _T_2743; // @[Mux.scala 27:72]
  wire  _T_2315 = btb_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_2744 = _T_2315 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_2999 = _T_2998 | _T_2744; // @[Mux.scala 27:72]
  wire  _T_2317 = btb_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_2745 = _T_2317 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3000 = _T_2999 | _T_2745; // @[Mux.scala 27:72]
  wire  _T_2319 = btb_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_2746 = _T_2319 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3001 = _T_3000 | _T_2746; // @[Mux.scala 27:72]
  wire  _T_2321 = btb_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_2747 = _T_2321 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3002 = _T_3001 | _T_2747; // @[Mux.scala 27:72]
  wire  _T_2323 = btb_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_2748 = _T_2323 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3003 = _T_3002 | _T_2748; // @[Mux.scala 27:72]
  wire  _T_2325 = btb_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_2749 = _T_2325 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3004 = _T_3003 | _T_2749; // @[Mux.scala 27:72]
  wire  _T_2327 = btb_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_2750 = _T_2327 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3005 = _T_3004 | _T_2750; // @[Mux.scala 27:72]
  wire  _T_2329 = btb_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_2751 = _T_2329 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3006 = _T_3005 | _T_2751; // @[Mux.scala 27:72]
  wire  _T_2331 = btb_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_2752 = _T_2331 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3007 = _T_3006 | _T_2752; // @[Mux.scala 27:72]
  wire  _T_2333 = btb_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_2753 = _T_2333 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3008 = _T_3007 | _T_2753; // @[Mux.scala 27:72]
  wire  _T_2335 = btb_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_2754 = _T_2335 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3009 = _T_3008 | _T_2754; // @[Mux.scala 27:72]
  wire  _T_2337 = btb_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_2755 = _T_2337 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3010 = _T_3009 | _T_2755; // @[Mux.scala 27:72]
  wire  _T_2339 = btb_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_2756 = _T_2339 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3011 = _T_3010 | _T_2756; // @[Mux.scala 27:72]
  wire  _T_2341 = btb_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_2757 = _T_2341 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3012 = _T_3011 | _T_2757; // @[Mux.scala 27:72]
  wire  _T_2343 = btb_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_2758 = _T_2343 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3013 = _T_3012 | _T_2758; // @[Mux.scala 27:72]
  wire  _T_2345 = btb_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_2759 = _T_2345 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3014 = _T_3013 | _T_2759; // @[Mux.scala 27:72]
  wire  _T_2347 = btb_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_2760 = _T_2347 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3015 = _T_3014 | _T_2760; // @[Mux.scala 27:72]
  wire  _T_2349 = btb_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_2761 = _T_2349 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3016 = _T_3015 | _T_2761; // @[Mux.scala 27:72]
  wire  _T_2351 = btb_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_2762 = _T_2351 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3017 = _T_3016 | _T_2762; // @[Mux.scala 27:72]
  wire  _T_2353 = btb_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_2763 = _T_2353 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3018 = _T_3017 | _T_2763; // @[Mux.scala 27:72]
  wire  _T_2355 = btb_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_2764 = _T_2355 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3019 = _T_3018 | _T_2764; // @[Mux.scala 27:72]
  wire  _T_2357 = btb_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_2765 = _T_2357 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3020 = _T_3019 | _T_2765; // @[Mux.scala 27:72]
  wire  _T_2359 = btb_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_2766 = _T_2359 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3021 = _T_3020 | _T_2766; // @[Mux.scala 27:72]
  wire  _T_2361 = btb_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_2767 = _T_2361 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3022 = _T_3021 | _T_2767; // @[Mux.scala 27:72]
  wire  _T_2363 = btb_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_2768 = _T_2363 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3023 = _T_3022 | _T_2768; // @[Mux.scala 27:72]
  wire  _T_2365 = btb_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_2769 = _T_2365 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3024 = _T_3023 | _T_2769; // @[Mux.scala 27:72]
  wire  _T_2367 = btb_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_2770 = _T_2367 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3025 = _T_3024 | _T_2770; // @[Mux.scala 27:72]
  wire  _T_2369 = btb_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_2771 = _T_2369 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3026 = _T_3025 | _T_2771; // @[Mux.scala 27:72]
  wire  _T_2371 = btb_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_2772 = _T_2371 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3027 = _T_3026 | _T_2772; // @[Mux.scala 27:72]
  wire  _T_2373 = btb_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_2773 = _T_2373 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3028 = _T_3027 | _T_2773; // @[Mux.scala 27:72]
  wire  _T_2375 = btb_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_2774 = _T_2375 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3029 = _T_3028 | _T_2774; // @[Mux.scala 27:72]
  wire  _T_2377 = btb_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_2775 = _T_2377 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3030 = _T_3029 | _T_2775; // @[Mux.scala 27:72]
  wire  _T_2379 = btb_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_2776 = _T_2379 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3031 = _T_3030 | _T_2776; // @[Mux.scala 27:72]
  wire  _T_2381 = btb_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_2777 = _T_2381 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3032 = _T_3031 | _T_2777; // @[Mux.scala 27:72]
  wire  _T_2383 = btb_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_2778 = _T_2383 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3033 = _T_3032 | _T_2778; // @[Mux.scala 27:72]
  wire  _T_2385 = btb_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_2779 = _T_2385 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3034 = _T_3033 | _T_2779; // @[Mux.scala 27:72]
  wire  _T_2387 = btb_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_2780 = _T_2387 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3035 = _T_3034 | _T_2780; // @[Mux.scala 27:72]
  wire  _T_2389 = btb_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_2781 = _T_2389 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3036 = _T_3035 | _T_2781; // @[Mux.scala 27:72]
  wire  _T_2391 = btb_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_2782 = _T_2391 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3037 = _T_3036 | _T_2782; // @[Mux.scala 27:72]
  wire  _T_2393 = btb_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_2783 = _T_2393 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3038 = _T_3037 | _T_2783; // @[Mux.scala 27:72]
  wire  _T_2395 = btb_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_2784 = _T_2395 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3039 = _T_3038 | _T_2784; // @[Mux.scala 27:72]
  wire  _T_2397 = btb_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_2785 = _T_2397 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3040 = _T_3039 | _T_2785; // @[Mux.scala 27:72]
  wire  _T_2399 = btb_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_2786 = _T_2399 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3041 = _T_3040 | _T_2786; // @[Mux.scala 27:72]
  wire  _T_2401 = btb_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_2787 = _T_2401 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3042 = _T_3041 | _T_2787; // @[Mux.scala 27:72]
  wire  _T_2403 = btb_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_2788 = _T_2403 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3043 = _T_3042 | _T_2788; // @[Mux.scala 27:72]
  wire  _T_2405 = btb_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_2789 = _T_2405 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3044 = _T_3043 | _T_2789; // @[Mux.scala 27:72]
  wire  _T_2407 = btb_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_2790 = _T_2407 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3045 = _T_3044 | _T_2790; // @[Mux.scala 27:72]
  wire  _T_2409 = btb_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_2791 = _T_2409 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3046 = _T_3045 | _T_2791; // @[Mux.scala 27:72]
  wire  _T_2411 = btb_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_2792 = _T_2411 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3047 = _T_3046 | _T_2792; // @[Mux.scala 27:72]
  wire  _T_2413 = btb_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_2793 = _T_2413 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3048 = _T_3047 | _T_2793; // @[Mux.scala 27:72]
  wire  _T_2415 = btb_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_2794 = _T_2415 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3049 = _T_3048 | _T_2794; // @[Mux.scala 27:72]
  wire  _T_2417 = btb_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_2795 = _T_2417 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3050 = _T_3049 | _T_2795; // @[Mux.scala 27:72]
  wire  _T_2419 = btb_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_2796 = _T_2419 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3051 = _T_3050 | _T_2796; // @[Mux.scala 27:72]
  wire  _T_2421 = btb_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_2797 = _T_2421 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3052 = _T_3051 | _T_2797; // @[Mux.scala 27:72]
  wire  _T_2423 = btb_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_2798 = _T_2423 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3053 = _T_3052 | _T_2798; // @[Mux.scala 27:72]
  wire  _T_2425 = btb_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_2799 = _T_2425 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3054 = _T_3053 | _T_2799; // @[Mux.scala 27:72]
  wire  _T_2427 = btb_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_2800 = _T_2427 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3055 = _T_3054 | _T_2800; // @[Mux.scala 27:72]
  wire  _T_2429 = btb_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_2801 = _T_2429 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3056 = _T_3055 | _T_2801; // @[Mux.scala 27:72]
  wire  _T_2431 = btb_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_2802 = _T_2431 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3057 = _T_3056 | _T_2802; // @[Mux.scala 27:72]
  wire  _T_2433 = btb_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_2803 = _T_2433 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3058 = _T_3057 | _T_2803; // @[Mux.scala 27:72]
  wire  _T_2435 = btb_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_2804 = _T_2435 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3059 = _T_3058 | _T_2804; // @[Mux.scala 27:72]
  wire  _T_2437 = btb_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_2805 = _T_2437 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3060 = _T_3059 | _T_2805; // @[Mux.scala 27:72]
  wire  _T_2439 = btb_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_2806 = _T_2439 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3061 = _T_3060 | _T_2806; // @[Mux.scala 27:72]
  wire  _T_2441 = btb_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_2807 = _T_2441 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3062 = _T_3061 | _T_2807; // @[Mux.scala 27:72]
  wire  _T_2443 = btb_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_2808 = _T_2443 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3063 = _T_3062 | _T_2808; // @[Mux.scala 27:72]
  wire  _T_2445 = btb_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_2809 = _T_2445 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3064 = _T_3063 | _T_2809; // @[Mux.scala 27:72]
  wire  _T_2447 = btb_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_2810 = _T_2447 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3065 = _T_3064 | _T_2810; // @[Mux.scala 27:72]
  wire  _T_2449 = btb_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_2811 = _T_2449 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3066 = _T_3065 | _T_2811; // @[Mux.scala 27:72]
  wire  _T_2451 = btb_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_2812 = _T_2451 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3067 = _T_3066 | _T_2812; // @[Mux.scala 27:72]
  wire  _T_2453 = btb_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_2813 = _T_2453 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3068 = _T_3067 | _T_2813; // @[Mux.scala 27:72]
  wire  _T_2455 = btb_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_2814 = _T_2455 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3069 = _T_3068 | _T_2814; // @[Mux.scala 27:72]
  wire  _T_2457 = btb_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_2815 = _T_2457 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3070 = _T_3069 | _T_2815; // @[Mux.scala 27:72]
  wire  _T_2459 = btb_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_2816 = _T_2459 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3071 = _T_3070 | _T_2816; // @[Mux.scala 27:72]
  wire  _T_2461 = btb_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_2817 = _T_2461 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3072 = _T_3071 | _T_2817; // @[Mux.scala 27:72]
  wire  _T_2463 = btb_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_2818 = _T_2463 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3073 = _T_3072 | _T_2818; // @[Mux.scala 27:72]
  wire  _T_2465 = btb_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_2819 = _T_2465 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3074 = _T_3073 | _T_2819; // @[Mux.scala 27:72]
  wire  _T_2467 = btb_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_2820 = _T_2467 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3075 = _T_3074 | _T_2820; // @[Mux.scala 27:72]
  wire  _T_2469 = btb_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_2821 = _T_2469 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3076 = _T_3075 | _T_2821; // @[Mux.scala 27:72]
  wire  _T_2471 = btb_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_2822 = _T_2471 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3077 = _T_3076 | _T_2822; // @[Mux.scala 27:72]
  wire  _T_2473 = btb_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_2823 = _T_2473 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3078 = _T_3077 | _T_2823; // @[Mux.scala 27:72]
  wire  _T_2475 = btb_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_2824 = _T_2475 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3079 = _T_3078 | _T_2824; // @[Mux.scala 27:72]
  wire  _T_2477 = btb_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_2825 = _T_2477 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3080 = _T_3079 | _T_2825; // @[Mux.scala 27:72]
  wire  _T_2479 = btb_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_2826 = _T_2479 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3081 = _T_3080 | _T_2826; // @[Mux.scala 27:72]
  wire  _T_2481 = btb_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_2827 = _T_2481 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3082 = _T_3081 | _T_2827; // @[Mux.scala 27:72]
  wire  _T_2483 = btb_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_2828 = _T_2483 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3083 = _T_3082 | _T_2828; // @[Mux.scala 27:72]
  wire  _T_2485 = btb_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_2829 = _T_2485 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3084 = _T_3083 | _T_2829; // @[Mux.scala 27:72]
  wire  _T_2487 = btb_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_2830 = _T_2487 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3085 = _T_3084 | _T_2830; // @[Mux.scala 27:72]
  wire  _T_2489 = btb_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_2831 = _T_2489 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3086 = _T_3085 | _T_2831; // @[Mux.scala 27:72]
  wire  _T_2491 = btb_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_2832 = _T_2491 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3087 = _T_3086 | _T_2832; // @[Mux.scala 27:72]
  wire  _T_2493 = btb_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_2833 = _T_2493 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3088 = _T_3087 | _T_2833; // @[Mux.scala 27:72]
  wire  _T_2495 = btb_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_2834 = _T_2495 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3089 = _T_3088 | _T_2834; // @[Mux.scala 27:72]
  wire  _T_2497 = btb_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_2835 = _T_2497 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3090 = _T_3089 | _T_2835; // @[Mux.scala 27:72]
  wire  _T_2499 = btb_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_2836 = _T_2499 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3091 = _T_3090 | _T_2836; // @[Mux.scala 27:72]
  wire  _T_2501 = btb_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_2837 = _T_2501 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3092 = _T_3091 | _T_2837; // @[Mux.scala 27:72]
  wire  _T_2503 = btb_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_2838 = _T_2503 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3093 = _T_3092 | _T_2838; // @[Mux.scala 27:72]
  wire  _T_2505 = btb_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_2839 = _T_2505 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3094 = _T_3093 | _T_2839; // @[Mux.scala 27:72]
  wire  _T_2507 = btb_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_2840 = _T_2507 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3095 = _T_3094 | _T_2840; // @[Mux.scala 27:72]
  wire  _T_2509 = btb_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_2841 = _T_2509 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3096 = _T_3095 | _T_2841; // @[Mux.scala 27:72]
  wire  _T_2511 = btb_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_2842 = _T_2511 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3097 = _T_3096 | _T_2842; // @[Mux.scala 27:72]
  wire  _T_2513 = btb_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_2843 = _T_2513 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3098 = _T_3097 | _T_2843; // @[Mux.scala 27:72]
  wire  _T_2515 = btb_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_2844 = _T_2515 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3099 = _T_3098 | _T_2844; // @[Mux.scala 27:72]
  wire  _T_2517 = btb_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_2845 = _T_2517 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3100 = _T_3099 | _T_2845; // @[Mux.scala 27:72]
  wire  _T_2519 = btb_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_2846 = _T_2519 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3101 = _T_3100 | _T_2846; // @[Mux.scala 27:72]
  wire  _T_2521 = btb_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_2847 = _T_2521 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3102 = _T_3101 | _T_2847; // @[Mux.scala 27:72]
  wire  _T_2523 = btb_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_2848 = _T_2523 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3103 = _T_3102 | _T_2848; // @[Mux.scala 27:72]
  wire  _T_2525 = btb_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_2849 = _T_2525 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3104 = _T_3103 | _T_2849; // @[Mux.scala 27:72]
  wire  _T_2527 = btb_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_2850 = _T_2527 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3105 = _T_3104 | _T_2850; // @[Mux.scala 27:72]
  wire  _T_2529 = btb_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_2851 = _T_2529 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3106 = _T_3105 | _T_2851; // @[Mux.scala 27:72]
  wire  _T_2531 = btb_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_2852 = _T_2531 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3107 = _T_3106 | _T_2852; // @[Mux.scala 27:72]
  wire  _T_2533 = btb_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_2853 = _T_2533 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3108 = _T_3107 | _T_2853; // @[Mux.scala 27:72]
  wire  _T_2535 = btb_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_2854 = _T_2535 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3109 = _T_3108 | _T_2854; // @[Mux.scala 27:72]
  wire  _T_2537 = btb_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_2855 = _T_2537 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3110 = _T_3109 | _T_2855; // @[Mux.scala 27:72]
  wire  _T_2539 = btb_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_2856 = _T_2539 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3111 = _T_3110 | _T_2856; // @[Mux.scala 27:72]
  wire  _T_2541 = btb_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_2857 = _T_2541 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3112 = _T_3111 | _T_2857; // @[Mux.scala 27:72]
  wire  _T_2543 = btb_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_2858 = _T_2543 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3113 = _T_3112 | _T_2858; // @[Mux.scala 27:72]
  wire  _T_2545 = btb_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_2859 = _T_2545 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3114 = _T_3113 | _T_2859; // @[Mux.scala 27:72]
  wire  _T_2547 = btb_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_2860 = _T_2547 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3115 = _T_3114 | _T_2860; // @[Mux.scala 27:72]
  wire  _T_2549 = btb_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_2861 = _T_2549 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3116 = _T_3115 | _T_2861; // @[Mux.scala 27:72]
  wire  _T_2551 = btb_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_2862 = _T_2551 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3117 = _T_3116 | _T_2862; // @[Mux.scala 27:72]
  wire  _T_2553 = btb_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_2863 = _T_2553 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3118 = _T_3117 | _T_2863; // @[Mux.scala 27:72]
  wire  _T_2555 = btb_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_2864 = _T_2555 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3119 = _T_3118 | _T_2864; // @[Mux.scala 27:72]
  wire  _T_2557 = btb_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_2865 = _T_2557 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3120 = _T_3119 | _T_2865; // @[Mux.scala 27:72]
  wire  _T_2559 = btb_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_2866 = _T_2559 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3121 = _T_3120 | _T_2866; // @[Mux.scala 27:72]
  wire  _T_2561 = btb_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_2867 = _T_2561 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3122 = _T_3121 | _T_2867; // @[Mux.scala 27:72]
  wire  _T_2563 = btb_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_2868 = _T_2563 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3123 = _T_3122 | _T_2868; // @[Mux.scala 27:72]
  wire  _T_2565 = btb_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_2869 = _T_2565 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3124 = _T_3123 | _T_2869; // @[Mux.scala 27:72]
  wire  _T_2567 = btb_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_2870 = _T_2567 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3125 = _T_3124 | _T_2870; // @[Mux.scala 27:72]
  wire  _T_2569 = btb_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_2871 = _T_2569 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3126 = _T_3125 | _T_2871; // @[Mux.scala 27:72]
  wire  _T_2571 = btb_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_2872 = _T_2571 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3127 = _T_3126 | _T_2872; // @[Mux.scala 27:72]
  wire  _T_2573 = btb_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_2873 = _T_2573 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3128 = _T_3127 | _T_2873; // @[Mux.scala 27:72]
  wire  _T_2575 = btb_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_2874 = _T_2575 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3129 = _T_3128 | _T_2874; // @[Mux.scala 27:72]
  wire  _T_2577 = btb_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_2875 = _T_2577 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3130 = _T_3129 | _T_2875; // @[Mux.scala 27:72]
  wire  _T_2579 = btb_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_2876 = _T_2579 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3131 = _T_3130 | _T_2876; // @[Mux.scala 27:72]
  wire  _T_2581 = btb_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_2877 = _T_2581 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3132 = _T_3131 | _T_2877; // @[Mux.scala 27:72]
  wire  _T_2583 = btb_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_2878 = _T_2583 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3133 = _T_3132 | _T_2878; // @[Mux.scala 27:72]
  wire  _T_2585 = btb_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_2879 = _T_2585 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3134 = _T_3133 | _T_2879; // @[Mux.scala 27:72]
  wire  _T_2587 = btb_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_2880 = _T_2587 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3135 = _T_3134 | _T_2880; // @[Mux.scala 27:72]
  wire  _T_2589 = btb_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_2881 = _T_2589 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3136 = _T_3135 | _T_2881; // @[Mux.scala 27:72]
  wire  _T_2591 = btb_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_2882 = _T_2591 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3137 = _T_3136 | _T_2882; // @[Mux.scala 27:72]
  wire  _T_2593 = btb_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_2883 = _T_2593 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3138 = _T_3137 | _T_2883; // @[Mux.scala 27:72]
  wire  _T_2595 = btb_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_2884 = _T_2595 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3139 = _T_3138 | _T_2884; // @[Mux.scala 27:72]
  wire  _T_2597 = btb_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_2885 = _T_2597 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3140 = _T_3139 | _T_2885; // @[Mux.scala 27:72]
  wire  _T_2599 = btb_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_2886 = _T_2599 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3141 = _T_3140 | _T_2886; // @[Mux.scala 27:72]
  wire  _T_2601 = btb_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_2887 = _T_2601 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3142 = _T_3141 | _T_2887; // @[Mux.scala 27:72]
  wire  _T_2603 = btb_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_2888 = _T_2603 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3143 = _T_3142 | _T_2888; // @[Mux.scala 27:72]
  wire  _T_2605 = btb_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_2889 = _T_2605 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3144 = _T_3143 | _T_2889; // @[Mux.scala 27:72]
  wire  _T_2607 = btb_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_2890 = _T_2607 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3145 = _T_3144 | _T_2890; // @[Mux.scala 27:72]
  wire  _T_2609 = btb_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_2891 = _T_2609 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3146 = _T_3145 | _T_2891; // @[Mux.scala 27:72]
  wire  _T_2611 = btb_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_2892 = _T_2611 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3147 = _T_3146 | _T_2892; // @[Mux.scala 27:72]
  wire  _T_2613 = btb_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_2893 = _T_2613 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3148 = _T_3147 | _T_2893; // @[Mux.scala 27:72]
  wire  _T_2615 = btb_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_2894 = _T_2615 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3149 = _T_3148 | _T_2894; // @[Mux.scala 27:72]
  wire  _T_2617 = btb_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_2895 = _T_2617 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3150 = _T_3149 | _T_2895; // @[Mux.scala 27:72]
  wire  _T_2619 = btb_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_2896 = _T_2619 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3151 = _T_3150 | _T_2896; // @[Mux.scala 27:72]
  wire  _T_2621 = btb_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_2897 = _T_2621 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3152 = _T_3151 | _T_2897; // @[Mux.scala 27:72]
  wire  _T_2623 = btb_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_2898 = _T_2623 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3153 = _T_3152 | _T_2898; // @[Mux.scala 27:72]
  wire  _T_2625 = btb_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_2899 = _T_2625 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3154 = _T_3153 | _T_2899; // @[Mux.scala 27:72]
  wire  _T_2627 = btb_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_2900 = _T_2627 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3155 = _T_3154 | _T_2900; // @[Mux.scala 27:72]
  wire  _T_2629 = btb_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_2901 = _T_2629 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3156 = _T_3155 | _T_2901; // @[Mux.scala 27:72]
  wire  _T_2631 = btb_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_2902 = _T_2631 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3157 = _T_3156 | _T_2902; // @[Mux.scala 27:72]
  wire  _T_2633 = btb_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_2903 = _T_2633 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3158 = _T_3157 | _T_2903; // @[Mux.scala 27:72]
  wire  _T_2635 = btb_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_2904 = _T_2635 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3159 = _T_3158 | _T_2904; // @[Mux.scala 27:72]
  wire  _T_2637 = btb_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_2905 = _T_2637 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3160 = _T_3159 | _T_2905; // @[Mux.scala 27:72]
  wire  _T_2639 = btb_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_2906 = _T_2639 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3161 = _T_3160 | _T_2906; // @[Mux.scala 27:72]
  wire  _T_2641 = btb_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_2907 = _T_2641 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3162 = _T_3161 | _T_2907; // @[Mux.scala 27:72]
  wire  _T_2643 = btb_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_2908 = _T_2643 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3163 = _T_3162 | _T_2908; // @[Mux.scala 27:72]
  wire  _T_2645 = btb_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_2909 = _T_2645 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3164 = _T_3163 | _T_2909; // @[Mux.scala 27:72]
  wire  _T_2647 = btb_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_2910 = _T_2647 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3165 = _T_3164 | _T_2910; // @[Mux.scala 27:72]
  wire  _T_2649 = btb_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_2911 = _T_2649 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3166 = _T_3165 | _T_2911; // @[Mux.scala 27:72]
  wire  _T_2651 = btb_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_2912 = _T_2651 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3167 = _T_3166 | _T_2912; // @[Mux.scala 27:72]
  wire  _T_2653 = btb_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_2913 = _T_2653 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3168 = _T_3167 | _T_2913; // @[Mux.scala 27:72]
  wire  _T_2655 = btb_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_2914 = _T_2655 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3169 = _T_3168 | _T_2914; // @[Mux.scala 27:72]
  wire  _T_2657 = btb_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_2915 = _T_2657 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3170 = _T_3169 | _T_2915; // @[Mux.scala 27:72]
  wire  _T_2659 = btb_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 435:80]
  reg [21:0] btb_bank0_rd_data_way0_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_2916 = _T_2659 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3171 = _T_3170 | _T_2916; // @[Mux.scala 27:72]
  wire [21:0] _T_3172 = _T_3171; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3171; // @[ifu_bp_ctl.scala 435:28]
  wire [4:0] _T_29 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_f = _T_29 ^ io_ifc_fetch_addr_f[23:19]; // @[lib.scala 42:111]
  wire  _T_46 = _T_3172[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 144:98]
  wire  _T_47 = _T_3172[0] & _T_46; // @[ifu_bp_ctl.scala 144:55]
  wire  _T_19 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_f; // @[ifu_bp_ctl.scala 125:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[ifu_bp_ctl.scala 125:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 129:63]
  wire  _T_48 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & branch_error_bank_conflict_f; // @[ifu_bp_ctl.scala 145:22]
  wire  _T_49 = ~_T_48; // @[ifu_bp_ctl.scala 145:5]
  wire  _T_50 = _T_47 & _T_49; // @[ifu_bp_ctl.scala 144:118]
  wire  _T_51 = _T_50 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 145:54]
  wire  tag_match_way0_f = _T_51 & _T; // @[ifu_bp_ctl.scala 145:75]
  wire  _T_82 = _T_3172[3] ^ _T_3172[4]; // @[ifu_bp_ctl.scala 159:90]
  wire  _T_83 = tag_match_way0_f & _T_82; // @[ifu_bp_ctl.scala 159:56]
  wire  _T_87 = ~_T_82; // @[ifu_bp_ctl.scala 160:24]
  wire  _T_88 = tag_match_way0_f & _T_87; // @[ifu_bp_ctl.scala 160:22]
  wire [1:0] tag_match_way0_expanded_f = {_T_83,_T_88}; // @[Cat.scala 29:58]
  wire [21:0] _T_129 = tag_match_way0_expanded_f[1] ? _T_3172 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_3685 = _T_2149 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_3686 = _T_2151 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3941 = _T_3685 | _T_3686; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_3687 = _T_2153 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3942 = _T_3941 | _T_3687; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_3688 = _T_2155 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3943 = _T_3942 | _T_3688; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_3689 = _T_2157 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3944 = _T_3943 | _T_3689; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_3690 = _T_2159 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3945 = _T_3944 | _T_3690; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_3691 = _T_2161 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3946 = _T_3945 | _T_3691; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_3692 = _T_2163 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3947 = _T_3946 | _T_3692; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_3693 = _T_2165 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3948 = _T_3947 | _T_3693; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_3694 = _T_2167 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3949 = _T_3948 | _T_3694; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_3695 = _T_2169 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3950 = _T_3949 | _T_3695; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_3696 = _T_2171 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3951 = _T_3950 | _T_3696; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_3697 = _T_2173 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3952 = _T_3951 | _T_3697; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_3698 = _T_2175 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3953 = _T_3952 | _T_3698; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_3699 = _T_2177 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3954 = _T_3953 | _T_3699; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_3700 = _T_2179 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3955 = _T_3954 | _T_3700; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_3701 = _T_2181 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3956 = _T_3955 | _T_3701; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_3702 = _T_2183 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3957 = _T_3956 | _T_3702; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_3703 = _T_2185 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3958 = _T_3957 | _T_3703; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_3704 = _T_2187 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3959 = _T_3958 | _T_3704; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_3705 = _T_2189 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3960 = _T_3959 | _T_3705; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_3706 = _T_2191 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3961 = _T_3960 | _T_3706; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_3707 = _T_2193 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3962 = _T_3961 | _T_3707; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_3708 = _T_2195 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3963 = _T_3962 | _T_3708; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_3709 = _T_2197 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3964 = _T_3963 | _T_3709; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_3710 = _T_2199 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3965 = _T_3964 | _T_3710; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_3711 = _T_2201 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3966 = _T_3965 | _T_3711; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_3712 = _T_2203 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3967 = _T_3966 | _T_3712; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_3713 = _T_2205 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3968 = _T_3967 | _T_3713; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_3714 = _T_2207 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3969 = _T_3968 | _T_3714; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_3715 = _T_2209 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3970 = _T_3969 | _T_3715; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_3716 = _T_2211 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3971 = _T_3970 | _T_3716; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_3717 = _T_2213 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3972 = _T_3971 | _T_3717; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_3718 = _T_2215 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3973 = _T_3972 | _T_3718; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_3719 = _T_2217 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3974 = _T_3973 | _T_3719; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_3720 = _T_2219 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3975 = _T_3974 | _T_3720; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_3721 = _T_2221 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3976 = _T_3975 | _T_3721; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_3722 = _T_2223 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3977 = _T_3976 | _T_3722; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_3723 = _T_2225 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3978 = _T_3977 | _T_3723; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_3724 = _T_2227 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3979 = _T_3978 | _T_3724; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_3725 = _T_2229 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3980 = _T_3979 | _T_3725; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_3726 = _T_2231 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3981 = _T_3980 | _T_3726; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_3727 = _T_2233 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3982 = _T_3981 | _T_3727; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_3728 = _T_2235 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3983 = _T_3982 | _T_3728; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_3729 = _T_2237 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3984 = _T_3983 | _T_3729; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_3730 = _T_2239 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3985 = _T_3984 | _T_3730; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_3731 = _T_2241 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3986 = _T_3985 | _T_3731; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_3732 = _T_2243 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3987 = _T_3986 | _T_3732; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_3733 = _T_2245 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3988 = _T_3987 | _T_3733; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_3734 = _T_2247 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3989 = _T_3988 | _T_3734; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_3735 = _T_2249 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3990 = _T_3989 | _T_3735; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_3736 = _T_2251 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3991 = _T_3990 | _T_3736; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_3737 = _T_2253 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3992 = _T_3991 | _T_3737; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_3738 = _T_2255 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3993 = _T_3992 | _T_3738; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_3739 = _T_2257 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3994 = _T_3993 | _T_3739; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_3740 = _T_2259 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3995 = _T_3994 | _T_3740; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_3741 = _T_2261 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3996 = _T_3995 | _T_3741; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_3742 = _T_2263 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3997 = _T_3996 | _T_3742; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_3743 = _T_2265 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3998 = _T_3997 | _T_3743; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_3744 = _T_2267 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3999 = _T_3998 | _T_3744; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_3745 = _T_2269 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4000 = _T_3999 | _T_3745; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_3746 = _T_2271 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4001 = _T_4000 | _T_3746; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_3747 = _T_2273 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4002 = _T_4001 | _T_3747; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_3748 = _T_2275 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4003 = _T_4002 | _T_3748; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_3749 = _T_2277 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4004 = _T_4003 | _T_3749; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_3750 = _T_2279 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4005 = _T_4004 | _T_3750; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_3751 = _T_2281 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4006 = _T_4005 | _T_3751; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_3752 = _T_2283 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4007 = _T_4006 | _T_3752; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_3753 = _T_2285 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4008 = _T_4007 | _T_3753; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_3754 = _T_2287 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4009 = _T_4008 | _T_3754; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_3755 = _T_2289 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4010 = _T_4009 | _T_3755; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_3756 = _T_2291 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4011 = _T_4010 | _T_3756; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_3757 = _T_2293 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4012 = _T_4011 | _T_3757; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_3758 = _T_2295 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4013 = _T_4012 | _T_3758; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_3759 = _T_2297 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4014 = _T_4013 | _T_3759; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_3760 = _T_2299 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4015 = _T_4014 | _T_3760; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_3761 = _T_2301 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4016 = _T_4015 | _T_3761; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_3762 = _T_2303 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4017 = _T_4016 | _T_3762; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_3763 = _T_2305 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4018 = _T_4017 | _T_3763; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_3764 = _T_2307 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4019 = _T_4018 | _T_3764; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_3765 = _T_2309 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4020 = _T_4019 | _T_3765; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_3766 = _T_2311 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4021 = _T_4020 | _T_3766; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_3767 = _T_2313 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4022 = _T_4021 | _T_3767; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_3768 = _T_2315 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4023 = _T_4022 | _T_3768; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_3769 = _T_2317 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4024 = _T_4023 | _T_3769; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_3770 = _T_2319 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4025 = _T_4024 | _T_3770; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_3771 = _T_2321 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4026 = _T_4025 | _T_3771; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_3772 = _T_2323 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4027 = _T_4026 | _T_3772; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_3773 = _T_2325 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4028 = _T_4027 | _T_3773; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_3774 = _T_2327 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4029 = _T_4028 | _T_3774; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_3775 = _T_2329 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4030 = _T_4029 | _T_3775; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_3776 = _T_2331 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4031 = _T_4030 | _T_3776; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_3777 = _T_2333 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4032 = _T_4031 | _T_3777; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_3778 = _T_2335 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4033 = _T_4032 | _T_3778; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_3779 = _T_2337 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4034 = _T_4033 | _T_3779; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_3780 = _T_2339 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4035 = _T_4034 | _T_3780; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_3781 = _T_2341 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4036 = _T_4035 | _T_3781; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_3782 = _T_2343 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4037 = _T_4036 | _T_3782; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_3783 = _T_2345 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4038 = _T_4037 | _T_3783; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_3784 = _T_2347 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4039 = _T_4038 | _T_3784; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_3785 = _T_2349 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4040 = _T_4039 | _T_3785; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_3786 = _T_2351 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4041 = _T_4040 | _T_3786; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_3787 = _T_2353 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4042 = _T_4041 | _T_3787; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_3788 = _T_2355 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4043 = _T_4042 | _T_3788; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_3789 = _T_2357 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4044 = _T_4043 | _T_3789; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_3790 = _T_2359 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4045 = _T_4044 | _T_3790; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_3791 = _T_2361 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4046 = _T_4045 | _T_3791; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_3792 = _T_2363 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4047 = _T_4046 | _T_3792; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_3793 = _T_2365 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4048 = _T_4047 | _T_3793; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_3794 = _T_2367 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4049 = _T_4048 | _T_3794; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_3795 = _T_2369 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4050 = _T_4049 | _T_3795; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_3796 = _T_2371 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4051 = _T_4050 | _T_3796; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_3797 = _T_2373 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4052 = _T_4051 | _T_3797; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_3798 = _T_2375 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4053 = _T_4052 | _T_3798; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_3799 = _T_2377 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4054 = _T_4053 | _T_3799; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_3800 = _T_2379 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4055 = _T_4054 | _T_3800; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_3801 = _T_2381 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4056 = _T_4055 | _T_3801; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_3802 = _T_2383 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4057 = _T_4056 | _T_3802; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_3803 = _T_2385 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4058 = _T_4057 | _T_3803; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_3804 = _T_2387 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4059 = _T_4058 | _T_3804; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_3805 = _T_2389 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4060 = _T_4059 | _T_3805; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_3806 = _T_2391 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4061 = _T_4060 | _T_3806; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_3807 = _T_2393 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4062 = _T_4061 | _T_3807; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_3808 = _T_2395 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4063 = _T_4062 | _T_3808; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_3809 = _T_2397 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4064 = _T_4063 | _T_3809; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_3810 = _T_2399 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4065 = _T_4064 | _T_3810; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_3811 = _T_2401 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4066 = _T_4065 | _T_3811; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_3812 = _T_2403 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4067 = _T_4066 | _T_3812; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_3813 = _T_2405 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4068 = _T_4067 | _T_3813; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_3814 = _T_2407 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4069 = _T_4068 | _T_3814; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_3815 = _T_2409 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4070 = _T_4069 | _T_3815; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_3816 = _T_2411 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4071 = _T_4070 | _T_3816; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_3817 = _T_2413 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4072 = _T_4071 | _T_3817; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_3818 = _T_2415 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4073 = _T_4072 | _T_3818; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_3819 = _T_2417 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4074 = _T_4073 | _T_3819; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_3820 = _T_2419 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4075 = _T_4074 | _T_3820; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_3821 = _T_2421 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4076 = _T_4075 | _T_3821; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_3822 = _T_2423 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4077 = _T_4076 | _T_3822; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_3823 = _T_2425 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4078 = _T_4077 | _T_3823; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_3824 = _T_2427 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4079 = _T_4078 | _T_3824; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_3825 = _T_2429 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4080 = _T_4079 | _T_3825; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_3826 = _T_2431 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4081 = _T_4080 | _T_3826; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_3827 = _T_2433 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4082 = _T_4081 | _T_3827; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_3828 = _T_2435 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4083 = _T_4082 | _T_3828; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_3829 = _T_2437 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4084 = _T_4083 | _T_3829; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_3830 = _T_2439 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4085 = _T_4084 | _T_3830; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_3831 = _T_2441 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4086 = _T_4085 | _T_3831; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_3832 = _T_2443 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4087 = _T_4086 | _T_3832; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_3833 = _T_2445 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4088 = _T_4087 | _T_3833; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_3834 = _T_2447 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4089 = _T_4088 | _T_3834; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_3835 = _T_2449 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4090 = _T_4089 | _T_3835; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_3836 = _T_2451 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4091 = _T_4090 | _T_3836; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_3837 = _T_2453 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4092 = _T_4091 | _T_3837; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_3838 = _T_2455 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4093 = _T_4092 | _T_3838; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_3839 = _T_2457 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4094 = _T_4093 | _T_3839; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_3840 = _T_2459 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4095 = _T_4094 | _T_3840; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_3841 = _T_2461 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4096 = _T_4095 | _T_3841; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_3842 = _T_2463 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4097 = _T_4096 | _T_3842; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_3843 = _T_2465 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4098 = _T_4097 | _T_3843; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_3844 = _T_2467 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4099 = _T_4098 | _T_3844; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_3845 = _T_2469 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4100 = _T_4099 | _T_3845; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_3846 = _T_2471 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4101 = _T_4100 | _T_3846; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_3847 = _T_2473 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4102 = _T_4101 | _T_3847; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_3848 = _T_2475 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4103 = _T_4102 | _T_3848; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_3849 = _T_2477 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4104 = _T_4103 | _T_3849; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_3850 = _T_2479 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4105 = _T_4104 | _T_3850; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_3851 = _T_2481 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4106 = _T_4105 | _T_3851; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_3852 = _T_2483 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4107 = _T_4106 | _T_3852; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_3853 = _T_2485 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4108 = _T_4107 | _T_3853; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_3854 = _T_2487 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4109 = _T_4108 | _T_3854; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_3855 = _T_2489 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4110 = _T_4109 | _T_3855; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_3856 = _T_2491 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4111 = _T_4110 | _T_3856; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_3857 = _T_2493 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4112 = _T_4111 | _T_3857; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_3858 = _T_2495 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4113 = _T_4112 | _T_3858; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_3859 = _T_2497 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4114 = _T_4113 | _T_3859; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_3860 = _T_2499 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4115 = _T_4114 | _T_3860; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_3861 = _T_2501 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4116 = _T_4115 | _T_3861; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_3862 = _T_2503 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4117 = _T_4116 | _T_3862; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_3863 = _T_2505 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4118 = _T_4117 | _T_3863; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_3864 = _T_2507 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4119 = _T_4118 | _T_3864; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_3865 = _T_2509 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4120 = _T_4119 | _T_3865; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_3866 = _T_2511 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4121 = _T_4120 | _T_3866; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_3867 = _T_2513 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4122 = _T_4121 | _T_3867; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_3868 = _T_2515 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4123 = _T_4122 | _T_3868; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_3869 = _T_2517 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4124 = _T_4123 | _T_3869; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_3870 = _T_2519 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4125 = _T_4124 | _T_3870; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_3871 = _T_2521 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4126 = _T_4125 | _T_3871; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_3872 = _T_2523 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4127 = _T_4126 | _T_3872; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_3873 = _T_2525 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4128 = _T_4127 | _T_3873; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_3874 = _T_2527 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4129 = _T_4128 | _T_3874; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_3875 = _T_2529 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4130 = _T_4129 | _T_3875; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_3876 = _T_2531 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4131 = _T_4130 | _T_3876; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_3877 = _T_2533 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4132 = _T_4131 | _T_3877; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_3878 = _T_2535 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4133 = _T_4132 | _T_3878; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_3879 = _T_2537 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4134 = _T_4133 | _T_3879; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_3880 = _T_2539 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4135 = _T_4134 | _T_3880; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_3881 = _T_2541 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4136 = _T_4135 | _T_3881; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_3882 = _T_2543 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4137 = _T_4136 | _T_3882; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_3883 = _T_2545 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4138 = _T_4137 | _T_3883; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_3884 = _T_2547 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4139 = _T_4138 | _T_3884; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_3885 = _T_2549 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4140 = _T_4139 | _T_3885; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_3886 = _T_2551 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4141 = _T_4140 | _T_3886; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_3887 = _T_2553 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4142 = _T_4141 | _T_3887; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_3888 = _T_2555 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4143 = _T_4142 | _T_3888; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_3889 = _T_2557 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4144 = _T_4143 | _T_3889; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_3890 = _T_2559 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4145 = _T_4144 | _T_3890; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_3891 = _T_2561 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4146 = _T_4145 | _T_3891; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_3892 = _T_2563 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4147 = _T_4146 | _T_3892; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_3893 = _T_2565 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4148 = _T_4147 | _T_3893; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_3894 = _T_2567 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4149 = _T_4148 | _T_3894; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_3895 = _T_2569 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4150 = _T_4149 | _T_3895; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_3896 = _T_2571 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4151 = _T_4150 | _T_3896; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_3897 = _T_2573 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4152 = _T_4151 | _T_3897; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_3898 = _T_2575 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4153 = _T_4152 | _T_3898; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_3899 = _T_2577 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4154 = _T_4153 | _T_3899; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_3900 = _T_2579 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4155 = _T_4154 | _T_3900; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_3901 = _T_2581 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4156 = _T_4155 | _T_3901; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_3902 = _T_2583 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4157 = _T_4156 | _T_3902; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_3903 = _T_2585 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4158 = _T_4157 | _T_3903; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_3904 = _T_2587 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4159 = _T_4158 | _T_3904; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_3905 = _T_2589 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4160 = _T_4159 | _T_3905; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_3906 = _T_2591 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4161 = _T_4160 | _T_3906; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_3907 = _T_2593 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4162 = _T_4161 | _T_3907; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_3908 = _T_2595 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4163 = _T_4162 | _T_3908; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_3909 = _T_2597 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4164 = _T_4163 | _T_3909; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_3910 = _T_2599 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4165 = _T_4164 | _T_3910; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_3911 = _T_2601 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4166 = _T_4165 | _T_3911; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_3912 = _T_2603 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4167 = _T_4166 | _T_3912; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_3913 = _T_2605 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4168 = _T_4167 | _T_3913; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_3914 = _T_2607 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4169 = _T_4168 | _T_3914; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_3915 = _T_2609 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4170 = _T_4169 | _T_3915; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_3916 = _T_2611 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4171 = _T_4170 | _T_3916; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_3917 = _T_2613 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4172 = _T_4171 | _T_3917; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_3918 = _T_2615 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4173 = _T_4172 | _T_3918; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_3919 = _T_2617 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4174 = _T_4173 | _T_3919; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_3920 = _T_2619 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4175 = _T_4174 | _T_3920; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_3921 = _T_2621 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4176 = _T_4175 | _T_3921; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_3922 = _T_2623 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4177 = _T_4176 | _T_3922; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_3923 = _T_2625 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4178 = _T_4177 | _T_3923; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_3924 = _T_2627 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4179 = _T_4178 | _T_3924; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_3925 = _T_2629 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4180 = _T_4179 | _T_3925; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_3926 = _T_2631 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4181 = _T_4180 | _T_3926; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_3927 = _T_2633 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4182 = _T_4181 | _T_3927; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_3928 = _T_2635 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4183 = _T_4182 | _T_3928; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_3929 = _T_2637 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4184 = _T_4183 | _T_3929; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_3930 = _T_2639 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4185 = _T_4184 | _T_3930; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_3931 = _T_2641 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4186 = _T_4185 | _T_3931; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_3932 = _T_2643 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4187 = _T_4186 | _T_3932; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_3933 = _T_2645 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4188 = _T_4187 | _T_3933; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_3934 = _T_2647 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4189 = _T_4188 | _T_3934; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_3935 = _T_2649 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4190 = _T_4189 | _T_3935; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_3936 = _T_2651 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4191 = _T_4190 | _T_3936; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_3937 = _T_2653 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4192 = _T_4191 | _T_3937; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_3938 = _T_2655 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4193 = _T_4192 | _T_3938; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_3939 = _T_2657 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4194 = _T_4193 | _T_3939; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_3940 = _T_2659 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4195 = _T_4194 | _T_3940; // @[Mux.scala 27:72]
  wire [21:0] _T_4196 = _T_4195; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4195; // @[ifu_bp_ctl.scala 438:28]
  wire  _T_55 = _T_4196[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 148:98]
  wire  _T_56 = _T_4196[0] & _T_55; // @[ifu_bp_ctl.scala 148:55]
  wire  _T_59 = _T_56 & _T_49; // @[ifu_bp_ctl.scala 148:118]
  wire  _T_60 = _T_59 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 149:54]
  wire  tag_match_way1_f = _T_60 & _T; // @[ifu_bp_ctl.scala 149:75]
  wire  _T_91 = _T_4196[3] ^ _T_4196[4]; // @[ifu_bp_ctl.scala 162:90]
  wire  _T_92 = tag_match_way1_f & _T_91; // @[ifu_bp_ctl.scala 162:56]
  wire  _T_96 = ~_T_91; // @[ifu_bp_ctl.scala 163:24]
  wire  _T_97 = tag_match_way1_f & _T_96; // @[ifu_bp_ctl.scala 163:22]
  wire [1:0] tag_match_way1_expanded_f = {_T_92,_T_97}; // @[Cat.scala 29:58]
  wire [21:0] _T_130 = tag_match_way1_expanded_f[1] ? _T_4196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0o_rd_data_f = _T_129 | _T_130; // @[Mux.scala 27:72]
  wire [21:0] _T_149 = _T_147 ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4197 = btb_rd_addr_p1_f == 8'h0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4709 = _T_4197 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4199 = btb_rd_addr_p1_f == 8'h1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4710 = _T_4199 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4965 = _T_4709 | _T_4710; // @[Mux.scala 27:72]
  wire  _T_4201 = btb_rd_addr_p1_f == 8'h2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4711 = _T_4201 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4966 = _T_4965 | _T_4711; // @[Mux.scala 27:72]
  wire  _T_4203 = btb_rd_addr_p1_f == 8'h3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4712 = _T_4203 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4967 = _T_4966 | _T_4712; // @[Mux.scala 27:72]
  wire  _T_4205 = btb_rd_addr_p1_f == 8'h4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4713 = _T_4205 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4968 = _T_4967 | _T_4713; // @[Mux.scala 27:72]
  wire  _T_4207 = btb_rd_addr_p1_f == 8'h5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4714 = _T_4207 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4969 = _T_4968 | _T_4714; // @[Mux.scala 27:72]
  wire  _T_4209 = btb_rd_addr_p1_f == 8'h6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4715 = _T_4209 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4970 = _T_4969 | _T_4715; // @[Mux.scala 27:72]
  wire  _T_4211 = btb_rd_addr_p1_f == 8'h7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4716 = _T_4211 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4971 = _T_4970 | _T_4716; // @[Mux.scala 27:72]
  wire  _T_4213 = btb_rd_addr_p1_f == 8'h8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4717 = _T_4213 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4972 = _T_4971 | _T_4717; // @[Mux.scala 27:72]
  wire  _T_4215 = btb_rd_addr_p1_f == 8'h9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4718 = _T_4215 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4973 = _T_4972 | _T_4718; // @[Mux.scala 27:72]
  wire  _T_4217 = btb_rd_addr_p1_f == 8'ha; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4719 = _T_4217 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4974 = _T_4973 | _T_4719; // @[Mux.scala 27:72]
  wire  _T_4219 = btb_rd_addr_p1_f == 8'hb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4720 = _T_4219 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4975 = _T_4974 | _T_4720; // @[Mux.scala 27:72]
  wire  _T_4221 = btb_rd_addr_p1_f == 8'hc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4721 = _T_4221 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4976 = _T_4975 | _T_4721; // @[Mux.scala 27:72]
  wire  _T_4223 = btb_rd_addr_p1_f == 8'hd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4722 = _T_4223 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4977 = _T_4976 | _T_4722; // @[Mux.scala 27:72]
  wire  _T_4225 = btb_rd_addr_p1_f == 8'he; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4723 = _T_4225 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4978 = _T_4977 | _T_4723; // @[Mux.scala 27:72]
  wire  _T_4227 = btb_rd_addr_p1_f == 8'hf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4724 = _T_4227 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4979 = _T_4978 | _T_4724; // @[Mux.scala 27:72]
  wire  _T_4229 = btb_rd_addr_p1_f == 8'h10; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4725 = _T_4229 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4980 = _T_4979 | _T_4725; // @[Mux.scala 27:72]
  wire  _T_4231 = btb_rd_addr_p1_f == 8'h11; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4726 = _T_4231 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4981 = _T_4980 | _T_4726; // @[Mux.scala 27:72]
  wire  _T_4233 = btb_rd_addr_p1_f == 8'h12; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4727 = _T_4233 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4982 = _T_4981 | _T_4727; // @[Mux.scala 27:72]
  wire  _T_4235 = btb_rd_addr_p1_f == 8'h13; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4728 = _T_4235 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4983 = _T_4982 | _T_4728; // @[Mux.scala 27:72]
  wire  _T_4237 = btb_rd_addr_p1_f == 8'h14; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4729 = _T_4237 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4984 = _T_4983 | _T_4729; // @[Mux.scala 27:72]
  wire  _T_4239 = btb_rd_addr_p1_f == 8'h15; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4730 = _T_4239 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4985 = _T_4984 | _T_4730; // @[Mux.scala 27:72]
  wire  _T_4241 = btb_rd_addr_p1_f == 8'h16; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4731 = _T_4241 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4986 = _T_4985 | _T_4731; // @[Mux.scala 27:72]
  wire  _T_4243 = btb_rd_addr_p1_f == 8'h17; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4732 = _T_4243 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4987 = _T_4986 | _T_4732; // @[Mux.scala 27:72]
  wire  _T_4245 = btb_rd_addr_p1_f == 8'h18; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4733 = _T_4245 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4988 = _T_4987 | _T_4733; // @[Mux.scala 27:72]
  wire  _T_4247 = btb_rd_addr_p1_f == 8'h19; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4734 = _T_4247 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4989 = _T_4988 | _T_4734; // @[Mux.scala 27:72]
  wire  _T_4249 = btb_rd_addr_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4735 = _T_4249 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4990 = _T_4989 | _T_4735; // @[Mux.scala 27:72]
  wire  _T_4251 = btb_rd_addr_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4736 = _T_4251 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4991 = _T_4990 | _T_4736; // @[Mux.scala 27:72]
  wire  _T_4253 = btb_rd_addr_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4737 = _T_4253 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4992 = _T_4991 | _T_4737; // @[Mux.scala 27:72]
  wire  _T_4255 = btb_rd_addr_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4738 = _T_4255 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4993 = _T_4992 | _T_4738; // @[Mux.scala 27:72]
  wire  _T_4257 = btb_rd_addr_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4739 = _T_4257 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4994 = _T_4993 | _T_4739; // @[Mux.scala 27:72]
  wire  _T_4259 = btb_rd_addr_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4740 = _T_4259 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4995 = _T_4994 | _T_4740; // @[Mux.scala 27:72]
  wire  _T_4261 = btb_rd_addr_p1_f == 8'h20; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4741 = _T_4261 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4996 = _T_4995 | _T_4741; // @[Mux.scala 27:72]
  wire  _T_4263 = btb_rd_addr_p1_f == 8'h21; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4742 = _T_4263 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4997 = _T_4996 | _T_4742; // @[Mux.scala 27:72]
  wire  _T_4265 = btb_rd_addr_p1_f == 8'h22; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4743 = _T_4265 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4998 = _T_4997 | _T_4743; // @[Mux.scala 27:72]
  wire  _T_4267 = btb_rd_addr_p1_f == 8'h23; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4744 = _T_4267 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4999 = _T_4998 | _T_4744; // @[Mux.scala 27:72]
  wire  _T_4269 = btb_rd_addr_p1_f == 8'h24; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4745 = _T_4269 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5000 = _T_4999 | _T_4745; // @[Mux.scala 27:72]
  wire  _T_4271 = btb_rd_addr_p1_f == 8'h25; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4746 = _T_4271 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5001 = _T_5000 | _T_4746; // @[Mux.scala 27:72]
  wire  _T_4273 = btb_rd_addr_p1_f == 8'h26; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4747 = _T_4273 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5002 = _T_5001 | _T_4747; // @[Mux.scala 27:72]
  wire  _T_4275 = btb_rd_addr_p1_f == 8'h27; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4748 = _T_4275 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5003 = _T_5002 | _T_4748; // @[Mux.scala 27:72]
  wire  _T_4277 = btb_rd_addr_p1_f == 8'h28; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4749 = _T_4277 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5004 = _T_5003 | _T_4749; // @[Mux.scala 27:72]
  wire  _T_4279 = btb_rd_addr_p1_f == 8'h29; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4750 = _T_4279 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5005 = _T_5004 | _T_4750; // @[Mux.scala 27:72]
  wire  _T_4281 = btb_rd_addr_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4751 = _T_4281 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5006 = _T_5005 | _T_4751; // @[Mux.scala 27:72]
  wire  _T_4283 = btb_rd_addr_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4752 = _T_4283 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5007 = _T_5006 | _T_4752; // @[Mux.scala 27:72]
  wire  _T_4285 = btb_rd_addr_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4753 = _T_4285 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5008 = _T_5007 | _T_4753; // @[Mux.scala 27:72]
  wire  _T_4287 = btb_rd_addr_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4754 = _T_4287 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5009 = _T_5008 | _T_4754; // @[Mux.scala 27:72]
  wire  _T_4289 = btb_rd_addr_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4755 = _T_4289 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5010 = _T_5009 | _T_4755; // @[Mux.scala 27:72]
  wire  _T_4291 = btb_rd_addr_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4756 = _T_4291 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5011 = _T_5010 | _T_4756; // @[Mux.scala 27:72]
  wire  _T_4293 = btb_rd_addr_p1_f == 8'h30; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4757 = _T_4293 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5012 = _T_5011 | _T_4757; // @[Mux.scala 27:72]
  wire  _T_4295 = btb_rd_addr_p1_f == 8'h31; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4758 = _T_4295 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5013 = _T_5012 | _T_4758; // @[Mux.scala 27:72]
  wire  _T_4297 = btb_rd_addr_p1_f == 8'h32; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4759 = _T_4297 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5014 = _T_5013 | _T_4759; // @[Mux.scala 27:72]
  wire  _T_4299 = btb_rd_addr_p1_f == 8'h33; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4760 = _T_4299 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5015 = _T_5014 | _T_4760; // @[Mux.scala 27:72]
  wire  _T_4301 = btb_rd_addr_p1_f == 8'h34; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4761 = _T_4301 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5016 = _T_5015 | _T_4761; // @[Mux.scala 27:72]
  wire  _T_4303 = btb_rd_addr_p1_f == 8'h35; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4762 = _T_4303 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5017 = _T_5016 | _T_4762; // @[Mux.scala 27:72]
  wire  _T_4305 = btb_rd_addr_p1_f == 8'h36; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4763 = _T_4305 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5018 = _T_5017 | _T_4763; // @[Mux.scala 27:72]
  wire  _T_4307 = btb_rd_addr_p1_f == 8'h37; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4764 = _T_4307 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5019 = _T_5018 | _T_4764; // @[Mux.scala 27:72]
  wire  _T_4309 = btb_rd_addr_p1_f == 8'h38; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4765 = _T_4309 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5020 = _T_5019 | _T_4765; // @[Mux.scala 27:72]
  wire  _T_4311 = btb_rd_addr_p1_f == 8'h39; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4766 = _T_4311 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5021 = _T_5020 | _T_4766; // @[Mux.scala 27:72]
  wire  _T_4313 = btb_rd_addr_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4767 = _T_4313 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5022 = _T_5021 | _T_4767; // @[Mux.scala 27:72]
  wire  _T_4315 = btb_rd_addr_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4768 = _T_4315 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5023 = _T_5022 | _T_4768; // @[Mux.scala 27:72]
  wire  _T_4317 = btb_rd_addr_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4769 = _T_4317 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5024 = _T_5023 | _T_4769; // @[Mux.scala 27:72]
  wire  _T_4319 = btb_rd_addr_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4770 = _T_4319 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5025 = _T_5024 | _T_4770; // @[Mux.scala 27:72]
  wire  _T_4321 = btb_rd_addr_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4771 = _T_4321 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5026 = _T_5025 | _T_4771; // @[Mux.scala 27:72]
  wire  _T_4323 = btb_rd_addr_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4772 = _T_4323 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5027 = _T_5026 | _T_4772; // @[Mux.scala 27:72]
  wire  _T_4325 = btb_rd_addr_p1_f == 8'h40; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4773 = _T_4325 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5028 = _T_5027 | _T_4773; // @[Mux.scala 27:72]
  wire  _T_4327 = btb_rd_addr_p1_f == 8'h41; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4774 = _T_4327 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5029 = _T_5028 | _T_4774; // @[Mux.scala 27:72]
  wire  _T_4329 = btb_rd_addr_p1_f == 8'h42; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4775 = _T_4329 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5030 = _T_5029 | _T_4775; // @[Mux.scala 27:72]
  wire  _T_4331 = btb_rd_addr_p1_f == 8'h43; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4776 = _T_4331 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5031 = _T_5030 | _T_4776; // @[Mux.scala 27:72]
  wire  _T_4333 = btb_rd_addr_p1_f == 8'h44; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4777 = _T_4333 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5032 = _T_5031 | _T_4777; // @[Mux.scala 27:72]
  wire  _T_4335 = btb_rd_addr_p1_f == 8'h45; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4778 = _T_4335 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5033 = _T_5032 | _T_4778; // @[Mux.scala 27:72]
  wire  _T_4337 = btb_rd_addr_p1_f == 8'h46; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4779 = _T_4337 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5034 = _T_5033 | _T_4779; // @[Mux.scala 27:72]
  wire  _T_4339 = btb_rd_addr_p1_f == 8'h47; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4780 = _T_4339 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5035 = _T_5034 | _T_4780; // @[Mux.scala 27:72]
  wire  _T_4341 = btb_rd_addr_p1_f == 8'h48; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4781 = _T_4341 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5036 = _T_5035 | _T_4781; // @[Mux.scala 27:72]
  wire  _T_4343 = btb_rd_addr_p1_f == 8'h49; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4782 = _T_4343 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5037 = _T_5036 | _T_4782; // @[Mux.scala 27:72]
  wire  _T_4345 = btb_rd_addr_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4783 = _T_4345 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5038 = _T_5037 | _T_4783; // @[Mux.scala 27:72]
  wire  _T_4347 = btb_rd_addr_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4784 = _T_4347 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5039 = _T_5038 | _T_4784; // @[Mux.scala 27:72]
  wire  _T_4349 = btb_rd_addr_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4785 = _T_4349 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5040 = _T_5039 | _T_4785; // @[Mux.scala 27:72]
  wire  _T_4351 = btb_rd_addr_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4786 = _T_4351 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5041 = _T_5040 | _T_4786; // @[Mux.scala 27:72]
  wire  _T_4353 = btb_rd_addr_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4787 = _T_4353 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5042 = _T_5041 | _T_4787; // @[Mux.scala 27:72]
  wire  _T_4355 = btb_rd_addr_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4788 = _T_4355 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5043 = _T_5042 | _T_4788; // @[Mux.scala 27:72]
  wire  _T_4357 = btb_rd_addr_p1_f == 8'h50; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4789 = _T_4357 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5044 = _T_5043 | _T_4789; // @[Mux.scala 27:72]
  wire  _T_4359 = btb_rd_addr_p1_f == 8'h51; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4790 = _T_4359 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5045 = _T_5044 | _T_4790; // @[Mux.scala 27:72]
  wire  _T_4361 = btb_rd_addr_p1_f == 8'h52; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4791 = _T_4361 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5046 = _T_5045 | _T_4791; // @[Mux.scala 27:72]
  wire  _T_4363 = btb_rd_addr_p1_f == 8'h53; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4792 = _T_4363 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5047 = _T_5046 | _T_4792; // @[Mux.scala 27:72]
  wire  _T_4365 = btb_rd_addr_p1_f == 8'h54; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4793 = _T_4365 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5048 = _T_5047 | _T_4793; // @[Mux.scala 27:72]
  wire  _T_4367 = btb_rd_addr_p1_f == 8'h55; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4794 = _T_4367 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5049 = _T_5048 | _T_4794; // @[Mux.scala 27:72]
  wire  _T_4369 = btb_rd_addr_p1_f == 8'h56; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4795 = _T_4369 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5050 = _T_5049 | _T_4795; // @[Mux.scala 27:72]
  wire  _T_4371 = btb_rd_addr_p1_f == 8'h57; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4796 = _T_4371 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5051 = _T_5050 | _T_4796; // @[Mux.scala 27:72]
  wire  _T_4373 = btb_rd_addr_p1_f == 8'h58; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4797 = _T_4373 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5052 = _T_5051 | _T_4797; // @[Mux.scala 27:72]
  wire  _T_4375 = btb_rd_addr_p1_f == 8'h59; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4798 = _T_4375 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5053 = _T_5052 | _T_4798; // @[Mux.scala 27:72]
  wire  _T_4377 = btb_rd_addr_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4799 = _T_4377 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5054 = _T_5053 | _T_4799; // @[Mux.scala 27:72]
  wire  _T_4379 = btb_rd_addr_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4800 = _T_4379 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5055 = _T_5054 | _T_4800; // @[Mux.scala 27:72]
  wire  _T_4381 = btb_rd_addr_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4801 = _T_4381 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5056 = _T_5055 | _T_4801; // @[Mux.scala 27:72]
  wire  _T_4383 = btb_rd_addr_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4802 = _T_4383 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5057 = _T_5056 | _T_4802; // @[Mux.scala 27:72]
  wire  _T_4385 = btb_rd_addr_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4803 = _T_4385 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5058 = _T_5057 | _T_4803; // @[Mux.scala 27:72]
  wire  _T_4387 = btb_rd_addr_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4804 = _T_4387 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5059 = _T_5058 | _T_4804; // @[Mux.scala 27:72]
  wire  _T_4389 = btb_rd_addr_p1_f == 8'h60; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4805 = _T_4389 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5060 = _T_5059 | _T_4805; // @[Mux.scala 27:72]
  wire  _T_4391 = btb_rd_addr_p1_f == 8'h61; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4806 = _T_4391 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5061 = _T_5060 | _T_4806; // @[Mux.scala 27:72]
  wire  _T_4393 = btb_rd_addr_p1_f == 8'h62; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4807 = _T_4393 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5062 = _T_5061 | _T_4807; // @[Mux.scala 27:72]
  wire  _T_4395 = btb_rd_addr_p1_f == 8'h63; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4808 = _T_4395 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5063 = _T_5062 | _T_4808; // @[Mux.scala 27:72]
  wire  _T_4397 = btb_rd_addr_p1_f == 8'h64; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4809 = _T_4397 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5064 = _T_5063 | _T_4809; // @[Mux.scala 27:72]
  wire  _T_4399 = btb_rd_addr_p1_f == 8'h65; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4810 = _T_4399 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5065 = _T_5064 | _T_4810; // @[Mux.scala 27:72]
  wire  _T_4401 = btb_rd_addr_p1_f == 8'h66; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4811 = _T_4401 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5066 = _T_5065 | _T_4811; // @[Mux.scala 27:72]
  wire  _T_4403 = btb_rd_addr_p1_f == 8'h67; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4812 = _T_4403 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5067 = _T_5066 | _T_4812; // @[Mux.scala 27:72]
  wire  _T_4405 = btb_rd_addr_p1_f == 8'h68; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4813 = _T_4405 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5068 = _T_5067 | _T_4813; // @[Mux.scala 27:72]
  wire  _T_4407 = btb_rd_addr_p1_f == 8'h69; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4814 = _T_4407 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5069 = _T_5068 | _T_4814; // @[Mux.scala 27:72]
  wire  _T_4409 = btb_rd_addr_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4815 = _T_4409 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5070 = _T_5069 | _T_4815; // @[Mux.scala 27:72]
  wire  _T_4411 = btb_rd_addr_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4816 = _T_4411 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5071 = _T_5070 | _T_4816; // @[Mux.scala 27:72]
  wire  _T_4413 = btb_rd_addr_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4817 = _T_4413 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5072 = _T_5071 | _T_4817; // @[Mux.scala 27:72]
  wire  _T_4415 = btb_rd_addr_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4818 = _T_4415 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5073 = _T_5072 | _T_4818; // @[Mux.scala 27:72]
  wire  _T_4417 = btb_rd_addr_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4819 = _T_4417 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5074 = _T_5073 | _T_4819; // @[Mux.scala 27:72]
  wire  _T_4419 = btb_rd_addr_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4820 = _T_4419 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5075 = _T_5074 | _T_4820; // @[Mux.scala 27:72]
  wire  _T_4421 = btb_rd_addr_p1_f == 8'h70; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4821 = _T_4421 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5076 = _T_5075 | _T_4821; // @[Mux.scala 27:72]
  wire  _T_4423 = btb_rd_addr_p1_f == 8'h71; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4822 = _T_4423 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5077 = _T_5076 | _T_4822; // @[Mux.scala 27:72]
  wire  _T_4425 = btb_rd_addr_p1_f == 8'h72; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4823 = _T_4425 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5078 = _T_5077 | _T_4823; // @[Mux.scala 27:72]
  wire  _T_4427 = btb_rd_addr_p1_f == 8'h73; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4824 = _T_4427 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5079 = _T_5078 | _T_4824; // @[Mux.scala 27:72]
  wire  _T_4429 = btb_rd_addr_p1_f == 8'h74; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4825 = _T_4429 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5080 = _T_5079 | _T_4825; // @[Mux.scala 27:72]
  wire  _T_4431 = btb_rd_addr_p1_f == 8'h75; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4826 = _T_4431 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5081 = _T_5080 | _T_4826; // @[Mux.scala 27:72]
  wire  _T_4433 = btb_rd_addr_p1_f == 8'h76; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4827 = _T_4433 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5082 = _T_5081 | _T_4827; // @[Mux.scala 27:72]
  wire  _T_4435 = btb_rd_addr_p1_f == 8'h77; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4828 = _T_4435 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5083 = _T_5082 | _T_4828; // @[Mux.scala 27:72]
  wire  _T_4437 = btb_rd_addr_p1_f == 8'h78; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4829 = _T_4437 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5084 = _T_5083 | _T_4829; // @[Mux.scala 27:72]
  wire  _T_4439 = btb_rd_addr_p1_f == 8'h79; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4830 = _T_4439 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5085 = _T_5084 | _T_4830; // @[Mux.scala 27:72]
  wire  _T_4441 = btb_rd_addr_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4831 = _T_4441 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5086 = _T_5085 | _T_4831; // @[Mux.scala 27:72]
  wire  _T_4443 = btb_rd_addr_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4832 = _T_4443 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5087 = _T_5086 | _T_4832; // @[Mux.scala 27:72]
  wire  _T_4445 = btb_rd_addr_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4833 = _T_4445 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5088 = _T_5087 | _T_4833; // @[Mux.scala 27:72]
  wire  _T_4447 = btb_rd_addr_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4834 = _T_4447 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5089 = _T_5088 | _T_4834; // @[Mux.scala 27:72]
  wire  _T_4449 = btb_rd_addr_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4835 = _T_4449 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5090 = _T_5089 | _T_4835; // @[Mux.scala 27:72]
  wire  _T_4451 = btb_rd_addr_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4836 = _T_4451 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5091 = _T_5090 | _T_4836; // @[Mux.scala 27:72]
  wire  _T_4453 = btb_rd_addr_p1_f == 8'h80; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4837 = _T_4453 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5092 = _T_5091 | _T_4837; // @[Mux.scala 27:72]
  wire  _T_4455 = btb_rd_addr_p1_f == 8'h81; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4838 = _T_4455 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5093 = _T_5092 | _T_4838; // @[Mux.scala 27:72]
  wire  _T_4457 = btb_rd_addr_p1_f == 8'h82; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4839 = _T_4457 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5094 = _T_5093 | _T_4839; // @[Mux.scala 27:72]
  wire  _T_4459 = btb_rd_addr_p1_f == 8'h83; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4840 = _T_4459 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5095 = _T_5094 | _T_4840; // @[Mux.scala 27:72]
  wire  _T_4461 = btb_rd_addr_p1_f == 8'h84; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4841 = _T_4461 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5096 = _T_5095 | _T_4841; // @[Mux.scala 27:72]
  wire  _T_4463 = btb_rd_addr_p1_f == 8'h85; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4842 = _T_4463 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5097 = _T_5096 | _T_4842; // @[Mux.scala 27:72]
  wire  _T_4465 = btb_rd_addr_p1_f == 8'h86; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4843 = _T_4465 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5098 = _T_5097 | _T_4843; // @[Mux.scala 27:72]
  wire  _T_4467 = btb_rd_addr_p1_f == 8'h87; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4844 = _T_4467 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5099 = _T_5098 | _T_4844; // @[Mux.scala 27:72]
  wire  _T_4469 = btb_rd_addr_p1_f == 8'h88; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4845 = _T_4469 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5100 = _T_5099 | _T_4845; // @[Mux.scala 27:72]
  wire  _T_4471 = btb_rd_addr_p1_f == 8'h89; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4846 = _T_4471 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5101 = _T_5100 | _T_4846; // @[Mux.scala 27:72]
  wire  _T_4473 = btb_rd_addr_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4847 = _T_4473 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5102 = _T_5101 | _T_4847; // @[Mux.scala 27:72]
  wire  _T_4475 = btb_rd_addr_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4848 = _T_4475 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5103 = _T_5102 | _T_4848; // @[Mux.scala 27:72]
  wire  _T_4477 = btb_rd_addr_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4849 = _T_4477 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5104 = _T_5103 | _T_4849; // @[Mux.scala 27:72]
  wire  _T_4479 = btb_rd_addr_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4850 = _T_4479 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5105 = _T_5104 | _T_4850; // @[Mux.scala 27:72]
  wire  _T_4481 = btb_rd_addr_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4851 = _T_4481 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5106 = _T_5105 | _T_4851; // @[Mux.scala 27:72]
  wire  _T_4483 = btb_rd_addr_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4852 = _T_4483 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5107 = _T_5106 | _T_4852; // @[Mux.scala 27:72]
  wire  _T_4485 = btb_rd_addr_p1_f == 8'h90; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4853 = _T_4485 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5108 = _T_5107 | _T_4853; // @[Mux.scala 27:72]
  wire  _T_4487 = btb_rd_addr_p1_f == 8'h91; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4854 = _T_4487 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5109 = _T_5108 | _T_4854; // @[Mux.scala 27:72]
  wire  _T_4489 = btb_rd_addr_p1_f == 8'h92; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4855 = _T_4489 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5110 = _T_5109 | _T_4855; // @[Mux.scala 27:72]
  wire  _T_4491 = btb_rd_addr_p1_f == 8'h93; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4856 = _T_4491 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5111 = _T_5110 | _T_4856; // @[Mux.scala 27:72]
  wire  _T_4493 = btb_rd_addr_p1_f == 8'h94; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4857 = _T_4493 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5112 = _T_5111 | _T_4857; // @[Mux.scala 27:72]
  wire  _T_4495 = btb_rd_addr_p1_f == 8'h95; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4858 = _T_4495 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5113 = _T_5112 | _T_4858; // @[Mux.scala 27:72]
  wire  _T_4497 = btb_rd_addr_p1_f == 8'h96; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4859 = _T_4497 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5114 = _T_5113 | _T_4859; // @[Mux.scala 27:72]
  wire  _T_4499 = btb_rd_addr_p1_f == 8'h97; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4860 = _T_4499 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5115 = _T_5114 | _T_4860; // @[Mux.scala 27:72]
  wire  _T_4501 = btb_rd_addr_p1_f == 8'h98; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4861 = _T_4501 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5116 = _T_5115 | _T_4861; // @[Mux.scala 27:72]
  wire  _T_4503 = btb_rd_addr_p1_f == 8'h99; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4862 = _T_4503 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5117 = _T_5116 | _T_4862; // @[Mux.scala 27:72]
  wire  _T_4505 = btb_rd_addr_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4863 = _T_4505 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5118 = _T_5117 | _T_4863; // @[Mux.scala 27:72]
  wire  _T_4507 = btb_rd_addr_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4864 = _T_4507 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5119 = _T_5118 | _T_4864; // @[Mux.scala 27:72]
  wire  _T_4509 = btb_rd_addr_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4865 = _T_4509 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5120 = _T_5119 | _T_4865; // @[Mux.scala 27:72]
  wire  _T_4511 = btb_rd_addr_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4866 = _T_4511 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5121 = _T_5120 | _T_4866; // @[Mux.scala 27:72]
  wire  _T_4513 = btb_rd_addr_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4867 = _T_4513 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5122 = _T_5121 | _T_4867; // @[Mux.scala 27:72]
  wire  _T_4515 = btb_rd_addr_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4868 = _T_4515 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5123 = _T_5122 | _T_4868; // @[Mux.scala 27:72]
  wire  _T_4517 = btb_rd_addr_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4869 = _T_4517 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5124 = _T_5123 | _T_4869; // @[Mux.scala 27:72]
  wire  _T_4519 = btb_rd_addr_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4870 = _T_4519 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5125 = _T_5124 | _T_4870; // @[Mux.scala 27:72]
  wire  _T_4521 = btb_rd_addr_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4871 = _T_4521 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5126 = _T_5125 | _T_4871; // @[Mux.scala 27:72]
  wire  _T_4523 = btb_rd_addr_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4872 = _T_4523 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5127 = _T_5126 | _T_4872; // @[Mux.scala 27:72]
  wire  _T_4525 = btb_rd_addr_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4873 = _T_4525 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5128 = _T_5127 | _T_4873; // @[Mux.scala 27:72]
  wire  _T_4527 = btb_rd_addr_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4874 = _T_4527 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5129 = _T_5128 | _T_4874; // @[Mux.scala 27:72]
  wire  _T_4529 = btb_rd_addr_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4875 = _T_4529 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5130 = _T_5129 | _T_4875; // @[Mux.scala 27:72]
  wire  _T_4531 = btb_rd_addr_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4876 = _T_4531 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5131 = _T_5130 | _T_4876; // @[Mux.scala 27:72]
  wire  _T_4533 = btb_rd_addr_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4877 = _T_4533 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5132 = _T_5131 | _T_4877; // @[Mux.scala 27:72]
  wire  _T_4535 = btb_rd_addr_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4878 = _T_4535 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5133 = _T_5132 | _T_4878; // @[Mux.scala 27:72]
  wire  _T_4537 = btb_rd_addr_p1_f == 8'haa; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4879 = _T_4537 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5134 = _T_5133 | _T_4879; // @[Mux.scala 27:72]
  wire  _T_4539 = btb_rd_addr_p1_f == 8'hab; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4880 = _T_4539 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5135 = _T_5134 | _T_4880; // @[Mux.scala 27:72]
  wire  _T_4541 = btb_rd_addr_p1_f == 8'hac; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4881 = _T_4541 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5136 = _T_5135 | _T_4881; // @[Mux.scala 27:72]
  wire  _T_4543 = btb_rd_addr_p1_f == 8'had; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4882 = _T_4543 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5137 = _T_5136 | _T_4882; // @[Mux.scala 27:72]
  wire  _T_4545 = btb_rd_addr_p1_f == 8'hae; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4883 = _T_4545 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5138 = _T_5137 | _T_4883; // @[Mux.scala 27:72]
  wire  _T_4547 = btb_rd_addr_p1_f == 8'haf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4884 = _T_4547 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5139 = _T_5138 | _T_4884; // @[Mux.scala 27:72]
  wire  _T_4549 = btb_rd_addr_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4885 = _T_4549 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5140 = _T_5139 | _T_4885; // @[Mux.scala 27:72]
  wire  _T_4551 = btb_rd_addr_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4886 = _T_4551 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5141 = _T_5140 | _T_4886; // @[Mux.scala 27:72]
  wire  _T_4553 = btb_rd_addr_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4887 = _T_4553 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5142 = _T_5141 | _T_4887; // @[Mux.scala 27:72]
  wire  _T_4555 = btb_rd_addr_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4888 = _T_4555 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5143 = _T_5142 | _T_4888; // @[Mux.scala 27:72]
  wire  _T_4557 = btb_rd_addr_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4889 = _T_4557 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5144 = _T_5143 | _T_4889; // @[Mux.scala 27:72]
  wire  _T_4559 = btb_rd_addr_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4890 = _T_4559 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5145 = _T_5144 | _T_4890; // @[Mux.scala 27:72]
  wire  _T_4561 = btb_rd_addr_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4891 = _T_4561 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5146 = _T_5145 | _T_4891; // @[Mux.scala 27:72]
  wire  _T_4563 = btb_rd_addr_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4892 = _T_4563 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5147 = _T_5146 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4565 = btb_rd_addr_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4893 = _T_4565 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5148 = _T_5147 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4567 = btb_rd_addr_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4894 = _T_4567 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5149 = _T_5148 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4569 = btb_rd_addr_p1_f == 8'hba; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4895 = _T_4569 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5150 = _T_5149 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4571 = btb_rd_addr_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4896 = _T_4571 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5151 = _T_5150 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4573 = btb_rd_addr_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4897 = _T_4573 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5152 = _T_5151 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4575 = btb_rd_addr_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4898 = _T_4575 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5153 = _T_5152 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4577 = btb_rd_addr_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4899 = _T_4577 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5154 = _T_5153 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4579 = btb_rd_addr_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4900 = _T_4579 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5155 = _T_5154 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4581 = btb_rd_addr_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4901 = _T_4581 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5156 = _T_5155 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4583 = btb_rd_addr_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4902 = _T_4583 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5157 = _T_5156 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4585 = btb_rd_addr_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4903 = _T_4585 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5158 = _T_5157 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4587 = btb_rd_addr_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4904 = _T_4587 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5159 = _T_5158 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4589 = btb_rd_addr_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4905 = _T_4589 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5160 = _T_5159 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4591 = btb_rd_addr_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4906 = _T_4591 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5161 = _T_5160 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4593 = btb_rd_addr_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4907 = _T_4593 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5162 = _T_5161 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4595 = btb_rd_addr_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4908 = _T_4595 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5163 = _T_5162 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4597 = btb_rd_addr_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4909 = _T_4597 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5164 = _T_5163 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4599 = btb_rd_addr_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4910 = _T_4599 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5165 = _T_5164 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4601 = btb_rd_addr_p1_f == 8'hca; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4911 = _T_4601 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5166 = _T_5165 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4603 = btb_rd_addr_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4912 = _T_4603 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5167 = _T_5166 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4605 = btb_rd_addr_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4913 = _T_4605 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5168 = _T_5167 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4607 = btb_rd_addr_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4914 = _T_4607 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5169 = _T_5168 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4609 = btb_rd_addr_p1_f == 8'hce; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4915 = _T_4609 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5170 = _T_5169 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4611 = btb_rd_addr_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4916 = _T_4611 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5171 = _T_5170 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4613 = btb_rd_addr_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4917 = _T_4613 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5172 = _T_5171 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4615 = btb_rd_addr_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4918 = _T_4615 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5173 = _T_5172 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4617 = btb_rd_addr_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4919 = _T_4617 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5174 = _T_5173 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4619 = btb_rd_addr_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4920 = _T_4619 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5175 = _T_5174 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4621 = btb_rd_addr_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4921 = _T_4621 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5176 = _T_5175 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4623 = btb_rd_addr_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4922 = _T_4623 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5177 = _T_5176 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4625 = btb_rd_addr_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4923 = _T_4625 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5178 = _T_5177 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4627 = btb_rd_addr_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4924 = _T_4627 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5179 = _T_5178 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4629 = btb_rd_addr_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4925 = _T_4629 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5180 = _T_5179 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_4631 = btb_rd_addr_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4926 = _T_4631 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5181 = _T_5180 | _T_4926; // @[Mux.scala 27:72]
  wire  _T_4633 = btb_rd_addr_p1_f == 8'hda; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4927 = _T_4633 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5182 = _T_5181 | _T_4927; // @[Mux.scala 27:72]
  wire  _T_4635 = btb_rd_addr_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4928 = _T_4635 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5183 = _T_5182 | _T_4928; // @[Mux.scala 27:72]
  wire  _T_4637 = btb_rd_addr_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4929 = _T_4637 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5184 = _T_5183 | _T_4929; // @[Mux.scala 27:72]
  wire  _T_4639 = btb_rd_addr_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4930 = _T_4639 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5185 = _T_5184 | _T_4930; // @[Mux.scala 27:72]
  wire  _T_4641 = btb_rd_addr_p1_f == 8'hde; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4931 = _T_4641 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5186 = _T_5185 | _T_4931; // @[Mux.scala 27:72]
  wire  _T_4643 = btb_rd_addr_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4932 = _T_4643 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5187 = _T_5186 | _T_4932; // @[Mux.scala 27:72]
  wire  _T_4645 = btb_rd_addr_p1_f == 8'he0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4933 = _T_4645 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5188 = _T_5187 | _T_4933; // @[Mux.scala 27:72]
  wire  _T_4647 = btb_rd_addr_p1_f == 8'he1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4934 = _T_4647 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5189 = _T_5188 | _T_4934; // @[Mux.scala 27:72]
  wire  _T_4649 = btb_rd_addr_p1_f == 8'he2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4935 = _T_4649 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5190 = _T_5189 | _T_4935; // @[Mux.scala 27:72]
  wire  _T_4651 = btb_rd_addr_p1_f == 8'he3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4936 = _T_4651 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5191 = _T_5190 | _T_4936; // @[Mux.scala 27:72]
  wire  _T_4653 = btb_rd_addr_p1_f == 8'he4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4937 = _T_4653 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5192 = _T_5191 | _T_4937; // @[Mux.scala 27:72]
  wire  _T_4655 = btb_rd_addr_p1_f == 8'he5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4938 = _T_4655 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5193 = _T_5192 | _T_4938; // @[Mux.scala 27:72]
  wire  _T_4657 = btb_rd_addr_p1_f == 8'he6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4939 = _T_4657 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5194 = _T_5193 | _T_4939; // @[Mux.scala 27:72]
  wire  _T_4659 = btb_rd_addr_p1_f == 8'he7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4940 = _T_4659 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5195 = _T_5194 | _T_4940; // @[Mux.scala 27:72]
  wire  _T_4661 = btb_rd_addr_p1_f == 8'he8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4941 = _T_4661 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5196 = _T_5195 | _T_4941; // @[Mux.scala 27:72]
  wire  _T_4663 = btb_rd_addr_p1_f == 8'he9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4942 = _T_4663 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5197 = _T_5196 | _T_4942; // @[Mux.scala 27:72]
  wire  _T_4665 = btb_rd_addr_p1_f == 8'hea; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4943 = _T_4665 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5198 = _T_5197 | _T_4943; // @[Mux.scala 27:72]
  wire  _T_4667 = btb_rd_addr_p1_f == 8'heb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4944 = _T_4667 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5199 = _T_5198 | _T_4944; // @[Mux.scala 27:72]
  wire  _T_4669 = btb_rd_addr_p1_f == 8'hec; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4945 = _T_4669 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5200 = _T_5199 | _T_4945; // @[Mux.scala 27:72]
  wire  _T_4671 = btb_rd_addr_p1_f == 8'hed; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4946 = _T_4671 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5201 = _T_5200 | _T_4946; // @[Mux.scala 27:72]
  wire  _T_4673 = btb_rd_addr_p1_f == 8'hee; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4947 = _T_4673 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5202 = _T_5201 | _T_4947; // @[Mux.scala 27:72]
  wire  _T_4675 = btb_rd_addr_p1_f == 8'hef; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4948 = _T_4675 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5203 = _T_5202 | _T_4948; // @[Mux.scala 27:72]
  wire  _T_4677 = btb_rd_addr_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4949 = _T_4677 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5204 = _T_5203 | _T_4949; // @[Mux.scala 27:72]
  wire  _T_4679 = btb_rd_addr_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4950 = _T_4679 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5205 = _T_5204 | _T_4950; // @[Mux.scala 27:72]
  wire  _T_4681 = btb_rd_addr_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4951 = _T_4681 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5206 = _T_5205 | _T_4951; // @[Mux.scala 27:72]
  wire  _T_4683 = btb_rd_addr_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4952 = _T_4683 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5207 = _T_5206 | _T_4952; // @[Mux.scala 27:72]
  wire  _T_4685 = btb_rd_addr_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4953 = _T_4685 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5208 = _T_5207 | _T_4953; // @[Mux.scala 27:72]
  wire  _T_4687 = btb_rd_addr_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4954 = _T_4687 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5209 = _T_5208 | _T_4954; // @[Mux.scala 27:72]
  wire  _T_4689 = btb_rd_addr_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4955 = _T_4689 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5210 = _T_5209 | _T_4955; // @[Mux.scala 27:72]
  wire  _T_4691 = btb_rd_addr_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4956 = _T_4691 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5211 = _T_5210 | _T_4956; // @[Mux.scala 27:72]
  wire  _T_4693 = btb_rd_addr_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4957 = _T_4693 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5212 = _T_5211 | _T_4957; // @[Mux.scala 27:72]
  wire  _T_4695 = btb_rd_addr_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4958 = _T_4695 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5213 = _T_5212 | _T_4958; // @[Mux.scala 27:72]
  wire  _T_4697 = btb_rd_addr_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4959 = _T_4697 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5214 = _T_5213 | _T_4959; // @[Mux.scala 27:72]
  wire  _T_4699 = btb_rd_addr_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4960 = _T_4699 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5215 = _T_5214 | _T_4960; // @[Mux.scala 27:72]
  wire  _T_4701 = btb_rd_addr_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4961 = _T_4701 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5216 = _T_5215 | _T_4961; // @[Mux.scala 27:72]
  wire  _T_4703 = btb_rd_addr_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4962 = _T_4703 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5217 = _T_5216 | _T_4962; // @[Mux.scala 27:72]
  wire  _T_4705 = btb_rd_addr_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4963 = _T_4705 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5218 = _T_5217 | _T_4963; // @[Mux.scala 27:72]
  wire  _T_4707 = btb_rd_addr_p1_f == 8'hff; // @[ifu_bp_ctl.scala 441:86]
  wire [21:0] _T_4964 = _T_4707 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5219 = _T_5218 | _T_4964; // @[Mux.scala 27:72]
  wire [21:0] _T_5220 = _T_5219; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5219; // @[ifu_bp_ctl.scala 441:31]
  wire [4:0] _T_35 = _T_8[13:9] ^ _T_8[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_p1_f = _T_35 ^ _T_8[23:19]; // @[lib.scala 42:111]
  wire  _T_64 = _T_5220[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 152:107]
  wire  _T_65 = _T_5220[0] & _T_64; // @[ifu_bp_ctl.scala 152:61]
  wire  _T_20 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 126:75]
  wire  branch_error_collision_p1_f = dec_tlu_error_wb & _T_20; // @[ifu_bp_ctl.scala 126:54]
  wire  branch_error_bank_conflict_p1_f = branch_error_collision_p1_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 130:69]
  wire  _T_66 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & branch_error_bank_conflict_p1_f; // @[ifu_bp_ctl.scala 153:22]
  wire  _T_67 = ~_T_66; // @[ifu_bp_ctl.scala 153:5]
  wire  _T_68 = _T_65 & _T_67; // @[ifu_bp_ctl.scala 152:130]
  wire  _T_69 = _T_68 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 153:57]
  wire  tag_match_way0_p1_f = _T_69 & _T; // @[ifu_bp_ctl.scala 153:78]
  wire  _T_100 = _T_5220[3] ^ _T_5220[4]; // @[ifu_bp_ctl.scala 165:99]
  wire  _T_101 = tag_match_way0_p1_f & _T_100; // @[ifu_bp_ctl.scala 165:62]
  wire  _T_105 = ~_T_100; // @[ifu_bp_ctl.scala 166:27]
  wire  _T_106 = tag_match_way0_p1_f & _T_105; // @[ifu_bp_ctl.scala 166:25]
  wire [1:0] tag_match_way0_expanded_p1_f = {_T_101,_T_106}; // @[Cat.scala 29:58]
  wire [21:0] _T_136 = tag_match_way0_expanded_p1_f[0] ? _T_5220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5733 = _T_4197 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5734 = _T_4199 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5989 = _T_5733 | _T_5734; // @[Mux.scala 27:72]
  wire [21:0] _T_5735 = _T_4201 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5990 = _T_5989 | _T_5735; // @[Mux.scala 27:72]
  wire [21:0] _T_5736 = _T_4203 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5991 = _T_5990 | _T_5736; // @[Mux.scala 27:72]
  wire [21:0] _T_5737 = _T_4205 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5992 = _T_5991 | _T_5737; // @[Mux.scala 27:72]
  wire [21:0] _T_5738 = _T_4207 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5993 = _T_5992 | _T_5738; // @[Mux.scala 27:72]
  wire [21:0] _T_5739 = _T_4209 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5994 = _T_5993 | _T_5739; // @[Mux.scala 27:72]
  wire [21:0] _T_5740 = _T_4211 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5995 = _T_5994 | _T_5740; // @[Mux.scala 27:72]
  wire [21:0] _T_5741 = _T_4213 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5996 = _T_5995 | _T_5741; // @[Mux.scala 27:72]
  wire [21:0] _T_5742 = _T_4215 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5997 = _T_5996 | _T_5742; // @[Mux.scala 27:72]
  wire [21:0] _T_5743 = _T_4217 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5998 = _T_5997 | _T_5743; // @[Mux.scala 27:72]
  wire [21:0] _T_5744 = _T_4219 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5999 = _T_5998 | _T_5744; // @[Mux.scala 27:72]
  wire [21:0] _T_5745 = _T_4221 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6000 = _T_5999 | _T_5745; // @[Mux.scala 27:72]
  wire [21:0] _T_5746 = _T_4223 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6001 = _T_6000 | _T_5746; // @[Mux.scala 27:72]
  wire [21:0] _T_5747 = _T_4225 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6002 = _T_6001 | _T_5747; // @[Mux.scala 27:72]
  wire [21:0] _T_5748 = _T_4227 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6003 = _T_6002 | _T_5748; // @[Mux.scala 27:72]
  wire [21:0] _T_5749 = _T_4229 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6004 = _T_6003 | _T_5749; // @[Mux.scala 27:72]
  wire [21:0] _T_5750 = _T_4231 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6005 = _T_6004 | _T_5750; // @[Mux.scala 27:72]
  wire [21:0] _T_5751 = _T_4233 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6006 = _T_6005 | _T_5751; // @[Mux.scala 27:72]
  wire [21:0] _T_5752 = _T_4235 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6007 = _T_6006 | _T_5752; // @[Mux.scala 27:72]
  wire [21:0] _T_5753 = _T_4237 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6008 = _T_6007 | _T_5753; // @[Mux.scala 27:72]
  wire [21:0] _T_5754 = _T_4239 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6009 = _T_6008 | _T_5754; // @[Mux.scala 27:72]
  wire [21:0] _T_5755 = _T_4241 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6010 = _T_6009 | _T_5755; // @[Mux.scala 27:72]
  wire [21:0] _T_5756 = _T_4243 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6011 = _T_6010 | _T_5756; // @[Mux.scala 27:72]
  wire [21:0] _T_5757 = _T_4245 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6012 = _T_6011 | _T_5757; // @[Mux.scala 27:72]
  wire [21:0] _T_5758 = _T_4247 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6013 = _T_6012 | _T_5758; // @[Mux.scala 27:72]
  wire [21:0] _T_5759 = _T_4249 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6014 = _T_6013 | _T_5759; // @[Mux.scala 27:72]
  wire [21:0] _T_5760 = _T_4251 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6015 = _T_6014 | _T_5760; // @[Mux.scala 27:72]
  wire [21:0] _T_5761 = _T_4253 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6016 = _T_6015 | _T_5761; // @[Mux.scala 27:72]
  wire [21:0] _T_5762 = _T_4255 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6017 = _T_6016 | _T_5762; // @[Mux.scala 27:72]
  wire [21:0] _T_5763 = _T_4257 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6018 = _T_6017 | _T_5763; // @[Mux.scala 27:72]
  wire [21:0] _T_5764 = _T_4259 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6019 = _T_6018 | _T_5764; // @[Mux.scala 27:72]
  wire [21:0] _T_5765 = _T_4261 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6020 = _T_6019 | _T_5765; // @[Mux.scala 27:72]
  wire [21:0] _T_5766 = _T_4263 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6021 = _T_6020 | _T_5766; // @[Mux.scala 27:72]
  wire [21:0] _T_5767 = _T_4265 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6022 = _T_6021 | _T_5767; // @[Mux.scala 27:72]
  wire [21:0] _T_5768 = _T_4267 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6023 = _T_6022 | _T_5768; // @[Mux.scala 27:72]
  wire [21:0] _T_5769 = _T_4269 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6024 = _T_6023 | _T_5769; // @[Mux.scala 27:72]
  wire [21:0] _T_5770 = _T_4271 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6025 = _T_6024 | _T_5770; // @[Mux.scala 27:72]
  wire [21:0] _T_5771 = _T_4273 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6026 = _T_6025 | _T_5771; // @[Mux.scala 27:72]
  wire [21:0] _T_5772 = _T_4275 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6027 = _T_6026 | _T_5772; // @[Mux.scala 27:72]
  wire [21:0] _T_5773 = _T_4277 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6028 = _T_6027 | _T_5773; // @[Mux.scala 27:72]
  wire [21:0] _T_5774 = _T_4279 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6029 = _T_6028 | _T_5774; // @[Mux.scala 27:72]
  wire [21:0] _T_5775 = _T_4281 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6030 = _T_6029 | _T_5775; // @[Mux.scala 27:72]
  wire [21:0] _T_5776 = _T_4283 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6031 = _T_6030 | _T_5776; // @[Mux.scala 27:72]
  wire [21:0] _T_5777 = _T_4285 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6032 = _T_6031 | _T_5777; // @[Mux.scala 27:72]
  wire [21:0] _T_5778 = _T_4287 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6033 = _T_6032 | _T_5778; // @[Mux.scala 27:72]
  wire [21:0] _T_5779 = _T_4289 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6034 = _T_6033 | _T_5779; // @[Mux.scala 27:72]
  wire [21:0] _T_5780 = _T_4291 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6035 = _T_6034 | _T_5780; // @[Mux.scala 27:72]
  wire [21:0] _T_5781 = _T_4293 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6036 = _T_6035 | _T_5781; // @[Mux.scala 27:72]
  wire [21:0] _T_5782 = _T_4295 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6037 = _T_6036 | _T_5782; // @[Mux.scala 27:72]
  wire [21:0] _T_5783 = _T_4297 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6038 = _T_6037 | _T_5783; // @[Mux.scala 27:72]
  wire [21:0] _T_5784 = _T_4299 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6039 = _T_6038 | _T_5784; // @[Mux.scala 27:72]
  wire [21:0] _T_5785 = _T_4301 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6040 = _T_6039 | _T_5785; // @[Mux.scala 27:72]
  wire [21:0] _T_5786 = _T_4303 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6041 = _T_6040 | _T_5786; // @[Mux.scala 27:72]
  wire [21:0] _T_5787 = _T_4305 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6042 = _T_6041 | _T_5787; // @[Mux.scala 27:72]
  wire [21:0] _T_5788 = _T_4307 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6043 = _T_6042 | _T_5788; // @[Mux.scala 27:72]
  wire [21:0] _T_5789 = _T_4309 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6044 = _T_6043 | _T_5789; // @[Mux.scala 27:72]
  wire [21:0] _T_5790 = _T_4311 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6045 = _T_6044 | _T_5790; // @[Mux.scala 27:72]
  wire [21:0] _T_5791 = _T_4313 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6046 = _T_6045 | _T_5791; // @[Mux.scala 27:72]
  wire [21:0] _T_5792 = _T_4315 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6047 = _T_6046 | _T_5792; // @[Mux.scala 27:72]
  wire [21:0] _T_5793 = _T_4317 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6048 = _T_6047 | _T_5793; // @[Mux.scala 27:72]
  wire [21:0] _T_5794 = _T_4319 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6049 = _T_6048 | _T_5794; // @[Mux.scala 27:72]
  wire [21:0] _T_5795 = _T_4321 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6050 = _T_6049 | _T_5795; // @[Mux.scala 27:72]
  wire [21:0] _T_5796 = _T_4323 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6051 = _T_6050 | _T_5796; // @[Mux.scala 27:72]
  wire [21:0] _T_5797 = _T_4325 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6052 = _T_6051 | _T_5797; // @[Mux.scala 27:72]
  wire [21:0] _T_5798 = _T_4327 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6053 = _T_6052 | _T_5798; // @[Mux.scala 27:72]
  wire [21:0] _T_5799 = _T_4329 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6054 = _T_6053 | _T_5799; // @[Mux.scala 27:72]
  wire [21:0] _T_5800 = _T_4331 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6055 = _T_6054 | _T_5800; // @[Mux.scala 27:72]
  wire [21:0] _T_5801 = _T_4333 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6056 = _T_6055 | _T_5801; // @[Mux.scala 27:72]
  wire [21:0] _T_5802 = _T_4335 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6057 = _T_6056 | _T_5802; // @[Mux.scala 27:72]
  wire [21:0] _T_5803 = _T_4337 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6058 = _T_6057 | _T_5803; // @[Mux.scala 27:72]
  wire [21:0] _T_5804 = _T_4339 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6059 = _T_6058 | _T_5804; // @[Mux.scala 27:72]
  wire [21:0] _T_5805 = _T_4341 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6060 = _T_6059 | _T_5805; // @[Mux.scala 27:72]
  wire [21:0] _T_5806 = _T_4343 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6061 = _T_6060 | _T_5806; // @[Mux.scala 27:72]
  wire [21:0] _T_5807 = _T_4345 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6062 = _T_6061 | _T_5807; // @[Mux.scala 27:72]
  wire [21:0] _T_5808 = _T_4347 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6063 = _T_6062 | _T_5808; // @[Mux.scala 27:72]
  wire [21:0] _T_5809 = _T_4349 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6064 = _T_6063 | _T_5809; // @[Mux.scala 27:72]
  wire [21:0] _T_5810 = _T_4351 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6065 = _T_6064 | _T_5810; // @[Mux.scala 27:72]
  wire [21:0] _T_5811 = _T_4353 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6066 = _T_6065 | _T_5811; // @[Mux.scala 27:72]
  wire [21:0] _T_5812 = _T_4355 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6067 = _T_6066 | _T_5812; // @[Mux.scala 27:72]
  wire [21:0] _T_5813 = _T_4357 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6068 = _T_6067 | _T_5813; // @[Mux.scala 27:72]
  wire [21:0] _T_5814 = _T_4359 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6069 = _T_6068 | _T_5814; // @[Mux.scala 27:72]
  wire [21:0] _T_5815 = _T_4361 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6070 = _T_6069 | _T_5815; // @[Mux.scala 27:72]
  wire [21:0] _T_5816 = _T_4363 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6071 = _T_6070 | _T_5816; // @[Mux.scala 27:72]
  wire [21:0] _T_5817 = _T_4365 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6072 = _T_6071 | _T_5817; // @[Mux.scala 27:72]
  wire [21:0] _T_5818 = _T_4367 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6073 = _T_6072 | _T_5818; // @[Mux.scala 27:72]
  wire [21:0] _T_5819 = _T_4369 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6074 = _T_6073 | _T_5819; // @[Mux.scala 27:72]
  wire [21:0] _T_5820 = _T_4371 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6075 = _T_6074 | _T_5820; // @[Mux.scala 27:72]
  wire [21:0] _T_5821 = _T_4373 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6076 = _T_6075 | _T_5821; // @[Mux.scala 27:72]
  wire [21:0] _T_5822 = _T_4375 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6077 = _T_6076 | _T_5822; // @[Mux.scala 27:72]
  wire [21:0] _T_5823 = _T_4377 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6078 = _T_6077 | _T_5823; // @[Mux.scala 27:72]
  wire [21:0] _T_5824 = _T_4379 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6079 = _T_6078 | _T_5824; // @[Mux.scala 27:72]
  wire [21:0] _T_5825 = _T_4381 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6080 = _T_6079 | _T_5825; // @[Mux.scala 27:72]
  wire [21:0] _T_5826 = _T_4383 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6081 = _T_6080 | _T_5826; // @[Mux.scala 27:72]
  wire [21:0] _T_5827 = _T_4385 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6082 = _T_6081 | _T_5827; // @[Mux.scala 27:72]
  wire [21:0] _T_5828 = _T_4387 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6083 = _T_6082 | _T_5828; // @[Mux.scala 27:72]
  wire [21:0] _T_5829 = _T_4389 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6084 = _T_6083 | _T_5829; // @[Mux.scala 27:72]
  wire [21:0] _T_5830 = _T_4391 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6085 = _T_6084 | _T_5830; // @[Mux.scala 27:72]
  wire [21:0] _T_5831 = _T_4393 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6086 = _T_6085 | _T_5831; // @[Mux.scala 27:72]
  wire [21:0] _T_5832 = _T_4395 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6087 = _T_6086 | _T_5832; // @[Mux.scala 27:72]
  wire [21:0] _T_5833 = _T_4397 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6088 = _T_6087 | _T_5833; // @[Mux.scala 27:72]
  wire [21:0] _T_5834 = _T_4399 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6089 = _T_6088 | _T_5834; // @[Mux.scala 27:72]
  wire [21:0] _T_5835 = _T_4401 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6090 = _T_6089 | _T_5835; // @[Mux.scala 27:72]
  wire [21:0] _T_5836 = _T_4403 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6091 = _T_6090 | _T_5836; // @[Mux.scala 27:72]
  wire [21:0] _T_5837 = _T_4405 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6092 = _T_6091 | _T_5837; // @[Mux.scala 27:72]
  wire [21:0] _T_5838 = _T_4407 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6093 = _T_6092 | _T_5838; // @[Mux.scala 27:72]
  wire [21:0] _T_5839 = _T_4409 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6094 = _T_6093 | _T_5839; // @[Mux.scala 27:72]
  wire [21:0] _T_5840 = _T_4411 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6095 = _T_6094 | _T_5840; // @[Mux.scala 27:72]
  wire [21:0] _T_5841 = _T_4413 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6096 = _T_6095 | _T_5841; // @[Mux.scala 27:72]
  wire [21:0] _T_5842 = _T_4415 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6097 = _T_6096 | _T_5842; // @[Mux.scala 27:72]
  wire [21:0] _T_5843 = _T_4417 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6098 = _T_6097 | _T_5843; // @[Mux.scala 27:72]
  wire [21:0] _T_5844 = _T_4419 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6099 = _T_6098 | _T_5844; // @[Mux.scala 27:72]
  wire [21:0] _T_5845 = _T_4421 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6100 = _T_6099 | _T_5845; // @[Mux.scala 27:72]
  wire [21:0] _T_5846 = _T_4423 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6101 = _T_6100 | _T_5846; // @[Mux.scala 27:72]
  wire [21:0] _T_5847 = _T_4425 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6102 = _T_6101 | _T_5847; // @[Mux.scala 27:72]
  wire [21:0] _T_5848 = _T_4427 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6103 = _T_6102 | _T_5848; // @[Mux.scala 27:72]
  wire [21:0] _T_5849 = _T_4429 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6104 = _T_6103 | _T_5849; // @[Mux.scala 27:72]
  wire [21:0] _T_5850 = _T_4431 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6105 = _T_6104 | _T_5850; // @[Mux.scala 27:72]
  wire [21:0] _T_5851 = _T_4433 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6106 = _T_6105 | _T_5851; // @[Mux.scala 27:72]
  wire [21:0] _T_5852 = _T_4435 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6107 = _T_6106 | _T_5852; // @[Mux.scala 27:72]
  wire [21:0] _T_5853 = _T_4437 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6108 = _T_6107 | _T_5853; // @[Mux.scala 27:72]
  wire [21:0] _T_5854 = _T_4439 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6109 = _T_6108 | _T_5854; // @[Mux.scala 27:72]
  wire [21:0] _T_5855 = _T_4441 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6110 = _T_6109 | _T_5855; // @[Mux.scala 27:72]
  wire [21:0] _T_5856 = _T_4443 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6111 = _T_6110 | _T_5856; // @[Mux.scala 27:72]
  wire [21:0] _T_5857 = _T_4445 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6112 = _T_6111 | _T_5857; // @[Mux.scala 27:72]
  wire [21:0] _T_5858 = _T_4447 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6113 = _T_6112 | _T_5858; // @[Mux.scala 27:72]
  wire [21:0] _T_5859 = _T_4449 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6114 = _T_6113 | _T_5859; // @[Mux.scala 27:72]
  wire [21:0] _T_5860 = _T_4451 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6115 = _T_6114 | _T_5860; // @[Mux.scala 27:72]
  wire [21:0] _T_5861 = _T_4453 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6116 = _T_6115 | _T_5861; // @[Mux.scala 27:72]
  wire [21:0] _T_5862 = _T_4455 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6117 = _T_6116 | _T_5862; // @[Mux.scala 27:72]
  wire [21:0] _T_5863 = _T_4457 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6118 = _T_6117 | _T_5863; // @[Mux.scala 27:72]
  wire [21:0] _T_5864 = _T_4459 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6119 = _T_6118 | _T_5864; // @[Mux.scala 27:72]
  wire [21:0] _T_5865 = _T_4461 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6120 = _T_6119 | _T_5865; // @[Mux.scala 27:72]
  wire [21:0] _T_5866 = _T_4463 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6121 = _T_6120 | _T_5866; // @[Mux.scala 27:72]
  wire [21:0] _T_5867 = _T_4465 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6122 = _T_6121 | _T_5867; // @[Mux.scala 27:72]
  wire [21:0] _T_5868 = _T_4467 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6123 = _T_6122 | _T_5868; // @[Mux.scala 27:72]
  wire [21:0] _T_5869 = _T_4469 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6124 = _T_6123 | _T_5869; // @[Mux.scala 27:72]
  wire [21:0] _T_5870 = _T_4471 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6125 = _T_6124 | _T_5870; // @[Mux.scala 27:72]
  wire [21:0] _T_5871 = _T_4473 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6126 = _T_6125 | _T_5871; // @[Mux.scala 27:72]
  wire [21:0] _T_5872 = _T_4475 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6127 = _T_6126 | _T_5872; // @[Mux.scala 27:72]
  wire [21:0] _T_5873 = _T_4477 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6128 = _T_6127 | _T_5873; // @[Mux.scala 27:72]
  wire [21:0] _T_5874 = _T_4479 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6129 = _T_6128 | _T_5874; // @[Mux.scala 27:72]
  wire [21:0] _T_5875 = _T_4481 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6130 = _T_6129 | _T_5875; // @[Mux.scala 27:72]
  wire [21:0] _T_5876 = _T_4483 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6131 = _T_6130 | _T_5876; // @[Mux.scala 27:72]
  wire [21:0] _T_5877 = _T_4485 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6132 = _T_6131 | _T_5877; // @[Mux.scala 27:72]
  wire [21:0] _T_5878 = _T_4487 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6133 = _T_6132 | _T_5878; // @[Mux.scala 27:72]
  wire [21:0] _T_5879 = _T_4489 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6134 = _T_6133 | _T_5879; // @[Mux.scala 27:72]
  wire [21:0] _T_5880 = _T_4491 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6135 = _T_6134 | _T_5880; // @[Mux.scala 27:72]
  wire [21:0] _T_5881 = _T_4493 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6136 = _T_6135 | _T_5881; // @[Mux.scala 27:72]
  wire [21:0] _T_5882 = _T_4495 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6137 = _T_6136 | _T_5882; // @[Mux.scala 27:72]
  wire [21:0] _T_5883 = _T_4497 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6138 = _T_6137 | _T_5883; // @[Mux.scala 27:72]
  wire [21:0] _T_5884 = _T_4499 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6139 = _T_6138 | _T_5884; // @[Mux.scala 27:72]
  wire [21:0] _T_5885 = _T_4501 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6140 = _T_6139 | _T_5885; // @[Mux.scala 27:72]
  wire [21:0] _T_5886 = _T_4503 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6141 = _T_6140 | _T_5886; // @[Mux.scala 27:72]
  wire [21:0] _T_5887 = _T_4505 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6142 = _T_6141 | _T_5887; // @[Mux.scala 27:72]
  wire [21:0] _T_5888 = _T_4507 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6143 = _T_6142 | _T_5888; // @[Mux.scala 27:72]
  wire [21:0] _T_5889 = _T_4509 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6144 = _T_6143 | _T_5889; // @[Mux.scala 27:72]
  wire [21:0] _T_5890 = _T_4511 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6145 = _T_6144 | _T_5890; // @[Mux.scala 27:72]
  wire [21:0] _T_5891 = _T_4513 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6146 = _T_6145 | _T_5891; // @[Mux.scala 27:72]
  wire [21:0] _T_5892 = _T_4515 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6147 = _T_6146 | _T_5892; // @[Mux.scala 27:72]
  wire [21:0] _T_5893 = _T_4517 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6148 = _T_6147 | _T_5893; // @[Mux.scala 27:72]
  wire [21:0] _T_5894 = _T_4519 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6149 = _T_6148 | _T_5894; // @[Mux.scala 27:72]
  wire [21:0] _T_5895 = _T_4521 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6150 = _T_6149 | _T_5895; // @[Mux.scala 27:72]
  wire [21:0] _T_5896 = _T_4523 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6151 = _T_6150 | _T_5896; // @[Mux.scala 27:72]
  wire [21:0] _T_5897 = _T_4525 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6152 = _T_6151 | _T_5897; // @[Mux.scala 27:72]
  wire [21:0] _T_5898 = _T_4527 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6153 = _T_6152 | _T_5898; // @[Mux.scala 27:72]
  wire [21:0] _T_5899 = _T_4529 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6154 = _T_6153 | _T_5899; // @[Mux.scala 27:72]
  wire [21:0] _T_5900 = _T_4531 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6155 = _T_6154 | _T_5900; // @[Mux.scala 27:72]
  wire [21:0] _T_5901 = _T_4533 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6156 = _T_6155 | _T_5901; // @[Mux.scala 27:72]
  wire [21:0] _T_5902 = _T_4535 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6157 = _T_6156 | _T_5902; // @[Mux.scala 27:72]
  wire [21:0] _T_5903 = _T_4537 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6158 = _T_6157 | _T_5903; // @[Mux.scala 27:72]
  wire [21:0] _T_5904 = _T_4539 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6159 = _T_6158 | _T_5904; // @[Mux.scala 27:72]
  wire [21:0] _T_5905 = _T_4541 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6160 = _T_6159 | _T_5905; // @[Mux.scala 27:72]
  wire [21:0] _T_5906 = _T_4543 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6161 = _T_6160 | _T_5906; // @[Mux.scala 27:72]
  wire [21:0] _T_5907 = _T_4545 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6162 = _T_6161 | _T_5907; // @[Mux.scala 27:72]
  wire [21:0] _T_5908 = _T_4547 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6163 = _T_6162 | _T_5908; // @[Mux.scala 27:72]
  wire [21:0] _T_5909 = _T_4549 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6164 = _T_6163 | _T_5909; // @[Mux.scala 27:72]
  wire [21:0] _T_5910 = _T_4551 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6165 = _T_6164 | _T_5910; // @[Mux.scala 27:72]
  wire [21:0] _T_5911 = _T_4553 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6166 = _T_6165 | _T_5911; // @[Mux.scala 27:72]
  wire [21:0] _T_5912 = _T_4555 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6167 = _T_6166 | _T_5912; // @[Mux.scala 27:72]
  wire [21:0] _T_5913 = _T_4557 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6168 = _T_6167 | _T_5913; // @[Mux.scala 27:72]
  wire [21:0] _T_5914 = _T_4559 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6169 = _T_6168 | _T_5914; // @[Mux.scala 27:72]
  wire [21:0] _T_5915 = _T_4561 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6170 = _T_6169 | _T_5915; // @[Mux.scala 27:72]
  wire [21:0] _T_5916 = _T_4563 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6171 = _T_6170 | _T_5916; // @[Mux.scala 27:72]
  wire [21:0] _T_5917 = _T_4565 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6172 = _T_6171 | _T_5917; // @[Mux.scala 27:72]
  wire [21:0] _T_5918 = _T_4567 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6173 = _T_6172 | _T_5918; // @[Mux.scala 27:72]
  wire [21:0] _T_5919 = _T_4569 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6174 = _T_6173 | _T_5919; // @[Mux.scala 27:72]
  wire [21:0] _T_5920 = _T_4571 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6175 = _T_6174 | _T_5920; // @[Mux.scala 27:72]
  wire [21:0] _T_5921 = _T_4573 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6176 = _T_6175 | _T_5921; // @[Mux.scala 27:72]
  wire [21:0] _T_5922 = _T_4575 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6177 = _T_6176 | _T_5922; // @[Mux.scala 27:72]
  wire [21:0] _T_5923 = _T_4577 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6178 = _T_6177 | _T_5923; // @[Mux.scala 27:72]
  wire [21:0] _T_5924 = _T_4579 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6179 = _T_6178 | _T_5924; // @[Mux.scala 27:72]
  wire [21:0] _T_5925 = _T_4581 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6180 = _T_6179 | _T_5925; // @[Mux.scala 27:72]
  wire [21:0] _T_5926 = _T_4583 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6181 = _T_6180 | _T_5926; // @[Mux.scala 27:72]
  wire [21:0] _T_5927 = _T_4585 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6182 = _T_6181 | _T_5927; // @[Mux.scala 27:72]
  wire [21:0] _T_5928 = _T_4587 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6183 = _T_6182 | _T_5928; // @[Mux.scala 27:72]
  wire [21:0] _T_5929 = _T_4589 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6184 = _T_6183 | _T_5929; // @[Mux.scala 27:72]
  wire [21:0] _T_5930 = _T_4591 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6185 = _T_6184 | _T_5930; // @[Mux.scala 27:72]
  wire [21:0] _T_5931 = _T_4593 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6186 = _T_6185 | _T_5931; // @[Mux.scala 27:72]
  wire [21:0] _T_5932 = _T_4595 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6187 = _T_6186 | _T_5932; // @[Mux.scala 27:72]
  wire [21:0] _T_5933 = _T_4597 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6188 = _T_6187 | _T_5933; // @[Mux.scala 27:72]
  wire [21:0] _T_5934 = _T_4599 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6189 = _T_6188 | _T_5934; // @[Mux.scala 27:72]
  wire [21:0] _T_5935 = _T_4601 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6190 = _T_6189 | _T_5935; // @[Mux.scala 27:72]
  wire [21:0] _T_5936 = _T_4603 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6191 = _T_6190 | _T_5936; // @[Mux.scala 27:72]
  wire [21:0] _T_5937 = _T_4605 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6192 = _T_6191 | _T_5937; // @[Mux.scala 27:72]
  wire [21:0] _T_5938 = _T_4607 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6193 = _T_6192 | _T_5938; // @[Mux.scala 27:72]
  wire [21:0] _T_5939 = _T_4609 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6194 = _T_6193 | _T_5939; // @[Mux.scala 27:72]
  wire [21:0] _T_5940 = _T_4611 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6195 = _T_6194 | _T_5940; // @[Mux.scala 27:72]
  wire [21:0] _T_5941 = _T_4613 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6196 = _T_6195 | _T_5941; // @[Mux.scala 27:72]
  wire [21:0] _T_5942 = _T_4615 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6197 = _T_6196 | _T_5942; // @[Mux.scala 27:72]
  wire [21:0] _T_5943 = _T_4617 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6198 = _T_6197 | _T_5943; // @[Mux.scala 27:72]
  wire [21:0] _T_5944 = _T_4619 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6199 = _T_6198 | _T_5944; // @[Mux.scala 27:72]
  wire [21:0] _T_5945 = _T_4621 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6200 = _T_6199 | _T_5945; // @[Mux.scala 27:72]
  wire [21:0] _T_5946 = _T_4623 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6201 = _T_6200 | _T_5946; // @[Mux.scala 27:72]
  wire [21:0] _T_5947 = _T_4625 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6202 = _T_6201 | _T_5947; // @[Mux.scala 27:72]
  wire [21:0] _T_5948 = _T_4627 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6203 = _T_6202 | _T_5948; // @[Mux.scala 27:72]
  wire [21:0] _T_5949 = _T_4629 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6204 = _T_6203 | _T_5949; // @[Mux.scala 27:72]
  wire [21:0] _T_5950 = _T_4631 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6205 = _T_6204 | _T_5950; // @[Mux.scala 27:72]
  wire [21:0] _T_5951 = _T_4633 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6206 = _T_6205 | _T_5951; // @[Mux.scala 27:72]
  wire [21:0] _T_5952 = _T_4635 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6207 = _T_6206 | _T_5952; // @[Mux.scala 27:72]
  wire [21:0] _T_5953 = _T_4637 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6208 = _T_6207 | _T_5953; // @[Mux.scala 27:72]
  wire [21:0] _T_5954 = _T_4639 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6209 = _T_6208 | _T_5954; // @[Mux.scala 27:72]
  wire [21:0] _T_5955 = _T_4641 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6210 = _T_6209 | _T_5955; // @[Mux.scala 27:72]
  wire [21:0] _T_5956 = _T_4643 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6211 = _T_6210 | _T_5956; // @[Mux.scala 27:72]
  wire [21:0] _T_5957 = _T_4645 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6212 = _T_6211 | _T_5957; // @[Mux.scala 27:72]
  wire [21:0] _T_5958 = _T_4647 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6213 = _T_6212 | _T_5958; // @[Mux.scala 27:72]
  wire [21:0] _T_5959 = _T_4649 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6214 = _T_6213 | _T_5959; // @[Mux.scala 27:72]
  wire [21:0] _T_5960 = _T_4651 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6215 = _T_6214 | _T_5960; // @[Mux.scala 27:72]
  wire [21:0] _T_5961 = _T_4653 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6216 = _T_6215 | _T_5961; // @[Mux.scala 27:72]
  wire [21:0] _T_5962 = _T_4655 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6217 = _T_6216 | _T_5962; // @[Mux.scala 27:72]
  wire [21:0] _T_5963 = _T_4657 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6218 = _T_6217 | _T_5963; // @[Mux.scala 27:72]
  wire [21:0] _T_5964 = _T_4659 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6219 = _T_6218 | _T_5964; // @[Mux.scala 27:72]
  wire [21:0] _T_5965 = _T_4661 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6220 = _T_6219 | _T_5965; // @[Mux.scala 27:72]
  wire [21:0] _T_5966 = _T_4663 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6221 = _T_6220 | _T_5966; // @[Mux.scala 27:72]
  wire [21:0] _T_5967 = _T_4665 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6222 = _T_6221 | _T_5967; // @[Mux.scala 27:72]
  wire [21:0] _T_5968 = _T_4667 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6223 = _T_6222 | _T_5968; // @[Mux.scala 27:72]
  wire [21:0] _T_5969 = _T_4669 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6224 = _T_6223 | _T_5969; // @[Mux.scala 27:72]
  wire [21:0] _T_5970 = _T_4671 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6225 = _T_6224 | _T_5970; // @[Mux.scala 27:72]
  wire [21:0] _T_5971 = _T_4673 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6226 = _T_6225 | _T_5971; // @[Mux.scala 27:72]
  wire [21:0] _T_5972 = _T_4675 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6227 = _T_6226 | _T_5972; // @[Mux.scala 27:72]
  wire [21:0] _T_5973 = _T_4677 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6228 = _T_6227 | _T_5973; // @[Mux.scala 27:72]
  wire [21:0] _T_5974 = _T_4679 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6229 = _T_6228 | _T_5974; // @[Mux.scala 27:72]
  wire [21:0] _T_5975 = _T_4681 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6230 = _T_6229 | _T_5975; // @[Mux.scala 27:72]
  wire [21:0] _T_5976 = _T_4683 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6231 = _T_6230 | _T_5976; // @[Mux.scala 27:72]
  wire [21:0] _T_5977 = _T_4685 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6232 = _T_6231 | _T_5977; // @[Mux.scala 27:72]
  wire [21:0] _T_5978 = _T_4687 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6233 = _T_6232 | _T_5978; // @[Mux.scala 27:72]
  wire [21:0] _T_5979 = _T_4689 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6234 = _T_6233 | _T_5979; // @[Mux.scala 27:72]
  wire [21:0] _T_5980 = _T_4691 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6235 = _T_6234 | _T_5980; // @[Mux.scala 27:72]
  wire [21:0] _T_5981 = _T_4693 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6236 = _T_6235 | _T_5981; // @[Mux.scala 27:72]
  wire [21:0] _T_5982 = _T_4695 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6237 = _T_6236 | _T_5982; // @[Mux.scala 27:72]
  wire [21:0] _T_5983 = _T_4697 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6238 = _T_6237 | _T_5983; // @[Mux.scala 27:72]
  wire [21:0] _T_5984 = _T_4699 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6239 = _T_6238 | _T_5984; // @[Mux.scala 27:72]
  wire [21:0] _T_5985 = _T_4701 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6240 = _T_6239 | _T_5985; // @[Mux.scala 27:72]
  wire [21:0] _T_5986 = _T_4703 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6241 = _T_6240 | _T_5986; // @[Mux.scala 27:72]
  wire [21:0] _T_5987 = _T_4705 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6242 = _T_6241 | _T_5987; // @[Mux.scala 27:72]
  wire [21:0] _T_5988 = _T_4707 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6243 = _T_6242 | _T_5988; // @[Mux.scala 27:72]
  wire [21:0] _T_6244 = _T_6243; // @[Mux.scala 27:72 Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6243; // @[ifu_bp_ctl.scala 444:31]
  wire  _T_73 = _T_6244[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 155:107]
  wire  _T_74 = _T_6244[0] & _T_73; // @[ifu_bp_ctl.scala 155:61]
  wire  _T_77 = _T_74 & _T_67; // @[ifu_bp_ctl.scala 155:130]
  wire  _T_78 = _T_77 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 156:57]
  wire  tag_match_way1_p1_f = _T_78 & _T; // @[ifu_bp_ctl.scala 156:78]
  wire  _T_109 = _T_6244[3] ^ _T_6244[4]; // @[ifu_bp_ctl.scala 168:99]
  wire  _T_110 = tag_match_way1_p1_f & _T_109; // @[ifu_bp_ctl.scala 168:62]
  wire  _T_114 = ~_T_109; // @[ifu_bp_ctl.scala 169:27]
  wire  _T_115 = tag_match_way1_p1_f & _T_114; // @[ifu_bp_ctl.scala 169:25]
  wire [1:0] tag_match_way1_expanded_p1_f = {_T_110,_T_115}; // @[Cat.scala 29:58]
  wire [21:0] _T_137 = tag_match_way1_expanded_p1_f[0] ? _T_6244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_p1_f = _T_136 | _T_137; // @[Mux.scala 27:72]
  wire [21:0] _T_150 = io_ifc_fetch_addr_f[0] ? btb_bank0e_rd_data_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_149 | _T_150; // @[Mux.scala 27:72]
  wire  _T_236 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 280:59]
  wire [21:0] _T_122 = tag_match_way0_expanded_f[0] ? _T_3172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_123 = tag_match_way1_expanded_f[0] ? _T_4196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_f = _T_122 | _T_123; // @[Mux.scala 27:72]
  wire [21:0] _T_142 = _T_147 ? btb_bank0e_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_143 = io_ifc_fetch_addr_f[0] ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_142 | _T_143; // @[Mux.scala 27:72]
  wire  _T_239 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 281:59]
  wire [1:0] bht_force_taken_f = {_T_236,_T_239}; // @[Cat.scala 29:58]
  wire [9:0] _T_582 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[Reg.scala 27:20]
  wire [7:0] bht_rd_addr_hashed_f = _T_582[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_21957 = bht_rd_addr_hashed_f == 8'h0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_22469 = _T_21957 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_21959 = bht_rd_addr_hashed_f == 8'h1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_22470 = _T_21959 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22725 = _T_22469 | _T_22470; // @[Mux.scala 27:72]
  wire  _T_21961 = bht_rd_addr_hashed_f == 8'h2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_22471 = _T_21961 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22726 = _T_22725 | _T_22471; // @[Mux.scala 27:72]
  wire  _T_21963 = bht_rd_addr_hashed_f == 8'h3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_22472 = _T_21963 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22727 = _T_22726 | _T_22472; // @[Mux.scala 27:72]
  wire  _T_21965 = bht_rd_addr_hashed_f == 8'h4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_22473 = _T_21965 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22728 = _T_22727 | _T_22473; // @[Mux.scala 27:72]
  wire  _T_21967 = bht_rd_addr_hashed_f == 8'h5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_22474 = _T_21967 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22729 = _T_22728 | _T_22474; // @[Mux.scala 27:72]
  wire  _T_21969 = bht_rd_addr_hashed_f == 8'h6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_22475 = _T_21969 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22730 = _T_22729 | _T_22475; // @[Mux.scala 27:72]
  wire  _T_21971 = bht_rd_addr_hashed_f == 8'h7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_22476 = _T_21971 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22731 = _T_22730 | _T_22476; // @[Mux.scala 27:72]
  wire  _T_21973 = bht_rd_addr_hashed_f == 8'h8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_22477 = _T_21973 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22732 = _T_22731 | _T_22477; // @[Mux.scala 27:72]
  wire  _T_21975 = bht_rd_addr_hashed_f == 8'h9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_22478 = _T_21975 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22733 = _T_22732 | _T_22478; // @[Mux.scala 27:72]
  wire  _T_21977 = bht_rd_addr_hashed_f == 8'ha; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_22479 = _T_21977 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22734 = _T_22733 | _T_22479; // @[Mux.scala 27:72]
  wire  _T_21979 = bht_rd_addr_hashed_f == 8'hb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_22480 = _T_21979 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22735 = _T_22734 | _T_22480; // @[Mux.scala 27:72]
  wire  _T_21981 = bht_rd_addr_hashed_f == 8'hc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_22481 = _T_21981 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22736 = _T_22735 | _T_22481; // @[Mux.scala 27:72]
  wire  _T_21983 = bht_rd_addr_hashed_f == 8'hd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_22482 = _T_21983 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22737 = _T_22736 | _T_22482; // @[Mux.scala 27:72]
  wire  _T_21985 = bht_rd_addr_hashed_f == 8'he; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_22483 = _T_21985 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22738 = _T_22737 | _T_22483; // @[Mux.scala 27:72]
  wire  _T_21987 = bht_rd_addr_hashed_f == 8'hf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_22484 = _T_21987 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22739 = _T_22738 | _T_22484; // @[Mux.scala 27:72]
  wire  _T_21989 = bht_rd_addr_hashed_f == 8'h10; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_22485 = _T_21989 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22740 = _T_22739 | _T_22485; // @[Mux.scala 27:72]
  wire  _T_21991 = bht_rd_addr_hashed_f == 8'h11; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_22486 = _T_21991 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22741 = _T_22740 | _T_22486; // @[Mux.scala 27:72]
  wire  _T_21993 = bht_rd_addr_hashed_f == 8'h12; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_22487 = _T_21993 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22742 = _T_22741 | _T_22487; // @[Mux.scala 27:72]
  wire  _T_21995 = bht_rd_addr_hashed_f == 8'h13; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_22488 = _T_21995 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22743 = _T_22742 | _T_22488; // @[Mux.scala 27:72]
  wire  _T_21997 = bht_rd_addr_hashed_f == 8'h14; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_22489 = _T_21997 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22744 = _T_22743 | _T_22489; // @[Mux.scala 27:72]
  wire  _T_21999 = bht_rd_addr_hashed_f == 8'h15; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_22490 = _T_21999 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22745 = _T_22744 | _T_22490; // @[Mux.scala 27:72]
  wire  _T_22001 = bht_rd_addr_hashed_f == 8'h16; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_22491 = _T_22001 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22746 = _T_22745 | _T_22491; // @[Mux.scala 27:72]
  wire  _T_22003 = bht_rd_addr_hashed_f == 8'h17; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_22492 = _T_22003 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22747 = _T_22746 | _T_22492; // @[Mux.scala 27:72]
  wire  _T_22005 = bht_rd_addr_hashed_f == 8'h18; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_22493 = _T_22005 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22748 = _T_22747 | _T_22493; // @[Mux.scala 27:72]
  wire  _T_22007 = bht_rd_addr_hashed_f == 8'h19; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_22494 = _T_22007 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22749 = _T_22748 | _T_22494; // @[Mux.scala 27:72]
  wire  _T_22009 = bht_rd_addr_hashed_f == 8'h1a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_22495 = _T_22009 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22750 = _T_22749 | _T_22495; // @[Mux.scala 27:72]
  wire  _T_22011 = bht_rd_addr_hashed_f == 8'h1b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_22496 = _T_22011 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22751 = _T_22750 | _T_22496; // @[Mux.scala 27:72]
  wire  _T_22013 = bht_rd_addr_hashed_f == 8'h1c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_22497 = _T_22013 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22752 = _T_22751 | _T_22497; // @[Mux.scala 27:72]
  wire  _T_22015 = bht_rd_addr_hashed_f == 8'h1d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_22498 = _T_22015 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22753 = _T_22752 | _T_22498; // @[Mux.scala 27:72]
  wire  _T_22017 = bht_rd_addr_hashed_f == 8'h1e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_22499 = _T_22017 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22754 = _T_22753 | _T_22499; // @[Mux.scala 27:72]
  wire  _T_22019 = bht_rd_addr_hashed_f == 8'h1f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_22500 = _T_22019 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22755 = _T_22754 | _T_22500; // @[Mux.scala 27:72]
  wire  _T_22021 = bht_rd_addr_hashed_f == 8'h20; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_22501 = _T_22021 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22756 = _T_22755 | _T_22501; // @[Mux.scala 27:72]
  wire  _T_22023 = bht_rd_addr_hashed_f == 8'h21; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_22502 = _T_22023 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22757 = _T_22756 | _T_22502; // @[Mux.scala 27:72]
  wire  _T_22025 = bht_rd_addr_hashed_f == 8'h22; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_22503 = _T_22025 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22758 = _T_22757 | _T_22503; // @[Mux.scala 27:72]
  wire  _T_22027 = bht_rd_addr_hashed_f == 8'h23; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_22504 = _T_22027 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22759 = _T_22758 | _T_22504; // @[Mux.scala 27:72]
  wire  _T_22029 = bht_rd_addr_hashed_f == 8'h24; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_22505 = _T_22029 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22760 = _T_22759 | _T_22505; // @[Mux.scala 27:72]
  wire  _T_22031 = bht_rd_addr_hashed_f == 8'h25; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_22506 = _T_22031 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22761 = _T_22760 | _T_22506; // @[Mux.scala 27:72]
  wire  _T_22033 = bht_rd_addr_hashed_f == 8'h26; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_22507 = _T_22033 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22762 = _T_22761 | _T_22507; // @[Mux.scala 27:72]
  wire  _T_22035 = bht_rd_addr_hashed_f == 8'h27; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_22508 = _T_22035 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22763 = _T_22762 | _T_22508; // @[Mux.scala 27:72]
  wire  _T_22037 = bht_rd_addr_hashed_f == 8'h28; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_22509 = _T_22037 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22764 = _T_22763 | _T_22509; // @[Mux.scala 27:72]
  wire  _T_22039 = bht_rd_addr_hashed_f == 8'h29; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_22510 = _T_22039 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22765 = _T_22764 | _T_22510; // @[Mux.scala 27:72]
  wire  _T_22041 = bht_rd_addr_hashed_f == 8'h2a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_22511 = _T_22041 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22766 = _T_22765 | _T_22511; // @[Mux.scala 27:72]
  wire  _T_22043 = bht_rd_addr_hashed_f == 8'h2b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_22512 = _T_22043 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22767 = _T_22766 | _T_22512; // @[Mux.scala 27:72]
  wire  _T_22045 = bht_rd_addr_hashed_f == 8'h2c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_22513 = _T_22045 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22768 = _T_22767 | _T_22513; // @[Mux.scala 27:72]
  wire  _T_22047 = bht_rd_addr_hashed_f == 8'h2d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_22514 = _T_22047 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22769 = _T_22768 | _T_22514; // @[Mux.scala 27:72]
  wire  _T_22049 = bht_rd_addr_hashed_f == 8'h2e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_22515 = _T_22049 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22770 = _T_22769 | _T_22515; // @[Mux.scala 27:72]
  wire  _T_22051 = bht_rd_addr_hashed_f == 8'h2f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_22516 = _T_22051 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22771 = _T_22770 | _T_22516; // @[Mux.scala 27:72]
  wire  _T_22053 = bht_rd_addr_hashed_f == 8'h30; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_22517 = _T_22053 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22772 = _T_22771 | _T_22517; // @[Mux.scala 27:72]
  wire  _T_22055 = bht_rd_addr_hashed_f == 8'h31; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_22518 = _T_22055 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22773 = _T_22772 | _T_22518; // @[Mux.scala 27:72]
  wire  _T_22057 = bht_rd_addr_hashed_f == 8'h32; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_22519 = _T_22057 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22774 = _T_22773 | _T_22519; // @[Mux.scala 27:72]
  wire  _T_22059 = bht_rd_addr_hashed_f == 8'h33; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_22520 = _T_22059 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22775 = _T_22774 | _T_22520; // @[Mux.scala 27:72]
  wire  _T_22061 = bht_rd_addr_hashed_f == 8'h34; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_22521 = _T_22061 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22776 = _T_22775 | _T_22521; // @[Mux.scala 27:72]
  wire  _T_22063 = bht_rd_addr_hashed_f == 8'h35; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_22522 = _T_22063 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22777 = _T_22776 | _T_22522; // @[Mux.scala 27:72]
  wire  _T_22065 = bht_rd_addr_hashed_f == 8'h36; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_22523 = _T_22065 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22778 = _T_22777 | _T_22523; // @[Mux.scala 27:72]
  wire  _T_22067 = bht_rd_addr_hashed_f == 8'h37; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_22524 = _T_22067 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22779 = _T_22778 | _T_22524; // @[Mux.scala 27:72]
  wire  _T_22069 = bht_rd_addr_hashed_f == 8'h38; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_22525 = _T_22069 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22780 = _T_22779 | _T_22525; // @[Mux.scala 27:72]
  wire  _T_22071 = bht_rd_addr_hashed_f == 8'h39; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_22526 = _T_22071 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22781 = _T_22780 | _T_22526; // @[Mux.scala 27:72]
  wire  _T_22073 = bht_rd_addr_hashed_f == 8'h3a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_22527 = _T_22073 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22782 = _T_22781 | _T_22527; // @[Mux.scala 27:72]
  wire  _T_22075 = bht_rd_addr_hashed_f == 8'h3b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_22528 = _T_22075 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22783 = _T_22782 | _T_22528; // @[Mux.scala 27:72]
  wire  _T_22077 = bht_rd_addr_hashed_f == 8'h3c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_22529 = _T_22077 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22784 = _T_22783 | _T_22529; // @[Mux.scala 27:72]
  wire  _T_22079 = bht_rd_addr_hashed_f == 8'h3d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_22530 = _T_22079 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22785 = _T_22784 | _T_22530; // @[Mux.scala 27:72]
  wire  _T_22081 = bht_rd_addr_hashed_f == 8'h3e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_22531 = _T_22081 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22786 = _T_22785 | _T_22531; // @[Mux.scala 27:72]
  wire  _T_22083 = bht_rd_addr_hashed_f == 8'h3f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_22532 = _T_22083 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22787 = _T_22786 | _T_22532; // @[Mux.scala 27:72]
  wire  _T_22085 = bht_rd_addr_hashed_f == 8'h40; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_22533 = _T_22085 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22788 = _T_22787 | _T_22533; // @[Mux.scala 27:72]
  wire  _T_22087 = bht_rd_addr_hashed_f == 8'h41; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_22534 = _T_22087 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22789 = _T_22788 | _T_22534; // @[Mux.scala 27:72]
  wire  _T_22089 = bht_rd_addr_hashed_f == 8'h42; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_22535 = _T_22089 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22790 = _T_22789 | _T_22535; // @[Mux.scala 27:72]
  wire  _T_22091 = bht_rd_addr_hashed_f == 8'h43; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_22536 = _T_22091 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22791 = _T_22790 | _T_22536; // @[Mux.scala 27:72]
  wire  _T_22093 = bht_rd_addr_hashed_f == 8'h44; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_22537 = _T_22093 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22792 = _T_22791 | _T_22537; // @[Mux.scala 27:72]
  wire  _T_22095 = bht_rd_addr_hashed_f == 8'h45; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_22538 = _T_22095 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22793 = _T_22792 | _T_22538; // @[Mux.scala 27:72]
  wire  _T_22097 = bht_rd_addr_hashed_f == 8'h46; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_22539 = _T_22097 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22794 = _T_22793 | _T_22539; // @[Mux.scala 27:72]
  wire  _T_22099 = bht_rd_addr_hashed_f == 8'h47; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_22540 = _T_22099 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22795 = _T_22794 | _T_22540; // @[Mux.scala 27:72]
  wire  _T_22101 = bht_rd_addr_hashed_f == 8'h48; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_22541 = _T_22101 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22796 = _T_22795 | _T_22541; // @[Mux.scala 27:72]
  wire  _T_22103 = bht_rd_addr_hashed_f == 8'h49; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_22542 = _T_22103 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22797 = _T_22796 | _T_22542; // @[Mux.scala 27:72]
  wire  _T_22105 = bht_rd_addr_hashed_f == 8'h4a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_22543 = _T_22105 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22798 = _T_22797 | _T_22543; // @[Mux.scala 27:72]
  wire  _T_22107 = bht_rd_addr_hashed_f == 8'h4b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_22544 = _T_22107 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22799 = _T_22798 | _T_22544; // @[Mux.scala 27:72]
  wire  _T_22109 = bht_rd_addr_hashed_f == 8'h4c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_22545 = _T_22109 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22800 = _T_22799 | _T_22545; // @[Mux.scala 27:72]
  wire  _T_22111 = bht_rd_addr_hashed_f == 8'h4d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_22546 = _T_22111 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22801 = _T_22800 | _T_22546; // @[Mux.scala 27:72]
  wire  _T_22113 = bht_rd_addr_hashed_f == 8'h4e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_22547 = _T_22113 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22802 = _T_22801 | _T_22547; // @[Mux.scala 27:72]
  wire  _T_22115 = bht_rd_addr_hashed_f == 8'h4f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_22548 = _T_22115 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22803 = _T_22802 | _T_22548; // @[Mux.scala 27:72]
  wire  _T_22117 = bht_rd_addr_hashed_f == 8'h50; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_22549 = _T_22117 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22804 = _T_22803 | _T_22549; // @[Mux.scala 27:72]
  wire  _T_22119 = bht_rd_addr_hashed_f == 8'h51; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_22550 = _T_22119 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22805 = _T_22804 | _T_22550; // @[Mux.scala 27:72]
  wire  _T_22121 = bht_rd_addr_hashed_f == 8'h52; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_22551 = _T_22121 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22806 = _T_22805 | _T_22551; // @[Mux.scala 27:72]
  wire  _T_22123 = bht_rd_addr_hashed_f == 8'h53; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_22552 = _T_22123 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22807 = _T_22806 | _T_22552; // @[Mux.scala 27:72]
  wire  _T_22125 = bht_rd_addr_hashed_f == 8'h54; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_22553 = _T_22125 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22808 = _T_22807 | _T_22553; // @[Mux.scala 27:72]
  wire  _T_22127 = bht_rd_addr_hashed_f == 8'h55; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_22554 = _T_22127 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22809 = _T_22808 | _T_22554; // @[Mux.scala 27:72]
  wire  _T_22129 = bht_rd_addr_hashed_f == 8'h56; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_22555 = _T_22129 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22810 = _T_22809 | _T_22555; // @[Mux.scala 27:72]
  wire  _T_22131 = bht_rd_addr_hashed_f == 8'h57; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_22556 = _T_22131 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22811 = _T_22810 | _T_22556; // @[Mux.scala 27:72]
  wire  _T_22133 = bht_rd_addr_hashed_f == 8'h58; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_22557 = _T_22133 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22812 = _T_22811 | _T_22557; // @[Mux.scala 27:72]
  wire  _T_22135 = bht_rd_addr_hashed_f == 8'h59; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_22558 = _T_22135 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22813 = _T_22812 | _T_22558; // @[Mux.scala 27:72]
  wire  _T_22137 = bht_rd_addr_hashed_f == 8'h5a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_22559 = _T_22137 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22814 = _T_22813 | _T_22559; // @[Mux.scala 27:72]
  wire  _T_22139 = bht_rd_addr_hashed_f == 8'h5b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_22560 = _T_22139 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22815 = _T_22814 | _T_22560; // @[Mux.scala 27:72]
  wire  _T_22141 = bht_rd_addr_hashed_f == 8'h5c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_22561 = _T_22141 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22816 = _T_22815 | _T_22561; // @[Mux.scala 27:72]
  wire  _T_22143 = bht_rd_addr_hashed_f == 8'h5d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_22562 = _T_22143 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22817 = _T_22816 | _T_22562; // @[Mux.scala 27:72]
  wire  _T_22145 = bht_rd_addr_hashed_f == 8'h5e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_22563 = _T_22145 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22818 = _T_22817 | _T_22563; // @[Mux.scala 27:72]
  wire  _T_22147 = bht_rd_addr_hashed_f == 8'h5f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_22564 = _T_22147 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22819 = _T_22818 | _T_22564; // @[Mux.scala 27:72]
  wire  _T_22149 = bht_rd_addr_hashed_f == 8'h60; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_22565 = _T_22149 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22820 = _T_22819 | _T_22565; // @[Mux.scala 27:72]
  wire  _T_22151 = bht_rd_addr_hashed_f == 8'h61; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_22566 = _T_22151 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22821 = _T_22820 | _T_22566; // @[Mux.scala 27:72]
  wire  _T_22153 = bht_rd_addr_hashed_f == 8'h62; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_22567 = _T_22153 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22822 = _T_22821 | _T_22567; // @[Mux.scala 27:72]
  wire  _T_22155 = bht_rd_addr_hashed_f == 8'h63; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_22568 = _T_22155 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22823 = _T_22822 | _T_22568; // @[Mux.scala 27:72]
  wire  _T_22157 = bht_rd_addr_hashed_f == 8'h64; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_22569 = _T_22157 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22824 = _T_22823 | _T_22569; // @[Mux.scala 27:72]
  wire  _T_22159 = bht_rd_addr_hashed_f == 8'h65; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_22570 = _T_22159 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22825 = _T_22824 | _T_22570; // @[Mux.scala 27:72]
  wire  _T_22161 = bht_rd_addr_hashed_f == 8'h66; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_22571 = _T_22161 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22826 = _T_22825 | _T_22571; // @[Mux.scala 27:72]
  wire  _T_22163 = bht_rd_addr_hashed_f == 8'h67; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_22572 = _T_22163 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22827 = _T_22826 | _T_22572; // @[Mux.scala 27:72]
  wire  _T_22165 = bht_rd_addr_hashed_f == 8'h68; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_22573 = _T_22165 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22828 = _T_22827 | _T_22573; // @[Mux.scala 27:72]
  wire  _T_22167 = bht_rd_addr_hashed_f == 8'h69; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_22574 = _T_22167 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22829 = _T_22828 | _T_22574; // @[Mux.scala 27:72]
  wire  _T_22169 = bht_rd_addr_hashed_f == 8'h6a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_22575 = _T_22169 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22830 = _T_22829 | _T_22575; // @[Mux.scala 27:72]
  wire  _T_22171 = bht_rd_addr_hashed_f == 8'h6b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_22576 = _T_22171 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22831 = _T_22830 | _T_22576; // @[Mux.scala 27:72]
  wire  _T_22173 = bht_rd_addr_hashed_f == 8'h6c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_22577 = _T_22173 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22832 = _T_22831 | _T_22577; // @[Mux.scala 27:72]
  wire  _T_22175 = bht_rd_addr_hashed_f == 8'h6d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_22578 = _T_22175 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22833 = _T_22832 | _T_22578; // @[Mux.scala 27:72]
  wire  _T_22177 = bht_rd_addr_hashed_f == 8'h6e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_22579 = _T_22177 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22834 = _T_22833 | _T_22579; // @[Mux.scala 27:72]
  wire  _T_22179 = bht_rd_addr_hashed_f == 8'h6f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_22580 = _T_22179 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22835 = _T_22834 | _T_22580; // @[Mux.scala 27:72]
  wire  _T_22181 = bht_rd_addr_hashed_f == 8'h70; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_22581 = _T_22181 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22836 = _T_22835 | _T_22581; // @[Mux.scala 27:72]
  wire  _T_22183 = bht_rd_addr_hashed_f == 8'h71; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_22582 = _T_22183 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22837 = _T_22836 | _T_22582; // @[Mux.scala 27:72]
  wire  _T_22185 = bht_rd_addr_hashed_f == 8'h72; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_22583 = _T_22185 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22838 = _T_22837 | _T_22583; // @[Mux.scala 27:72]
  wire  _T_22187 = bht_rd_addr_hashed_f == 8'h73; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_22584 = _T_22187 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22839 = _T_22838 | _T_22584; // @[Mux.scala 27:72]
  wire  _T_22189 = bht_rd_addr_hashed_f == 8'h74; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_22585 = _T_22189 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22840 = _T_22839 | _T_22585; // @[Mux.scala 27:72]
  wire  _T_22191 = bht_rd_addr_hashed_f == 8'h75; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_22586 = _T_22191 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22841 = _T_22840 | _T_22586; // @[Mux.scala 27:72]
  wire  _T_22193 = bht_rd_addr_hashed_f == 8'h76; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_22587 = _T_22193 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22842 = _T_22841 | _T_22587; // @[Mux.scala 27:72]
  wire  _T_22195 = bht_rd_addr_hashed_f == 8'h77; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_22588 = _T_22195 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22843 = _T_22842 | _T_22588; // @[Mux.scala 27:72]
  wire  _T_22197 = bht_rd_addr_hashed_f == 8'h78; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_22589 = _T_22197 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22844 = _T_22843 | _T_22589; // @[Mux.scala 27:72]
  wire  _T_22199 = bht_rd_addr_hashed_f == 8'h79; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_22590 = _T_22199 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22845 = _T_22844 | _T_22590; // @[Mux.scala 27:72]
  wire  _T_22201 = bht_rd_addr_hashed_f == 8'h7a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_22591 = _T_22201 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22846 = _T_22845 | _T_22591; // @[Mux.scala 27:72]
  wire  _T_22203 = bht_rd_addr_hashed_f == 8'h7b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_22592 = _T_22203 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22847 = _T_22846 | _T_22592; // @[Mux.scala 27:72]
  wire  _T_22205 = bht_rd_addr_hashed_f == 8'h7c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_22593 = _T_22205 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22848 = _T_22847 | _T_22593; // @[Mux.scala 27:72]
  wire  _T_22207 = bht_rd_addr_hashed_f == 8'h7d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_22594 = _T_22207 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22849 = _T_22848 | _T_22594; // @[Mux.scala 27:72]
  wire  _T_22209 = bht_rd_addr_hashed_f == 8'h7e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_22595 = _T_22209 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22850 = _T_22849 | _T_22595; // @[Mux.scala 27:72]
  wire  _T_22211 = bht_rd_addr_hashed_f == 8'h7f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_22596 = _T_22211 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22851 = _T_22850 | _T_22596; // @[Mux.scala 27:72]
  wire  _T_22213 = bht_rd_addr_hashed_f == 8'h80; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_22597 = _T_22213 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22852 = _T_22851 | _T_22597; // @[Mux.scala 27:72]
  wire  _T_22215 = bht_rd_addr_hashed_f == 8'h81; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_22598 = _T_22215 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22853 = _T_22852 | _T_22598; // @[Mux.scala 27:72]
  wire  _T_22217 = bht_rd_addr_hashed_f == 8'h82; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_22599 = _T_22217 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22854 = _T_22853 | _T_22599; // @[Mux.scala 27:72]
  wire  _T_22219 = bht_rd_addr_hashed_f == 8'h83; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_22600 = _T_22219 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22855 = _T_22854 | _T_22600; // @[Mux.scala 27:72]
  wire  _T_22221 = bht_rd_addr_hashed_f == 8'h84; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_22601 = _T_22221 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22856 = _T_22855 | _T_22601; // @[Mux.scala 27:72]
  wire  _T_22223 = bht_rd_addr_hashed_f == 8'h85; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_22602 = _T_22223 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22857 = _T_22856 | _T_22602; // @[Mux.scala 27:72]
  wire  _T_22225 = bht_rd_addr_hashed_f == 8'h86; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_22603 = _T_22225 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22858 = _T_22857 | _T_22603; // @[Mux.scala 27:72]
  wire  _T_22227 = bht_rd_addr_hashed_f == 8'h87; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_22604 = _T_22227 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22859 = _T_22858 | _T_22604; // @[Mux.scala 27:72]
  wire  _T_22229 = bht_rd_addr_hashed_f == 8'h88; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_22605 = _T_22229 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22860 = _T_22859 | _T_22605; // @[Mux.scala 27:72]
  wire  _T_22231 = bht_rd_addr_hashed_f == 8'h89; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_22606 = _T_22231 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22861 = _T_22860 | _T_22606; // @[Mux.scala 27:72]
  wire  _T_22233 = bht_rd_addr_hashed_f == 8'h8a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_22607 = _T_22233 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22862 = _T_22861 | _T_22607; // @[Mux.scala 27:72]
  wire  _T_22235 = bht_rd_addr_hashed_f == 8'h8b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_22608 = _T_22235 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22863 = _T_22862 | _T_22608; // @[Mux.scala 27:72]
  wire  _T_22237 = bht_rd_addr_hashed_f == 8'h8c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_22609 = _T_22237 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22864 = _T_22863 | _T_22609; // @[Mux.scala 27:72]
  wire  _T_22239 = bht_rd_addr_hashed_f == 8'h8d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_22610 = _T_22239 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22865 = _T_22864 | _T_22610; // @[Mux.scala 27:72]
  wire  _T_22241 = bht_rd_addr_hashed_f == 8'h8e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_22611 = _T_22241 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22866 = _T_22865 | _T_22611; // @[Mux.scala 27:72]
  wire  _T_22243 = bht_rd_addr_hashed_f == 8'h8f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_22612 = _T_22243 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22867 = _T_22866 | _T_22612; // @[Mux.scala 27:72]
  wire  _T_22245 = bht_rd_addr_hashed_f == 8'h90; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_22613 = _T_22245 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22868 = _T_22867 | _T_22613; // @[Mux.scala 27:72]
  wire  _T_22247 = bht_rd_addr_hashed_f == 8'h91; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_22614 = _T_22247 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22869 = _T_22868 | _T_22614; // @[Mux.scala 27:72]
  wire  _T_22249 = bht_rd_addr_hashed_f == 8'h92; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_22615 = _T_22249 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22870 = _T_22869 | _T_22615; // @[Mux.scala 27:72]
  wire  _T_22251 = bht_rd_addr_hashed_f == 8'h93; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_22616 = _T_22251 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22871 = _T_22870 | _T_22616; // @[Mux.scala 27:72]
  wire  _T_22253 = bht_rd_addr_hashed_f == 8'h94; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_22617 = _T_22253 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22872 = _T_22871 | _T_22617; // @[Mux.scala 27:72]
  wire  _T_22255 = bht_rd_addr_hashed_f == 8'h95; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_22618 = _T_22255 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22873 = _T_22872 | _T_22618; // @[Mux.scala 27:72]
  wire  _T_22257 = bht_rd_addr_hashed_f == 8'h96; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_22619 = _T_22257 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22874 = _T_22873 | _T_22619; // @[Mux.scala 27:72]
  wire  _T_22259 = bht_rd_addr_hashed_f == 8'h97; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_22620 = _T_22259 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22875 = _T_22874 | _T_22620; // @[Mux.scala 27:72]
  wire  _T_22261 = bht_rd_addr_hashed_f == 8'h98; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_22621 = _T_22261 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22876 = _T_22875 | _T_22621; // @[Mux.scala 27:72]
  wire  _T_22263 = bht_rd_addr_hashed_f == 8'h99; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_22622 = _T_22263 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22877 = _T_22876 | _T_22622; // @[Mux.scala 27:72]
  wire  _T_22265 = bht_rd_addr_hashed_f == 8'h9a; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_22623 = _T_22265 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22878 = _T_22877 | _T_22623; // @[Mux.scala 27:72]
  wire  _T_22267 = bht_rd_addr_hashed_f == 8'h9b; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_22624 = _T_22267 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22879 = _T_22878 | _T_22624; // @[Mux.scala 27:72]
  wire  _T_22269 = bht_rd_addr_hashed_f == 8'h9c; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_22625 = _T_22269 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22880 = _T_22879 | _T_22625; // @[Mux.scala 27:72]
  wire  _T_22271 = bht_rd_addr_hashed_f == 8'h9d; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_22626 = _T_22271 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22881 = _T_22880 | _T_22626; // @[Mux.scala 27:72]
  wire  _T_22273 = bht_rd_addr_hashed_f == 8'h9e; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_22627 = _T_22273 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22882 = _T_22881 | _T_22627; // @[Mux.scala 27:72]
  wire  _T_22275 = bht_rd_addr_hashed_f == 8'h9f; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_22628 = _T_22275 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22883 = _T_22882 | _T_22628; // @[Mux.scala 27:72]
  wire  _T_22277 = bht_rd_addr_hashed_f == 8'ha0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_22629 = _T_22277 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22884 = _T_22883 | _T_22629; // @[Mux.scala 27:72]
  wire  _T_22279 = bht_rd_addr_hashed_f == 8'ha1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_22630 = _T_22279 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22885 = _T_22884 | _T_22630; // @[Mux.scala 27:72]
  wire  _T_22281 = bht_rd_addr_hashed_f == 8'ha2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_22631 = _T_22281 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22886 = _T_22885 | _T_22631; // @[Mux.scala 27:72]
  wire  _T_22283 = bht_rd_addr_hashed_f == 8'ha3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_22632 = _T_22283 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22887 = _T_22886 | _T_22632; // @[Mux.scala 27:72]
  wire  _T_22285 = bht_rd_addr_hashed_f == 8'ha4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_22633 = _T_22285 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22888 = _T_22887 | _T_22633; // @[Mux.scala 27:72]
  wire  _T_22287 = bht_rd_addr_hashed_f == 8'ha5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_22634 = _T_22287 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22889 = _T_22888 | _T_22634; // @[Mux.scala 27:72]
  wire  _T_22289 = bht_rd_addr_hashed_f == 8'ha6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_22635 = _T_22289 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22890 = _T_22889 | _T_22635; // @[Mux.scala 27:72]
  wire  _T_22291 = bht_rd_addr_hashed_f == 8'ha7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_22636 = _T_22291 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22891 = _T_22890 | _T_22636; // @[Mux.scala 27:72]
  wire  _T_22293 = bht_rd_addr_hashed_f == 8'ha8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_22637 = _T_22293 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22892 = _T_22891 | _T_22637; // @[Mux.scala 27:72]
  wire  _T_22295 = bht_rd_addr_hashed_f == 8'ha9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_22638 = _T_22295 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22893 = _T_22892 | _T_22638; // @[Mux.scala 27:72]
  wire  _T_22297 = bht_rd_addr_hashed_f == 8'haa; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_22639 = _T_22297 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22894 = _T_22893 | _T_22639; // @[Mux.scala 27:72]
  wire  _T_22299 = bht_rd_addr_hashed_f == 8'hab; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_22640 = _T_22299 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22895 = _T_22894 | _T_22640; // @[Mux.scala 27:72]
  wire  _T_22301 = bht_rd_addr_hashed_f == 8'hac; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_22641 = _T_22301 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22896 = _T_22895 | _T_22641; // @[Mux.scala 27:72]
  wire  _T_22303 = bht_rd_addr_hashed_f == 8'had; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_22642 = _T_22303 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22897 = _T_22896 | _T_22642; // @[Mux.scala 27:72]
  wire  _T_22305 = bht_rd_addr_hashed_f == 8'hae; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_22643 = _T_22305 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22898 = _T_22897 | _T_22643; // @[Mux.scala 27:72]
  wire  _T_22307 = bht_rd_addr_hashed_f == 8'haf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_22644 = _T_22307 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22899 = _T_22898 | _T_22644; // @[Mux.scala 27:72]
  wire  _T_22309 = bht_rd_addr_hashed_f == 8'hb0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_22645 = _T_22309 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22900 = _T_22899 | _T_22645; // @[Mux.scala 27:72]
  wire  _T_22311 = bht_rd_addr_hashed_f == 8'hb1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_22646 = _T_22311 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22901 = _T_22900 | _T_22646; // @[Mux.scala 27:72]
  wire  _T_22313 = bht_rd_addr_hashed_f == 8'hb2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_22647 = _T_22313 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22902 = _T_22901 | _T_22647; // @[Mux.scala 27:72]
  wire  _T_22315 = bht_rd_addr_hashed_f == 8'hb3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_22648 = _T_22315 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22903 = _T_22902 | _T_22648; // @[Mux.scala 27:72]
  wire  _T_22317 = bht_rd_addr_hashed_f == 8'hb4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_22649 = _T_22317 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22904 = _T_22903 | _T_22649; // @[Mux.scala 27:72]
  wire  _T_22319 = bht_rd_addr_hashed_f == 8'hb5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_22650 = _T_22319 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22905 = _T_22904 | _T_22650; // @[Mux.scala 27:72]
  wire  _T_22321 = bht_rd_addr_hashed_f == 8'hb6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_22651 = _T_22321 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22906 = _T_22905 | _T_22651; // @[Mux.scala 27:72]
  wire  _T_22323 = bht_rd_addr_hashed_f == 8'hb7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_22652 = _T_22323 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22907 = _T_22906 | _T_22652; // @[Mux.scala 27:72]
  wire  _T_22325 = bht_rd_addr_hashed_f == 8'hb8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_22653 = _T_22325 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22908 = _T_22907 | _T_22653; // @[Mux.scala 27:72]
  wire  _T_22327 = bht_rd_addr_hashed_f == 8'hb9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_22654 = _T_22327 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22909 = _T_22908 | _T_22654; // @[Mux.scala 27:72]
  wire  _T_22329 = bht_rd_addr_hashed_f == 8'hba; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_22655 = _T_22329 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22910 = _T_22909 | _T_22655; // @[Mux.scala 27:72]
  wire  _T_22331 = bht_rd_addr_hashed_f == 8'hbb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_22656 = _T_22331 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22911 = _T_22910 | _T_22656; // @[Mux.scala 27:72]
  wire  _T_22333 = bht_rd_addr_hashed_f == 8'hbc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_22657 = _T_22333 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22912 = _T_22911 | _T_22657; // @[Mux.scala 27:72]
  wire  _T_22335 = bht_rd_addr_hashed_f == 8'hbd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_22658 = _T_22335 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22913 = _T_22912 | _T_22658; // @[Mux.scala 27:72]
  wire  _T_22337 = bht_rd_addr_hashed_f == 8'hbe; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_22659 = _T_22337 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22914 = _T_22913 | _T_22659; // @[Mux.scala 27:72]
  wire  _T_22339 = bht_rd_addr_hashed_f == 8'hbf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_22660 = _T_22339 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22915 = _T_22914 | _T_22660; // @[Mux.scala 27:72]
  wire  _T_22341 = bht_rd_addr_hashed_f == 8'hc0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_22661 = _T_22341 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22916 = _T_22915 | _T_22661; // @[Mux.scala 27:72]
  wire  _T_22343 = bht_rd_addr_hashed_f == 8'hc1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_22662 = _T_22343 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22917 = _T_22916 | _T_22662; // @[Mux.scala 27:72]
  wire  _T_22345 = bht_rd_addr_hashed_f == 8'hc2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_22663 = _T_22345 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22918 = _T_22917 | _T_22663; // @[Mux.scala 27:72]
  wire  _T_22347 = bht_rd_addr_hashed_f == 8'hc3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_22664 = _T_22347 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22919 = _T_22918 | _T_22664; // @[Mux.scala 27:72]
  wire  _T_22349 = bht_rd_addr_hashed_f == 8'hc4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_22665 = _T_22349 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22920 = _T_22919 | _T_22665; // @[Mux.scala 27:72]
  wire  _T_22351 = bht_rd_addr_hashed_f == 8'hc5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_22666 = _T_22351 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22921 = _T_22920 | _T_22666; // @[Mux.scala 27:72]
  wire  _T_22353 = bht_rd_addr_hashed_f == 8'hc6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_22667 = _T_22353 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22922 = _T_22921 | _T_22667; // @[Mux.scala 27:72]
  wire  _T_22355 = bht_rd_addr_hashed_f == 8'hc7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_22668 = _T_22355 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22923 = _T_22922 | _T_22668; // @[Mux.scala 27:72]
  wire  _T_22357 = bht_rd_addr_hashed_f == 8'hc8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_22669 = _T_22357 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22924 = _T_22923 | _T_22669; // @[Mux.scala 27:72]
  wire  _T_22359 = bht_rd_addr_hashed_f == 8'hc9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_22670 = _T_22359 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22925 = _T_22924 | _T_22670; // @[Mux.scala 27:72]
  wire  _T_22361 = bht_rd_addr_hashed_f == 8'hca; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_22671 = _T_22361 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22926 = _T_22925 | _T_22671; // @[Mux.scala 27:72]
  wire  _T_22363 = bht_rd_addr_hashed_f == 8'hcb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_22672 = _T_22363 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22927 = _T_22926 | _T_22672; // @[Mux.scala 27:72]
  wire  _T_22365 = bht_rd_addr_hashed_f == 8'hcc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_22673 = _T_22365 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22928 = _T_22927 | _T_22673; // @[Mux.scala 27:72]
  wire  _T_22367 = bht_rd_addr_hashed_f == 8'hcd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_22674 = _T_22367 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22929 = _T_22928 | _T_22674; // @[Mux.scala 27:72]
  wire  _T_22369 = bht_rd_addr_hashed_f == 8'hce; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_22675 = _T_22369 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22930 = _T_22929 | _T_22675; // @[Mux.scala 27:72]
  wire  _T_22371 = bht_rd_addr_hashed_f == 8'hcf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_22676 = _T_22371 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22931 = _T_22930 | _T_22676; // @[Mux.scala 27:72]
  wire  _T_22373 = bht_rd_addr_hashed_f == 8'hd0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_22677 = _T_22373 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22932 = _T_22931 | _T_22677; // @[Mux.scala 27:72]
  wire  _T_22375 = bht_rd_addr_hashed_f == 8'hd1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_22678 = _T_22375 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22933 = _T_22932 | _T_22678; // @[Mux.scala 27:72]
  wire  _T_22377 = bht_rd_addr_hashed_f == 8'hd2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_22679 = _T_22377 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22934 = _T_22933 | _T_22679; // @[Mux.scala 27:72]
  wire  _T_22379 = bht_rd_addr_hashed_f == 8'hd3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_22680 = _T_22379 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22935 = _T_22934 | _T_22680; // @[Mux.scala 27:72]
  wire  _T_22381 = bht_rd_addr_hashed_f == 8'hd4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_22681 = _T_22381 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22936 = _T_22935 | _T_22681; // @[Mux.scala 27:72]
  wire  _T_22383 = bht_rd_addr_hashed_f == 8'hd5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_22682 = _T_22383 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22937 = _T_22936 | _T_22682; // @[Mux.scala 27:72]
  wire  _T_22385 = bht_rd_addr_hashed_f == 8'hd6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_22683 = _T_22385 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22938 = _T_22937 | _T_22683; // @[Mux.scala 27:72]
  wire  _T_22387 = bht_rd_addr_hashed_f == 8'hd7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_22684 = _T_22387 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22939 = _T_22938 | _T_22684; // @[Mux.scala 27:72]
  wire  _T_22389 = bht_rd_addr_hashed_f == 8'hd8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_22685 = _T_22389 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22940 = _T_22939 | _T_22685; // @[Mux.scala 27:72]
  wire  _T_22391 = bht_rd_addr_hashed_f == 8'hd9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_22686 = _T_22391 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22941 = _T_22940 | _T_22686; // @[Mux.scala 27:72]
  wire  _T_22393 = bht_rd_addr_hashed_f == 8'hda; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_22687 = _T_22393 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22942 = _T_22941 | _T_22687; // @[Mux.scala 27:72]
  wire  _T_22395 = bht_rd_addr_hashed_f == 8'hdb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_22688 = _T_22395 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22943 = _T_22942 | _T_22688; // @[Mux.scala 27:72]
  wire  _T_22397 = bht_rd_addr_hashed_f == 8'hdc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_22689 = _T_22397 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22944 = _T_22943 | _T_22689; // @[Mux.scala 27:72]
  wire  _T_22399 = bht_rd_addr_hashed_f == 8'hdd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_22690 = _T_22399 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22945 = _T_22944 | _T_22690; // @[Mux.scala 27:72]
  wire  _T_22401 = bht_rd_addr_hashed_f == 8'hde; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_22691 = _T_22401 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22946 = _T_22945 | _T_22691; // @[Mux.scala 27:72]
  wire  _T_22403 = bht_rd_addr_hashed_f == 8'hdf; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_22692 = _T_22403 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22947 = _T_22946 | _T_22692; // @[Mux.scala 27:72]
  wire  _T_22405 = bht_rd_addr_hashed_f == 8'he0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_22693 = _T_22405 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22948 = _T_22947 | _T_22693; // @[Mux.scala 27:72]
  wire  _T_22407 = bht_rd_addr_hashed_f == 8'he1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_22694 = _T_22407 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22949 = _T_22948 | _T_22694; // @[Mux.scala 27:72]
  wire  _T_22409 = bht_rd_addr_hashed_f == 8'he2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_22695 = _T_22409 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22950 = _T_22949 | _T_22695; // @[Mux.scala 27:72]
  wire  _T_22411 = bht_rd_addr_hashed_f == 8'he3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_22696 = _T_22411 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22951 = _T_22950 | _T_22696; // @[Mux.scala 27:72]
  wire  _T_22413 = bht_rd_addr_hashed_f == 8'he4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_22697 = _T_22413 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22952 = _T_22951 | _T_22697; // @[Mux.scala 27:72]
  wire  _T_22415 = bht_rd_addr_hashed_f == 8'he5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_22698 = _T_22415 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22953 = _T_22952 | _T_22698; // @[Mux.scala 27:72]
  wire  _T_22417 = bht_rd_addr_hashed_f == 8'he6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_22699 = _T_22417 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22954 = _T_22953 | _T_22699; // @[Mux.scala 27:72]
  wire  _T_22419 = bht_rd_addr_hashed_f == 8'he7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_22700 = _T_22419 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22955 = _T_22954 | _T_22700; // @[Mux.scala 27:72]
  wire  _T_22421 = bht_rd_addr_hashed_f == 8'he8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_22701 = _T_22421 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22956 = _T_22955 | _T_22701; // @[Mux.scala 27:72]
  wire  _T_22423 = bht_rd_addr_hashed_f == 8'he9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_22702 = _T_22423 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22957 = _T_22956 | _T_22702; // @[Mux.scala 27:72]
  wire  _T_22425 = bht_rd_addr_hashed_f == 8'hea; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_22703 = _T_22425 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22958 = _T_22957 | _T_22703; // @[Mux.scala 27:72]
  wire  _T_22427 = bht_rd_addr_hashed_f == 8'heb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_22704 = _T_22427 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22959 = _T_22958 | _T_22704; // @[Mux.scala 27:72]
  wire  _T_22429 = bht_rd_addr_hashed_f == 8'hec; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_22705 = _T_22429 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22960 = _T_22959 | _T_22705; // @[Mux.scala 27:72]
  wire  _T_22431 = bht_rd_addr_hashed_f == 8'hed; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_22706 = _T_22431 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22961 = _T_22960 | _T_22706; // @[Mux.scala 27:72]
  wire  _T_22433 = bht_rd_addr_hashed_f == 8'hee; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_22707 = _T_22433 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22962 = _T_22961 | _T_22707; // @[Mux.scala 27:72]
  wire  _T_22435 = bht_rd_addr_hashed_f == 8'hef; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_22708 = _T_22435 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22963 = _T_22962 | _T_22708; // @[Mux.scala 27:72]
  wire  _T_22437 = bht_rd_addr_hashed_f == 8'hf0; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_22709 = _T_22437 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22964 = _T_22963 | _T_22709; // @[Mux.scala 27:72]
  wire  _T_22439 = bht_rd_addr_hashed_f == 8'hf1; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_22710 = _T_22439 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22965 = _T_22964 | _T_22710; // @[Mux.scala 27:72]
  wire  _T_22441 = bht_rd_addr_hashed_f == 8'hf2; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_22711 = _T_22441 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22966 = _T_22965 | _T_22711; // @[Mux.scala 27:72]
  wire  _T_22443 = bht_rd_addr_hashed_f == 8'hf3; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_22712 = _T_22443 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22967 = _T_22966 | _T_22712; // @[Mux.scala 27:72]
  wire  _T_22445 = bht_rd_addr_hashed_f == 8'hf4; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_22713 = _T_22445 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22968 = _T_22967 | _T_22713; // @[Mux.scala 27:72]
  wire  _T_22447 = bht_rd_addr_hashed_f == 8'hf5; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_22714 = _T_22447 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22969 = _T_22968 | _T_22714; // @[Mux.scala 27:72]
  wire  _T_22449 = bht_rd_addr_hashed_f == 8'hf6; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_22715 = _T_22449 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22970 = _T_22969 | _T_22715; // @[Mux.scala 27:72]
  wire  _T_22451 = bht_rd_addr_hashed_f == 8'hf7; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_22716 = _T_22451 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22971 = _T_22970 | _T_22716; // @[Mux.scala 27:72]
  wire  _T_22453 = bht_rd_addr_hashed_f == 8'hf8; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_22717 = _T_22453 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22972 = _T_22971 | _T_22717; // @[Mux.scala 27:72]
  wire  _T_22455 = bht_rd_addr_hashed_f == 8'hf9; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_22718 = _T_22455 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22973 = _T_22972 | _T_22718; // @[Mux.scala 27:72]
  wire  _T_22457 = bht_rd_addr_hashed_f == 8'hfa; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_22719 = _T_22457 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22974 = _T_22973 | _T_22719; // @[Mux.scala 27:72]
  wire  _T_22459 = bht_rd_addr_hashed_f == 8'hfb; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_22720 = _T_22459 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22975 = _T_22974 | _T_22720; // @[Mux.scala 27:72]
  wire  _T_22461 = bht_rd_addr_hashed_f == 8'hfc; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_22721 = _T_22461 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22976 = _T_22975 | _T_22721; // @[Mux.scala 27:72]
  wire  _T_22463 = bht_rd_addr_hashed_f == 8'hfd; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_22722 = _T_22463 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22977 = _T_22976 | _T_22722; // @[Mux.scala 27:72]
  wire  _T_22465 = bht_rd_addr_hashed_f == 8'hfe; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_22723 = _T_22465 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22978 = _T_22977 | _T_22723; // @[Mux.scala 27:72]
  wire  _T_22467 = bht_rd_addr_hashed_f == 8'hff; // @[ifu_bp_ctl.scala 536:79]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_22724 = _T_22467 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_22978 | _T_22724; // @[Mux.scala 27:72]
  wire [1:0] _T_253 = _T_147 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_585 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_585[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_22981 = bht_rd_addr_hashed_p1_f == 8'h0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_23493 = _T_22981 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22983 = bht_rd_addr_hashed_p1_f == 8'h1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_23494 = _T_22983 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23749 = _T_23493 | _T_23494; // @[Mux.scala 27:72]
  wire  _T_22985 = bht_rd_addr_hashed_p1_f == 8'h2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_23495 = _T_22985 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23750 = _T_23749 | _T_23495; // @[Mux.scala 27:72]
  wire  _T_22987 = bht_rd_addr_hashed_p1_f == 8'h3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_23496 = _T_22987 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23751 = _T_23750 | _T_23496; // @[Mux.scala 27:72]
  wire  _T_22989 = bht_rd_addr_hashed_p1_f == 8'h4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_23497 = _T_22989 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23752 = _T_23751 | _T_23497; // @[Mux.scala 27:72]
  wire  _T_22991 = bht_rd_addr_hashed_p1_f == 8'h5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_23498 = _T_22991 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23753 = _T_23752 | _T_23498; // @[Mux.scala 27:72]
  wire  _T_22993 = bht_rd_addr_hashed_p1_f == 8'h6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_23499 = _T_22993 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23754 = _T_23753 | _T_23499; // @[Mux.scala 27:72]
  wire  _T_22995 = bht_rd_addr_hashed_p1_f == 8'h7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_23500 = _T_22995 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23755 = _T_23754 | _T_23500; // @[Mux.scala 27:72]
  wire  _T_22997 = bht_rd_addr_hashed_p1_f == 8'h8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_23501 = _T_22997 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23756 = _T_23755 | _T_23501; // @[Mux.scala 27:72]
  wire  _T_22999 = bht_rd_addr_hashed_p1_f == 8'h9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_23502 = _T_22999 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23757 = _T_23756 | _T_23502; // @[Mux.scala 27:72]
  wire  _T_23001 = bht_rd_addr_hashed_p1_f == 8'ha; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_23503 = _T_23001 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23758 = _T_23757 | _T_23503; // @[Mux.scala 27:72]
  wire  _T_23003 = bht_rd_addr_hashed_p1_f == 8'hb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_23504 = _T_23003 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23759 = _T_23758 | _T_23504; // @[Mux.scala 27:72]
  wire  _T_23005 = bht_rd_addr_hashed_p1_f == 8'hc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_23505 = _T_23005 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23760 = _T_23759 | _T_23505; // @[Mux.scala 27:72]
  wire  _T_23007 = bht_rd_addr_hashed_p1_f == 8'hd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_23506 = _T_23007 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23761 = _T_23760 | _T_23506; // @[Mux.scala 27:72]
  wire  _T_23009 = bht_rd_addr_hashed_p1_f == 8'he; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_23507 = _T_23009 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23762 = _T_23761 | _T_23507; // @[Mux.scala 27:72]
  wire  _T_23011 = bht_rd_addr_hashed_p1_f == 8'hf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_23508 = _T_23011 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23763 = _T_23762 | _T_23508; // @[Mux.scala 27:72]
  wire  _T_23013 = bht_rd_addr_hashed_p1_f == 8'h10; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_23509 = _T_23013 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23764 = _T_23763 | _T_23509; // @[Mux.scala 27:72]
  wire  _T_23015 = bht_rd_addr_hashed_p1_f == 8'h11; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_23510 = _T_23015 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23765 = _T_23764 | _T_23510; // @[Mux.scala 27:72]
  wire  _T_23017 = bht_rd_addr_hashed_p1_f == 8'h12; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_23511 = _T_23017 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23766 = _T_23765 | _T_23511; // @[Mux.scala 27:72]
  wire  _T_23019 = bht_rd_addr_hashed_p1_f == 8'h13; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_23512 = _T_23019 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23767 = _T_23766 | _T_23512; // @[Mux.scala 27:72]
  wire  _T_23021 = bht_rd_addr_hashed_p1_f == 8'h14; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_23513 = _T_23021 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23768 = _T_23767 | _T_23513; // @[Mux.scala 27:72]
  wire  _T_23023 = bht_rd_addr_hashed_p1_f == 8'h15; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_23514 = _T_23023 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23769 = _T_23768 | _T_23514; // @[Mux.scala 27:72]
  wire  _T_23025 = bht_rd_addr_hashed_p1_f == 8'h16; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_23515 = _T_23025 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23770 = _T_23769 | _T_23515; // @[Mux.scala 27:72]
  wire  _T_23027 = bht_rd_addr_hashed_p1_f == 8'h17; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_23516 = _T_23027 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23771 = _T_23770 | _T_23516; // @[Mux.scala 27:72]
  wire  _T_23029 = bht_rd_addr_hashed_p1_f == 8'h18; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_23517 = _T_23029 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23772 = _T_23771 | _T_23517; // @[Mux.scala 27:72]
  wire  _T_23031 = bht_rd_addr_hashed_p1_f == 8'h19; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_23518 = _T_23031 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23773 = _T_23772 | _T_23518; // @[Mux.scala 27:72]
  wire  _T_23033 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_23519 = _T_23033 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23774 = _T_23773 | _T_23519; // @[Mux.scala 27:72]
  wire  _T_23035 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_23520 = _T_23035 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23775 = _T_23774 | _T_23520; // @[Mux.scala 27:72]
  wire  _T_23037 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_23521 = _T_23037 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23776 = _T_23775 | _T_23521; // @[Mux.scala 27:72]
  wire  _T_23039 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_23522 = _T_23039 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23777 = _T_23776 | _T_23522; // @[Mux.scala 27:72]
  wire  _T_23041 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_23523 = _T_23041 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23778 = _T_23777 | _T_23523; // @[Mux.scala 27:72]
  wire  _T_23043 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_23524 = _T_23043 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23779 = _T_23778 | _T_23524; // @[Mux.scala 27:72]
  wire  _T_23045 = bht_rd_addr_hashed_p1_f == 8'h20; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_23525 = _T_23045 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23780 = _T_23779 | _T_23525; // @[Mux.scala 27:72]
  wire  _T_23047 = bht_rd_addr_hashed_p1_f == 8'h21; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_23526 = _T_23047 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23781 = _T_23780 | _T_23526; // @[Mux.scala 27:72]
  wire  _T_23049 = bht_rd_addr_hashed_p1_f == 8'h22; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_23527 = _T_23049 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23782 = _T_23781 | _T_23527; // @[Mux.scala 27:72]
  wire  _T_23051 = bht_rd_addr_hashed_p1_f == 8'h23; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_23528 = _T_23051 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23783 = _T_23782 | _T_23528; // @[Mux.scala 27:72]
  wire  _T_23053 = bht_rd_addr_hashed_p1_f == 8'h24; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_23529 = _T_23053 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23784 = _T_23783 | _T_23529; // @[Mux.scala 27:72]
  wire  _T_23055 = bht_rd_addr_hashed_p1_f == 8'h25; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_23530 = _T_23055 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23785 = _T_23784 | _T_23530; // @[Mux.scala 27:72]
  wire  _T_23057 = bht_rd_addr_hashed_p1_f == 8'h26; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_23531 = _T_23057 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23786 = _T_23785 | _T_23531; // @[Mux.scala 27:72]
  wire  _T_23059 = bht_rd_addr_hashed_p1_f == 8'h27; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_23532 = _T_23059 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23787 = _T_23786 | _T_23532; // @[Mux.scala 27:72]
  wire  _T_23061 = bht_rd_addr_hashed_p1_f == 8'h28; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_23533 = _T_23061 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23788 = _T_23787 | _T_23533; // @[Mux.scala 27:72]
  wire  _T_23063 = bht_rd_addr_hashed_p1_f == 8'h29; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_23534 = _T_23063 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23789 = _T_23788 | _T_23534; // @[Mux.scala 27:72]
  wire  _T_23065 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_23535 = _T_23065 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23790 = _T_23789 | _T_23535; // @[Mux.scala 27:72]
  wire  _T_23067 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_23536 = _T_23067 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23791 = _T_23790 | _T_23536; // @[Mux.scala 27:72]
  wire  _T_23069 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_23537 = _T_23069 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23792 = _T_23791 | _T_23537; // @[Mux.scala 27:72]
  wire  _T_23071 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_23538 = _T_23071 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23793 = _T_23792 | _T_23538; // @[Mux.scala 27:72]
  wire  _T_23073 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_23539 = _T_23073 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23794 = _T_23793 | _T_23539; // @[Mux.scala 27:72]
  wire  _T_23075 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_23540 = _T_23075 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23795 = _T_23794 | _T_23540; // @[Mux.scala 27:72]
  wire  _T_23077 = bht_rd_addr_hashed_p1_f == 8'h30; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_23541 = _T_23077 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23796 = _T_23795 | _T_23541; // @[Mux.scala 27:72]
  wire  _T_23079 = bht_rd_addr_hashed_p1_f == 8'h31; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_23542 = _T_23079 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23797 = _T_23796 | _T_23542; // @[Mux.scala 27:72]
  wire  _T_23081 = bht_rd_addr_hashed_p1_f == 8'h32; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_23543 = _T_23081 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23798 = _T_23797 | _T_23543; // @[Mux.scala 27:72]
  wire  _T_23083 = bht_rd_addr_hashed_p1_f == 8'h33; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_23544 = _T_23083 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23799 = _T_23798 | _T_23544; // @[Mux.scala 27:72]
  wire  _T_23085 = bht_rd_addr_hashed_p1_f == 8'h34; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_23545 = _T_23085 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23800 = _T_23799 | _T_23545; // @[Mux.scala 27:72]
  wire  _T_23087 = bht_rd_addr_hashed_p1_f == 8'h35; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_23546 = _T_23087 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23801 = _T_23800 | _T_23546; // @[Mux.scala 27:72]
  wire  _T_23089 = bht_rd_addr_hashed_p1_f == 8'h36; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_23547 = _T_23089 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23802 = _T_23801 | _T_23547; // @[Mux.scala 27:72]
  wire  _T_23091 = bht_rd_addr_hashed_p1_f == 8'h37; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_23548 = _T_23091 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23803 = _T_23802 | _T_23548; // @[Mux.scala 27:72]
  wire  _T_23093 = bht_rd_addr_hashed_p1_f == 8'h38; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_23549 = _T_23093 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23804 = _T_23803 | _T_23549; // @[Mux.scala 27:72]
  wire  _T_23095 = bht_rd_addr_hashed_p1_f == 8'h39; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_23550 = _T_23095 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23805 = _T_23804 | _T_23550; // @[Mux.scala 27:72]
  wire  _T_23097 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_23551 = _T_23097 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23806 = _T_23805 | _T_23551; // @[Mux.scala 27:72]
  wire  _T_23099 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_23552 = _T_23099 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23807 = _T_23806 | _T_23552; // @[Mux.scala 27:72]
  wire  _T_23101 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_23553 = _T_23101 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23808 = _T_23807 | _T_23553; // @[Mux.scala 27:72]
  wire  _T_23103 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_23554 = _T_23103 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23809 = _T_23808 | _T_23554; // @[Mux.scala 27:72]
  wire  _T_23105 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_23555 = _T_23105 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23810 = _T_23809 | _T_23555; // @[Mux.scala 27:72]
  wire  _T_23107 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_23556 = _T_23107 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23811 = _T_23810 | _T_23556; // @[Mux.scala 27:72]
  wire  _T_23109 = bht_rd_addr_hashed_p1_f == 8'h40; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_23557 = _T_23109 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23812 = _T_23811 | _T_23557; // @[Mux.scala 27:72]
  wire  _T_23111 = bht_rd_addr_hashed_p1_f == 8'h41; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_23558 = _T_23111 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23813 = _T_23812 | _T_23558; // @[Mux.scala 27:72]
  wire  _T_23113 = bht_rd_addr_hashed_p1_f == 8'h42; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_23559 = _T_23113 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23814 = _T_23813 | _T_23559; // @[Mux.scala 27:72]
  wire  _T_23115 = bht_rd_addr_hashed_p1_f == 8'h43; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_23560 = _T_23115 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23815 = _T_23814 | _T_23560; // @[Mux.scala 27:72]
  wire  _T_23117 = bht_rd_addr_hashed_p1_f == 8'h44; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_23561 = _T_23117 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23816 = _T_23815 | _T_23561; // @[Mux.scala 27:72]
  wire  _T_23119 = bht_rd_addr_hashed_p1_f == 8'h45; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_23562 = _T_23119 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23817 = _T_23816 | _T_23562; // @[Mux.scala 27:72]
  wire  _T_23121 = bht_rd_addr_hashed_p1_f == 8'h46; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_23563 = _T_23121 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23818 = _T_23817 | _T_23563; // @[Mux.scala 27:72]
  wire  _T_23123 = bht_rd_addr_hashed_p1_f == 8'h47; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_23564 = _T_23123 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23819 = _T_23818 | _T_23564; // @[Mux.scala 27:72]
  wire  _T_23125 = bht_rd_addr_hashed_p1_f == 8'h48; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_23565 = _T_23125 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23820 = _T_23819 | _T_23565; // @[Mux.scala 27:72]
  wire  _T_23127 = bht_rd_addr_hashed_p1_f == 8'h49; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_23566 = _T_23127 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23821 = _T_23820 | _T_23566; // @[Mux.scala 27:72]
  wire  _T_23129 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_23567 = _T_23129 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23822 = _T_23821 | _T_23567; // @[Mux.scala 27:72]
  wire  _T_23131 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_23568 = _T_23131 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23823 = _T_23822 | _T_23568; // @[Mux.scala 27:72]
  wire  _T_23133 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_23569 = _T_23133 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23824 = _T_23823 | _T_23569; // @[Mux.scala 27:72]
  wire  _T_23135 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_23570 = _T_23135 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23825 = _T_23824 | _T_23570; // @[Mux.scala 27:72]
  wire  _T_23137 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_23571 = _T_23137 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23826 = _T_23825 | _T_23571; // @[Mux.scala 27:72]
  wire  _T_23139 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_23572 = _T_23139 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23827 = _T_23826 | _T_23572; // @[Mux.scala 27:72]
  wire  _T_23141 = bht_rd_addr_hashed_p1_f == 8'h50; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_23573 = _T_23141 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23828 = _T_23827 | _T_23573; // @[Mux.scala 27:72]
  wire  _T_23143 = bht_rd_addr_hashed_p1_f == 8'h51; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_23574 = _T_23143 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23829 = _T_23828 | _T_23574; // @[Mux.scala 27:72]
  wire  _T_23145 = bht_rd_addr_hashed_p1_f == 8'h52; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_23575 = _T_23145 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23830 = _T_23829 | _T_23575; // @[Mux.scala 27:72]
  wire  _T_23147 = bht_rd_addr_hashed_p1_f == 8'h53; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_23576 = _T_23147 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23831 = _T_23830 | _T_23576; // @[Mux.scala 27:72]
  wire  _T_23149 = bht_rd_addr_hashed_p1_f == 8'h54; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_23577 = _T_23149 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23832 = _T_23831 | _T_23577; // @[Mux.scala 27:72]
  wire  _T_23151 = bht_rd_addr_hashed_p1_f == 8'h55; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_23578 = _T_23151 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23833 = _T_23832 | _T_23578; // @[Mux.scala 27:72]
  wire  _T_23153 = bht_rd_addr_hashed_p1_f == 8'h56; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_23579 = _T_23153 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23834 = _T_23833 | _T_23579; // @[Mux.scala 27:72]
  wire  _T_23155 = bht_rd_addr_hashed_p1_f == 8'h57; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_23580 = _T_23155 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23835 = _T_23834 | _T_23580; // @[Mux.scala 27:72]
  wire  _T_23157 = bht_rd_addr_hashed_p1_f == 8'h58; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_23581 = _T_23157 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23836 = _T_23835 | _T_23581; // @[Mux.scala 27:72]
  wire  _T_23159 = bht_rd_addr_hashed_p1_f == 8'h59; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_23582 = _T_23159 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23837 = _T_23836 | _T_23582; // @[Mux.scala 27:72]
  wire  _T_23161 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_23583 = _T_23161 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23838 = _T_23837 | _T_23583; // @[Mux.scala 27:72]
  wire  _T_23163 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_23584 = _T_23163 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23839 = _T_23838 | _T_23584; // @[Mux.scala 27:72]
  wire  _T_23165 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_23585 = _T_23165 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23840 = _T_23839 | _T_23585; // @[Mux.scala 27:72]
  wire  _T_23167 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_23586 = _T_23167 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23841 = _T_23840 | _T_23586; // @[Mux.scala 27:72]
  wire  _T_23169 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_23587 = _T_23169 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23842 = _T_23841 | _T_23587; // @[Mux.scala 27:72]
  wire  _T_23171 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_23588 = _T_23171 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23843 = _T_23842 | _T_23588; // @[Mux.scala 27:72]
  wire  _T_23173 = bht_rd_addr_hashed_p1_f == 8'h60; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_23589 = _T_23173 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23844 = _T_23843 | _T_23589; // @[Mux.scala 27:72]
  wire  _T_23175 = bht_rd_addr_hashed_p1_f == 8'h61; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_23590 = _T_23175 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23845 = _T_23844 | _T_23590; // @[Mux.scala 27:72]
  wire  _T_23177 = bht_rd_addr_hashed_p1_f == 8'h62; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_23591 = _T_23177 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23846 = _T_23845 | _T_23591; // @[Mux.scala 27:72]
  wire  _T_23179 = bht_rd_addr_hashed_p1_f == 8'h63; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_23592 = _T_23179 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23847 = _T_23846 | _T_23592; // @[Mux.scala 27:72]
  wire  _T_23181 = bht_rd_addr_hashed_p1_f == 8'h64; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_23593 = _T_23181 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23848 = _T_23847 | _T_23593; // @[Mux.scala 27:72]
  wire  _T_23183 = bht_rd_addr_hashed_p1_f == 8'h65; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_23594 = _T_23183 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23849 = _T_23848 | _T_23594; // @[Mux.scala 27:72]
  wire  _T_23185 = bht_rd_addr_hashed_p1_f == 8'h66; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_23595 = _T_23185 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23850 = _T_23849 | _T_23595; // @[Mux.scala 27:72]
  wire  _T_23187 = bht_rd_addr_hashed_p1_f == 8'h67; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_23596 = _T_23187 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23851 = _T_23850 | _T_23596; // @[Mux.scala 27:72]
  wire  _T_23189 = bht_rd_addr_hashed_p1_f == 8'h68; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_23597 = _T_23189 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23852 = _T_23851 | _T_23597; // @[Mux.scala 27:72]
  wire  _T_23191 = bht_rd_addr_hashed_p1_f == 8'h69; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_23598 = _T_23191 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23853 = _T_23852 | _T_23598; // @[Mux.scala 27:72]
  wire  _T_23193 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_23599 = _T_23193 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23854 = _T_23853 | _T_23599; // @[Mux.scala 27:72]
  wire  _T_23195 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_23600 = _T_23195 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23855 = _T_23854 | _T_23600; // @[Mux.scala 27:72]
  wire  _T_23197 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_23601 = _T_23197 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23856 = _T_23855 | _T_23601; // @[Mux.scala 27:72]
  wire  _T_23199 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_23602 = _T_23199 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23857 = _T_23856 | _T_23602; // @[Mux.scala 27:72]
  wire  _T_23201 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_23603 = _T_23201 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23858 = _T_23857 | _T_23603; // @[Mux.scala 27:72]
  wire  _T_23203 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_23604 = _T_23203 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23859 = _T_23858 | _T_23604; // @[Mux.scala 27:72]
  wire  _T_23205 = bht_rd_addr_hashed_p1_f == 8'h70; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_23605 = _T_23205 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23860 = _T_23859 | _T_23605; // @[Mux.scala 27:72]
  wire  _T_23207 = bht_rd_addr_hashed_p1_f == 8'h71; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_23606 = _T_23207 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23861 = _T_23860 | _T_23606; // @[Mux.scala 27:72]
  wire  _T_23209 = bht_rd_addr_hashed_p1_f == 8'h72; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_23607 = _T_23209 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23862 = _T_23861 | _T_23607; // @[Mux.scala 27:72]
  wire  _T_23211 = bht_rd_addr_hashed_p1_f == 8'h73; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_23608 = _T_23211 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23863 = _T_23862 | _T_23608; // @[Mux.scala 27:72]
  wire  _T_23213 = bht_rd_addr_hashed_p1_f == 8'h74; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_23609 = _T_23213 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23864 = _T_23863 | _T_23609; // @[Mux.scala 27:72]
  wire  _T_23215 = bht_rd_addr_hashed_p1_f == 8'h75; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_23610 = _T_23215 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23865 = _T_23864 | _T_23610; // @[Mux.scala 27:72]
  wire  _T_23217 = bht_rd_addr_hashed_p1_f == 8'h76; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_23611 = _T_23217 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23866 = _T_23865 | _T_23611; // @[Mux.scala 27:72]
  wire  _T_23219 = bht_rd_addr_hashed_p1_f == 8'h77; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_23612 = _T_23219 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23867 = _T_23866 | _T_23612; // @[Mux.scala 27:72]
  wire  _T_23221 = bht_rd_addr_hashed_p1_f == 8'h78; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_23613 = _T_23221 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23868 = _T_23867 | _T_23613; // @[Mux.scala 27:72]
  wire  _T_23223 = bht_rd_addr_hashed_p1_f == 8'h79; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_23614 = _T_23223 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23869 = _T_23868 | _T_23614; // @[Mux.scala 27:72]
  wire  _T_23225 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_23615 = _T_23225 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23870 = _T_23869 | _T_23615; // @[Mux.scala 27:72]
  wire  _T_23227 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_23616 = _T_23227 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23871 = _T_23870 | _T_23616; // @[Mux.scala 27:72]
  wire  _T_23229 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_23617 = _T_23229 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23872 = _T_23871 | _T_23617; // @[Mux.scala 27:72]
  wire  _T_23231 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_23618 = _T_23231 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23873 = _T_23872 | _T_23618; // @[Mux.scala 27:72]
  wire  _T_23233 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_23619 = _T_23233 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23874 = _T_23873 | _T_23619; // @[Mux.scala 27:72]
  wire  _T_23235 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_23620 = _T_23235 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23875 = _T_23874 | _T_23620; // @[Mux.scala 27:72]
  wire  _T_23237 = bht_rd_addr_hashed_p1_f == 8'h80; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_23621 = _T_23237 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23876 = _T_23875 | _T_23621; // @[Mux.scala 27:72]
  wire  _T_23239 = bht_rd_addr_hashed_p1_f == 8'h81; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_23622 = _T_23239 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23877 = _T_23876 | _T_23622; // @[Mux.scala 27:72]
  wire  _T_23241 = bht_rd_addr_hashed_p1_f == 8'h82; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_23623 = _T_23241 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23878 = _T_23877 | _T_23623; // @[Mux.scala 27:72]
  wire  _T_23243 = bht_rd_addr_hashed_p1_f == 8'h83; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_23624 = _T_23243 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23879 = _T_23878 | _T_23624; // @[Mux.scala 27:72]
  wire  _T_23245 = bht_rd_addr_hashed_p1_f == 8'h84; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_23625 = _T_23245 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23880 = _T_23879 | _T_23625; // @[Mux.scala 27:72]
  wire  _T_23247 = bht_rd_addr_hashed_p1_f == 8'h85; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_23626 = _T_23247 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23881 = _T_23880 | _T_23626; // @[Mux.scala 27:72]
  wire  _T_23249 = bht_rd_addr_hashed_p1_f == 8'h86; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_23627 = _T_23249 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23882 = _T_23881 | _T_23627; // @[Mux.scala 27:72]
  wire  _T_23251 = bht_rd_addr_hashed_p1_f == 8'h87; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_23628 = _T_23251 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23883 = _T_23882 | _T_23628; // @[Mux.scala 27:72]
  wire  _T_23253 = bht_rd_addr_hashed_p1_f == 8'h88; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_23629 = _T_23253 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23884 = _T_23883 | _T_23629; // @[Mux.scala 27:72]
  wire  _T_23255 = bht_rd_addr_hashed_p1_f == 8'h89; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_23630 = _T_23255 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23885 = _T_23884 | _T_23630; // @[Mux.scala 27:72]
  wire  _T_23257 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_23631 = _T_23257 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23886 = _T_23885 | _T_23631; // @[Mux.scala 27:72]
  wire  _T_23259 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_23632 = _T_23259 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23887 = _T_23886 | _T_23632; // @[Mux.scala 27:72]
  wire  _T_23261 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_23633 = _T_23261 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23888 = _T_23887 | _T_23633; // @[Mux.scala 27:72]
  wire  _T_23263 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_23634 = _T_23263 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23889 = _T_23888 | _T_23634; // @[Mux.scala 27:72]
  wire  _T_23265 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_23635 = _T_23265 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23890 = _T_23889 | _T_23635; // @[Mux.scala 27:72]
  wire  _T_23267 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_23636 = _T_23267 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23891 = _T_23890 | _T_23636; // @[Mux.scala 27:72]
  wire  _T_23269 = bht_rd_addr_hashed_p1_f == 8'h90; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_23637 = _T_23269 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23892 = _T_23891 | _T_23637; // @[Mux.scala 27:72]
  wire  _T_23271 = bht_rd_addr_hashed_p1_f == 8'h91; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_23638 = _T_23271 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23893 = _T_23892 | _T_23638; // @[Mux.scala 27:72]
  wire  _T_23273 = bht_rd_addr_hashed_p1_f == 8'h92; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_23639 = _T_23273 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23894 = _T_23893 | _T_23639; // @[Mux.scala 27:72]
  wire  _T_23275 = bht_rd_addr_hashed_p1_f == 8'h93; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_23640 = _T_23275 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23895 = _T_23894 | _T_23640; // @[Mux.scala 27:72]
  wire  _T_23277 = bht_rd_addr_hashed_p1_f == 8'h94; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_23641 = _T_23277 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23896 = _T_23895 | _T_23641; // @[Mux.scala 27:72]
  wire  _T_23279 = bht_rd_addr_hashed_p1_f == 8'h95; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_23642 = _T_23279 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23897 = _T_23896 | _T_23642; // @[Mux.scala 27:72]
  wire  _T_23281 = bht_rd_addr_hashed_p1_f == 8'h96; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_23643 = _T_23281 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23898 = _T_23897 | _T_23643; // @[Mux.scala 27:72]
  wire  _T_23283 = bht_rd_addr_hashed_p1_f == 8'h97; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_23644 = _T_23283 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23899 = _T_23898 | _T_23644; // @[Mux.scala 27:72]
  wire  _T_23285 = bht_rd_addr_hashed_p1_f == 8'h98; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_23645 = _T_23285 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23900 = _T_23899 | _T_23645; // @[Mux.scala 27:72]
  wire  _T_23287 = bht_rd_addr_hashed_p1_f == 8'h99; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_23646 = _T_23287 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23901 = _T_23900 | _T_23646; // @[Mux.scala 27:72]
  wire  _T_23289 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_23647 = _T_23289 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23902 = _T_23901 | _T_23647; // @[Mux.scala 27:72]
  wire  _T_23291 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_23648 = _T_23291 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23903 = _T_23902 | _T_23648; // @[Mux.scala 27:72]
  wire  _T_23293 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_23649 = _T_23293 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23904 = _T_23903 | _T_23649; // @[Mux.scala 27:72]
  wire  _T_23295 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_23650 = _T_23295 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23905 = _T_23904 | _T_23650; // @[Mux.scala 27:72]
  wire  _T_23297 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_23651 = _T_23297 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23906 = _T_23905 | _T_23651; // @[Mux.scala 27:72]
  wire  _T_23299 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_23652 = _T_23299 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23907 = _T_23906 | _T_23652; // @[Mux.scala 27:72]
  wire  _T_23301 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_23653 = _T_23301 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23908 = _T_23907 | _T_23653; // @[Mux.scala 27:72]
  wire  _T_23303 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_23654 = _T_23303 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23909 = _T_23908 | _T_23654; // @[Mux.scala 27:72]
  wire  _T_23305 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_23655 = _T_23305 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23910 = _T_23909 | _T_23655; // @[Mux.scala 27:72]
  wire  _T_23307 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_23656 = _T_23307 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23911 = _T_23910 | _T_23656; // @[Mux.scala 27:72]
  wire  _T_23309 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_23657 = _T_23309 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23912 = _T_23911 | _T_23657; // @[Mux.scala 27:72]
  wire  _T_23311 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_23658 = _T_23311 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23913 = _T_23912 | _T_23658; // @[Mux.scala 27:72]
  wire  _T_23313 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_23659 = _T_23313 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23914 = _T_23913 | _T_23659; // @[Mux.scala 27:72]
  wire  _T_23315 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_23660 = _T_23315 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23915 = _T_23914 | _T_23660; // @[Mux.scala 27:72]
  wire  _T_23317 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_23661 = _T_23317 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23916 = _T_23915 | _T_23661; // @[Mux.scala 27:72]
  wire  _T_23319 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_23662 = _T_23319 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23917 = _T_23916 | _T_23662; // @[Mux.scala 27:72]
  wire  _T_23321 = bht_rd_addr_hashed_p1_f == 8'haa; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_23663 = _T_23321 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23918 = _T_23917 | _T_23663; // @[Mux.scala 27:72]
  wire  _T_23323 = bht_rd_addr_hashed_p1_f == 8'hab; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_23664 = _T_23323 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23919 = _T_23918 | _T_23664; // @[Mux.scala 27:72]
  wire  _T_23325 = bht_rd_addr_hashed_p1_f == 8'hac; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_23665 = _T_23325 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23920 = _T_23919 | _T_23665; // @[Mux.scala 27:72]
  wire  _T_23327 = bht_rd_addr_hashed_p1_f == 8'had; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_23666 = _T_23327 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23921 = _T_23920 | _T_23666; // @[Mux.scala 27:72]
  wire  _T_23329 = bht_rd_addr_hashed_p1_f == 8'hae; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_23667 = _T_23329 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23922 = _T_23921 | _T_23667; // @[Mux.scala 27:72]
  wire  _T_23331 = bht_rd_addr_hashed_p1_f == 8'haf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_23668 = _T_23331 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23923 = _T_23922 | _T_23668; // @[Mux.scala 27:72]
  wire  _T_23333 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_23669 = _T_23333 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23924 = _T_23923 | _T_23669; // @[Mux.scala 27:72]
  wire  _T_23335 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_23670 = _T_23335 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23925 = _T_23924 | _T_23670; // @[Mux.scala 27:72]
  wire  _T_23337 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_23671 = _T_23337 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23926 = _T_23925 | _T_23671; // @[Mux.scala 27:72]
  wire  _T_23339 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_23672 = _T_23339 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23927 = _T_23926 | _T_23672; // @[Mux.scala 27:72]
  wire  _T_23341 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_23673 = _T_23341 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23928 = _T_23927 | _T_23673; // @[Mux.scala 27:72]
  wire  _T_23343 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_23674 = _T_23343 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23929 = _T_23928 | _T_23674; // @[Mux.scala 27:72]
  wire  _T_23345 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_23675 = _T_23345 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23930 = _T_23929 | _T_23675; // @[Mux.scala 27:72]
  wire  _T_23347 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_23676 = _T_23347 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23931 = _T_23930 | _T_23676; // @[Mux.scala 27:72]
  wire  _T_23349 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_23677 = _T_23349 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23932 = _T_23931 | _T_23677; // @[Mux.scala 27:72]
  wire  _T_23351 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_23678 = _T_23351 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23933 = _T_23932 | _T_23678; // @[Mux.scala 27:72]
  wire  _T_23353 = bht_rd_addr_hashed_p1_f == 8'hba; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_23679 = _T_23353 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23934 = _T_23933 | _T_23679; // @[Mux.scala 27:72]
  wire  _T_23355 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_23680 = _T_23355 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23935 = _T_23934 | _T_23680; // @[Mux.scala 27:72]
  wire  _T_23357 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_23681 = _T_23357 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23936 = _T_23935 | _T_23681; // @[Mux.scala 27:72]
  wire  _T_23359 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_23682 = _T_23359 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23937 = _T_23936 | _T_23682; // @[Mux.scala 27:72]
  wire  _T_23361 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_23683 = _T_23361 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23938 = _T_23937 | _T_23683; // @[Mux.scala 27:72]
  wire  _T_23363 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_23684 = _T_23363 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23939 = _T_23938 | _T_23684; // @[Mux.scala 27:72]
  wire  _T_23365 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_23685 = _T_23365 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23940 = _T_23939 | _T_23685; // @[Mux.scala 27:72]
  wire  _T_23367 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_23686 = _T_23367 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23941 = _T_23940 | _T_23686; // @[Mux.scala 27:72]
  wire  _T_23369 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_23687 = _T_23369 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23942 = _T_23941 | _T_23687; // @[Mux.scala 27:72]
  wire  _T_23371 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_23688 = _T_23371 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23943 = _T_23942 | _T_23688; // @[Mux.scala 27:72]
  wire  _T_23373 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_23689 = _T_23373 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23944 = _T_23943 | _T_23689; // @[Mux.scala 27:72]
  wire  _T_23375 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_23690 = _T_23375 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23945 = _T_23944 | _T_23690; // @[Mux.scala 27:72]
  wire  _T_23377 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_23691 = _T_23377 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23946 = _T_23945 | _T_23691; // @[Mux.scala 27:72]
  wire  _T_23379 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_23692 = _T_23379 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23947 = _T_23946 | _T_23692; // @[Mux.scala 27:72]
  wire  _T_23381 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_23693 = _T_23381 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23948 = _T_23947 | _T_23693; // @[Mux.scala 27:72]
  wire  _T_23383 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_23694 = _T_23383 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23949 = _T_23948 | _T_23694; // @[Mux.scala 27:72]
  wire  _T_23385 = bht_rd_addr_hashed_p1_f == 8'hca; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_23695 = _T_23385 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23950 = _T_23949 | _T_23695; // @[Mux.scala 27:72]
  wire  _T_23387 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_23696 = _T_23387 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23951 = _T_23950 | _T_23696; // @[Mux.scala 27:72]
  wire  _T_23389 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_23697 = _T_23389 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23952 = _T_23951 | _T_23697; // @[Mux.scala 27:72]
  wire  _T_23391 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_23698 = _T_23391 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23953 = _T_23952 | _T_23698; // @[Mux.scala 27:72]
  wire  _T_23393 = bht_rd_addr_hashed_p1_f == 8'hce; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_23699 = _T_23393 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23954 = _T_23953 | _T_23699; // @[Mux.scala 27:72]
  wire  _T_23395 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_23700 = _T_23395 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23955 = _T_23954 | _T_23700; // @[Mux.scala 27:72]
  wire  _T_23397 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_23701 = _T_23397 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23956 = _T_23955 | _T_23701; // @[Mux.scala 27:72]
  wire  _T_23399 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_23702 = _T_23399 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23957 = _T_23956 | _T_23702; // @[Mux.scala 27:72]
  wire  _T_23401 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_23703 = _T_23401 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23958 = _T_23957 | _T_23703; // @[Mux.scala 27:72]
  wire  _T_23403 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_23704 = _T_23403 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23959 = _T_23958 | _T_23704; // @[Mux.scala 27:72]
  wire  _T_23405 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_23705 = _T_23405 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23960 = _T_23959 | _T_23705; // @[Mux.scala 27:72]
  wire  _T_23407 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_23706 = _T_23407 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23961 = _T_23960 | _T_23706; // @[Mux.scala 27:72]
  wire  _T_23409 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_23707 = _T_23409 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23962 = _T_23961 | _T_23707; // @[Mux.scala 27:72]
  wire  _T_23411 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_23708 = _T_23411 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23963 = _T_23962 | _T_23708; // @[Mux.scala 27:72]
  wire  _T_23413 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_23709 = _T_23413 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23964 = _T_23963 | _T_23709; // @[Mux.scala 27:72]
  wire  _T_23415 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_23710 = _T_23415 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23965 = _T_23964 | _T_23710; // @[Mux.scala 27:72]
  wire  _T_23417 = bht_rd_addr_hashed_p1_f == 8'hda; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_23711 = _T_23417 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23966 = _T_23965 | _T_23711; // @[Mux.scala 27:72]
  wire  _T_23419 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_23712 = _T_23419 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23967 = _T_23966 | _T_23712; // @[Mux.scala 27:72]
  wire  _T_23421 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_23713 = _T_23421 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23968 = _T_23967 | _T_23713; // @[Mux.scala 27:72]
  wire  _T_23423 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_23714 = _T_23423 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23969 = _T_23968 | _T_23714; // @[Mux.scala 27:72]
  wire  _T_23425 = bht_rd_addr_hashed_p1_f == 8'hde; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_23715 = _T_23425 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23970 = _T_23969 | _T_23715; // @[Mux.scala 27:72]
  wire  _T_23427 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_23716 = _T_23427 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23971 = _T_23970 | _T_23716; // @[Mux.scala 27:72]
  wire  _T_23429 = bht_rd_addr_hashed_p1_f == 8'he0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_23717 = _T_23429 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23972 = _T_23971 | _T_23717; // @[Mux.scala 27:72]
  wire  _T_23431 = bht_rd_addr_hashed_p1_f == 8'he1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_23718 = _T_23431 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23973 = _T_23972 | _T_23718; // @[Mux.scala 27:72]
  wire  _T_23433 = bht_rd_addr_hashed_p1_f == 8'he2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_23719 = _T_23433 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23974 = _T_23973 | _T_23719; // @[Mux.scala 27:72]
  wire  _T_23435 = bht_rd_addr_hashed_p1_f == 8'he3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_23720 = _T_23435 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23975 = _T_23974 | _T_23720; // @[Mux.scala 27:72]
  wire  _T_23437 = bht_rd_addr_hashed_p1_f == 8'he4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_23721 = _T_23437 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23976 = _T_23975 | _T_23721; // @[Mux.scala 27:72]
  wire  _T_23439 = bht_rd_addr_hashed_p1_f == 8'he5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_23722 = _T_23439 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23977 = _T_23976 | _T_23722; // @[Mux.scala 27:72]
  wire  _T_23441 = bht_rd_addr_hashed_p1_f == 8'he6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_23723 = _T_23441 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23978 = _T_23977 | _T_23723; // @[Mux.scala 27:72]
  wire  _T_23443 = bht_rd_addr_hashed_p1_f == 8'he7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_23724 = _T_23443 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23979 = _T_23978 | _T_23724; // @[Mux.scala 27:72]
  wire  _T_23445 = bht_rd_addr_hashed_p1_f == 8'he8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_23725 = _T_23445 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23980 = _T_23979 | _T_23725; // @[Mux.scala 27:72]
  wire  _T_23447 = bht_rd_addr_hashed_p1_f == 8'he9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_23726 = _T_23447 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23981 = _T_23980 | _T_23726; // @[Mux.scala 27:72]
  wire  _T_23449 = bht_rd_addr_hashed_p1_f == 8'hea; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_23727 = _T_23449 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23982 = _T_23981 | _T_23727; // @[Mux.scala 27:72]
  wire  _T_23451 = bht_rd_addr_hashed_p1_f == 8'heb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_23728 = _T_23451 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23983 = _T_23982 | _T_23728; // @[Mux.scala 27:72]
  wire  _T_23453 = bht_rd_addr_hashed_p1_f == 8'hec; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_23729 = _T_23453 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23984 = _T_23983 | _T_23729; // @[Mux.scala 27:72]
  wire  _T_23455 = bht_rd_addr_hashed_p1_f == 8'hed; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_23730 = _T_23455 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23985 = _T_23984 | _T_23730; // @[Mux.scala 27:72]
  wire  _T_23457 = bht_rd_addr_hashed_p1_f == 8'hee; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_23731 = _T_23457 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23986 = _T_23985 | _T_23731; // @[Mux.scala 27:72]
  wire  _T_23459 = bht_rd_addr_hashed_p1_f == 8'hef; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_23732 = _T_23459 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23987 = _T_23986 | _T_23732; // @[Mux.scala 27:72]
  wire  _T_23461 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_23733 = _T_23461 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23988 = _T_23987 | _T_23733; // @[Mux.scala 27:72]
  wire  _T_23463 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_23734 = _T_23463 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23989 = _T_23988 | _T_23734; // @[Mux.scala 27:72]
  wire  _T_23465 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_23735 = _T_23465 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23990 = _T_23989 | _T_23735; // @[Mux.scala 27:72]
  wire  _T_23467 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_23736 = _T_23467 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23991 = _T_23990 | _T_23736; // @[Mux.scala 27:72]
  wire  _T_23469 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_23737 = _T_23469 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23992 = _T_23991 | _T_23737; // @[Mux.scala 27:72]
  wire  _T_23471 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_23738 = _T_23471 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23993 = _T_23992 | _T_23738; // @[Mux.scala 27:72]
  wire  _T_23473 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_23739 = _T_23473 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23994 = _T_23993 | _T_23739; // @[Mux.scala 27:72]
  wire  _T_23475 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_23740 = _T_23475 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23995 = _T_23994 | _T_23740; // @[Mux.scala 27:72]
  wire  _T_23477 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_23741 = _T_23477 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23996 = _T_23995 | _T_23741; // @[Mux.scala 27:72]
  wire  _T_23479 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_23742 = _T_23479 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23997 = _T_23996 | _T_23742; // @[Mux.scala 27:72]
  wire  _T_23481 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_23743 = _T_23481 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23998 = _T_23997 | _T_23743; // @[Mux.scala 27:72]
  wire  _T_23483 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_23744 = _T_23483 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23999 = _T_23998 | _T_23744; // @[Mux.scala 27:72]
  wire  _T_23485 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_23745 = _T_23485 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24000 = _T_23999 | _T_23745; // @[Mux.scala 27:72]
  wire  _T_23487 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_23746 = _T_23487 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24001 = _T_24000 | _T_23746; // @[Mux.scala 27:72]
  wire  _T_23489 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_23747 = _T_23489 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24002 = _T_24001 | _T_23747; // @[Mux.scala 27:72]
  wire  _T_23491 = bht_rd_addr_hashed_p1_f == 8'hff; // @[ifu_bp_ctl.scala 537:85]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_23748 = _T_23491 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_24002 | _T_23748; // @[Mux.scala 27:72]
  wire [1:0] _T_254 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_253 | _T_254; // @[Mux.scala 27:72]
  wire  _T_258 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 298:42]
  wire [1:0] wayhit_f = tag_match_way0_expanded_f | tag_match_way1_expanded_f; // @[ifu_bp_ctl.scala 172:41]
  wire [1:0] _T_607 = _T_147 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = tag_match_way0_expanded_p1_f | tag_match_way1_expanded_p1_f; // @[ifu_bp_ctl.scala 174:47]
  wire [1:0] _T_606 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_608 = io_ifc_fetch_addr_f[0] ? _T_606 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_609 = _T_607 | _T_608; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[ifu_bp_ctl.scala 258:64]
  wire  _T_212 = ~eoc_near; // @[ifu_bp_ctl.scala 260:15]
  wire [1:0] _T_214 = ~io_ifc_fetch_addr_f[1:0]; // @[ifu_bp_ctl.scala 260:28]
  wire  _T_215 = |_T_214; // @[ifu_bp_ctl.scala 260:58]
  wire  eoc_mask = _T_212 | _T_215; // @[ifu_bp_ctl.scala 260:25]
  wire [1:0] _T_611 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] vwayhit_f = _T_609 & _T_611; // @[ifu_bp_ctl.scala 431:71]
  wire  _T_260 = _T_258 & vwayhit_f[1]; // @[ifu_bp_ctl.scala 298:69]
  wire [1:0] _T_21445 = _T_21957 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21446 = _T_21959 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21701 = _T_21445 | _T_21446; // @[Mux.scala 27:72]
  wire [1:0] _T_21447 = _T_21961 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21702 = _T_21701 | _T_21447; // @[Mux.scala 27:72]
  wire [1:0] _T_21448 = _T_21963 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21703 = _T_21702 | _T_21448; // @[Mux.scala 27:72]
  wire [1:0] _T_21449 = _T_21965 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21704 = _T_21703 | _T_21449; // @[Mux.scala 27:72]
  wire [1:0] _T_21450 = _T_21967 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21705 = _T_21704 | _T_21450; // @[Mux.scala 27:72]
  wire [1:0] _T_21451 = _T_21969 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21706 = _T_21705 | _T_21451; // @[Mux.scala 27:72]
  wire [1:0] _T_21452 = _T_21971 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21707 = _T_21706 | _T_21452; // @[Mux.scala 27:72]
  wire [1:0] _T_21453 = _T_21973 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21708 = _T_21707 | _T_21453; // @[Mux.scala 27:72]
  wire [1:0] _T_21454 = _T_21975 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21709 = _T_21708 | _T_21454; // @[Mux.scala 27:72]
  wire [1:0] _T_21455 = _T_21977 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21710 = _T_21709 | _T_21455; // @[Mux.scala 27:72]
  wire [1:0] _T_21456 = _T_21979 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21711 = _T_21710 | _T_21456; // @[Mux.scala 27:72]
  wire [1:0] _T_21457 = _T_21981 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21712 = _T_21711 | _T_21457; // @[Mux.scala 27:72]
  wire [1:0] _T_21458 = _T_21983 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21713 = _T_21712 | _T_21458; // @[Mux.scala 27:72]
  wire [1:0] _T_21459 = _T_21985 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21714 = _T_21713 | _T_21459; // @[Mux.scala 27:72]
  wire [1:0] _T_21460 = _T_21987 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21715 = _T_21714 | _T_21460; // @[Mux.scala 27:72]
  wire [1:0] _T_21461 = _T_21989 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21716 = _T_21715 | _T_21461; // @[Mux.scala 27:72]
  wire [1:0] _T_21462 = _T_21991 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21717 = _T_21716 | _T_21462; // @[Mux.scala 27:72]
  wire [1:0] _T_21463 = _T_21993 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21718 = _T_21717 | _T_21463; // @[Mux.scala 27:72]
  wire [1:0] _T_21464 = _T_21995 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21719 = _T_21718 | _T_21464; // @[Mux.scala 27:72]
  wire [1:0] _T_21465 = _T_21997 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21720 = _T_21719 | _T_21465; // @[Mux.scala 27:72]
  wire [1:0] _T_21466 = _T_21999 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21721 = _T_21720 | _T_21466; // @[Mux.scala 27:72]
  wire [1:0] _T_21467 = _T_22001 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21722 = _T_21721 | _T_21467; // @[Mux.scala 27:72]
  wire [1:0] _T_21468 = _T_22003 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21723 = _T_21722 | _T_21468; // @[Mux.scala 27:72]
  wire [1:0] _T_21469 = _T_22005 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21724 = _T_21723 | _T_21469; // @[Mux.scala 27:72]
  wire [1:0] _T_21470 = _T_22007 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21725 = _T_21724 | _T_21470; // @[Mux.scala 27:72]
  wire [1:0] _T_21471 = _T_22009 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21726 = _T_21725 | _T_21471; // @[Mux.scala 27:72]
  wire [1:0] _T_21472 = _T_22011 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21727 = _T_21726 | _T_21472; // @[Mux.scala 27:72]
  wire [1:0] _T_21473 = _T_22013 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21728 = _T_21727 | _T_21473; // @[Mux.scala 27:72]
  wire [1:0] _T_21474 = _T_22015 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21729 = _T_21728 | _T_21474; // @[Mux.scala 27:72]
  wire [1:0] _T_21475 = _T_22017 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21730 = _T_21729 | _T_21475; // @[Mux.scala 27:72]
  wire [1:0] _T_21476 = _T_22019 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21731 = _T_21730 | _T_21476; // @[Mux.scala 27:72]
  wire [1:0] _T_21477 = _T_22021 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21732 = _T_21731 | _T_21477; // @[Mux.scala 27:72]
  wire [1:0] _T_21478 = _T_22023 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21733 = _T_21732 | _T_21478; // @[Mux.scala 27:72]
  wire [1:0] _T_21479 = _T_22025 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21734 = _T_21733 | _T_21479; // @[Mux.scala 27:72]
  wire [1:0] _T_21480 = _T_22027 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21735 = _T_21734 | _T_21480; // @[Mux.scala 27:72]
  wire [1:0] _T_21481 = _T_22029 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21736 = _T_21735 | _T_21481; // @[Mux.scala 27:72]
  wire [1:0] _T_21482 = _T_22031 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21737 = _T_21736 | _T_21482; // @[Mux.scala 27:72]
  wire [1:0] _T_21483 = _T_22033 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21738 = _T_21737 | _T_21483; // @[Mux.scala 27:72]
  wire [1:0] _T_21484 = _T_22035 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21739 = _T_21738 | _T_21484; // @[Mux.scala 27:72]
  wire [1:0] _T_21485 = _T_22037 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21740 = _T_21739 | _T_21485; // @[Mux.scala 27:72]
  wire [1:0] _T_21486 = _T_22039 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21741 = _T_21740 | _T_21486; // @[Mux.scala 27:72]
  wire [1:0] _T_21487 = _T_22041 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21742 = _T_21741 | _T_21487; // @[Mux.scala 27:72]
  wire [1:0] _T_21488 = _T_22043 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21743 = _T_21742 | _T_21488; // @[Mux.scala 27:72]
  wire [1:0] _T_21489 = _T_22045 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21744 = _T_21743 | _T_21489; // @[Mux.scala 27:72]
  wire [1:0] _T_21490 = _T_22047 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21745 = _T_21744 | _T_21490; // @[Mux.scala 27:72]
  wire [1:0] _T_21491 = _T_22049 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21746 = _T_21745 | _T_21491; // @[Mux.scala 27:72]
  wire [1:0] _T_21492 = _T_22051 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21747 = _T_21746 | _T_21492; // @[Mux.scala 27:72]
  wire [1:0] _T_21493 = _T_22053 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21748 = _T_21747 | _T_21493; // @[Mux.scala 27:72]
  wire [1:0] _T_21494 = _T_22055 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21749 = _T_21748 | _T_21494; // @[Mux.scala 27:72]
  wire [1:0] _T_21495 = _T_22057 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21750 = _T_21749 | _T_21495; // @[Mux.scala 27:72]
  wire [1:0] _T_21496 = _T_22059 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21751 = _T_21750 | _T_21496; // @[Mux.scala 27:72]
  wire [1:0] _T_21497 = _T_22061 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21752 = _T_21751 | _T_21497; // @[Mux.scala 27:72]
  wire [1:0] _T_21498 = _T_22063 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21753 = _T_21752 | _T_21498; // @[Mux.scala 27:72]
  wire [1:0] _T_21499 = _T_22065 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21754 = _T_21753 | _T_21499; // @[Mux.scala 27:72]
  wire [1:0] _T_21500 = _T_22067 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21755 = _T_21754 | _T_21500; // @[Mux.scala 27:72]
  wire [1:0] _T_21501 = _T_22069 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21756 = _T_21755 | _T_21501; // @[Mux.scala 27:72]
  wire [1:0] _T_21502 = _T_22071 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21757 = _T_21756 | _T_21502; // @[Mux.scala 27:72]
  wire [1:0] _T_21503 = _T_22073 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21758 = _T_21757 | _T_21503; // @[Mux.scala 27:72]
  wire [1:0] _T_21504 = _T_22075 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21759 = _T_21758 | _T_21504; // @[Mux.scala 27:72]
  wire [1:0] _T_21505 = _T_22077 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21760 = _T_21759 | _T_21505; // @[Mux.scala 27:72]
  wire [1:0] _T_21506 = _T_22079 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21761 = _T_21760 | _T_21506; // @[Mux.scala 27:72]
  wire [1:0] _T_21507 = _T_22081 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21762 = _T_21761 | _T_21507; // @[Mux.scala 27:72]
  wire [1:0] _T_21508 = _T_22083 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21763 = _T_21762 | _T_21508; // @[Mux.scala 27:72]
  wire [1:0] _T_21509 = _T_22085 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21764 = _T_21763 | _T_21509; // @[Mux.scala 27:72]
  wire [1:0] _T_21510 = _T_22087 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21765 = _T_21764 | _T_21510; // @[Mux.scala 27:72]
  wire [1:0] _T_21511 = _T_22089 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21766 = _T_21765 | _T_21511; // @[Mux.scala 27:72]
  wire [1:0] _T_21512 = _T_22091 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21767 = _T_21766 | _T_21512; // @[Mux.scala 27:72]
  wire [1:0] _T_21513 = _T_22093 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21768 = _T_21767 | _T_21513; // @[Mux.scala 27:72]
  wire [1:0] _T_21514 = _T_22095 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21769 = _T_21768 | _T_21514; // @[Mux.scala 27:72]
  wire [1:0] _T_21515 = _T_22097 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21770 = _T_21769 | _T_21515; // @[Mux.scala 27:72]
  wire [1:0] _T_21516 = _T_22099 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21771 = _T_21770 | _T_21516; // @[Mux.scala 27:72]
  wire [1:0] _T_21517 = _T_22101 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21772 = _T_21771 | _T_21517; // @[Mux.scala 27:72]
  wire [1:0] _T_21518 = _T_22103 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21773 = _T_21772 | _T_21518; // @[Mux.scala 27:72]
  wire [1:0] _T_21519 = _T_22105 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21774 = _T_21773 | _T_21519; // @[Mux.scala 27:72]
  wire [1:0] _T_21520 = _T_22107 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21775 = _T_21774 | _T_21520; // @[Mux.scala 27:72]
  wire [1:0] _T_21521 = _T_22109 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21776 = _T_21775 | _T_21521; // @[Mux.scala 27:72]
  wire [1:0] _T_21522 = _T_22111 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21777 = _T_21776 | _T_21522; // @[Mux.scala 27:72]
  wire [1:0] _T_21523 = _T_22113 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21778 = _T_21777 | _T_21523; // @[Mux.scala 27:72]
  wire [1:0] _T_21524 = _T_22115 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21779 = _T_21778 | _T_21524; // @[Mux.scala 27:72]
  wire [1:0] _T_21525 = _T_22117 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21780 = _T_21779 | _T_21525; // @[Mux.scala 27:72]
  wire [1:0] _T_21526 = _T_22119 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21781 = _T_21780 | _T_21526; // @[Mux.scala 27:72]
  wire [1:0] _T_21527 = _T_22121 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21782 = _T_21781 | _T_21527; // @[Mux.scala 27:72]
  wire [1:0] _T_21528 = _T_22123 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21783 = _T_21782 | _T_21528; // @[Mux.scala 27:72]
  wire [1:0] _T_21529 = _T_22125 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21784 = _T_21783 | _T_21529; // @[Mux.scala 27:72]
  wire [1:0] _T_21530 = _T_22127 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21785 = _T_21784 | _T_21530; // @[Mux.scala 27:72]
  wire [1:0] _T_21531 = _T_22129 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21786 = _T_21785 | _T_21531; // @[Mux.scala 27:72]
  wire [1:0] _T_21532 = _T_22131 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21787 = _T_21786 | _T_21532; // @[Mux.scala 27:72]
  wire [1:0] _T_21533 = _T_22133 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21788 = _T_21787 | _T_21533; // @[Mux.scala 27:72]
  wire [1:0] _T_21534 = _T_22135 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21789 = _T_21788 | _T_21534; // @[Mux.scala 27:72]
  wire [1:0] _T_21535 = _T_22137 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21790 = _T_21789 | _T_21535; // @[Mux.scala 27:72]
  wire [1:0] _T_21536 = _T_22139 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21791 = _T_21790 | _T_21536; // @[Mux.scala 27:72]
  wire [1:0] _T_21537 = _T_22141 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21792 = _T_21791 | _T_21537; // @[Mux.scala 27:72]
  wire [1:0] _T_21538 = _T_22143 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21793 = _T_21792 | _T_21538; // @[Mux.scala 27:72]
  wire [1:0] _T_21539 = _T_22145 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21794 = _T_21793 | _T_21539; // @[Mux.scala 27:72]
  wire [1:0] _T_21540 = _T_22147 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21795 = _T_21794 | _T_21540; // @[Mux.scala 27:72]
  wire [1:0] _T_21541 = _T_22149 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21796 = _T_21795 | _T_21541; // @[Mux.scala 27:72]
  wire [1:0] _T_21542 = _T_22151 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21797 = _T_21796 | _T_21542; // @[Mux.scala 27:72]
  wire [1:0] _T_21543 = _T_22153 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21798 = _T_21797 | _T_21543; // @[Mux.scala 27:72]
  wire [1:0] _T_21544 = _T_22155 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21799 = _T_21798 | _T_21544; // @[Mux.scala 27:72]
  wire [1:0] _T_21545 = _T_22157 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21800 = _T_21799 | _T_21545; // @[Mux.scala 27:72]
  wire [1:0] _T_21546 = _T_22159 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21801 = _T_21800 | _T_21546; // @[Mux.scala 27:72]
  wire [1:0] _T_21547 = _T_22161 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21802 = _T_21801 | _T_21547; // @[Mux.scala 27:72]
  wire [1:0] _T_21548 = _T_22163 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21803 = _T_21802 | _T_21548; // @[Mux.scala 27:72]
  wire [1:0] _T_21549 = _T_22165 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21804 = _T_21803 | _T_21549; // @[Mux.scala 27:72]
  wire [1:0] _T_21550 = _T_22167 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21805 = _T_21804 | _T_21550; // @[Mux.scala 27:72]
  wire [1:0] _T_21551 = _T_22169 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21806 = _T_21805 | _T_21551; // @[Mux.scala 27:72]
  wire [1:0] _T_21552 = _T_22171 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21807 = _T_21806 | _T_21552; // @[Mux.scala 27:72]
  wire [1:0] _T_21553 = _T_22173 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21808 = _T_21807 | _T_21553; // @[Mux.scala 27:72]
  wire [1:0] _T_21554 = _T_22175 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21809 = _T_21808 | _T_21554; // @[Mux.scala 27:72]
  wire [1:0] _T_21555 = _T_22177 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21810 = _T_21809 | _T_21555; // @[Mux.scala 27:72]
  wire [1:0] _T_21556 = _T_22179 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21811 = _T_21810 | _T_21556; // @[Mux.scala 27:72]
  wire [1:0] _T_21557 = _T_22181 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21812 = _T_21811 | _T_21557; // @[Mux.scala 27:72]
  wire [1:0] _T_21558 = _T_22183 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21813 = _T_21812 | _T_21558; // @[Mux.scala 27:72]
  wire [1:0] _T_21559 = _T_22185 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21814 = _T_21813 | _T_21559; // @[Mux.scala 27:72]
  wire [1:0] _T_21560 = _T_22187 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21815 = _T_21814 | _T_21560; // @[Mux.scala 27:72]
  wire [1:0] _T_21561 = _T_22189 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21816 = _T_21815 | _T_21561; // @[Mux.scala 27:72]
  wire [1:0] _T_21562 = _T_22191 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21817 = _T_21816 | _T_21562; // @[Mux.scala 27:72]
  wire [1:0] _T_21563 = _T_22193 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21818 = _T_21817 | _T_21563; // @[Mux.scala 27:72]
  wire [1:0] _T_21564 = _T_22195 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21819 = _T_21818 | _T_21564; // @[Mux.scala 27:72]
  wire [1:0] _T_21565 = _T_22197 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21820 = _T_21819 | _T_21565; // @[Mux.scala 27:72]
  wire [1:0] _T_21566 = _T_22199 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21821 = _T_21820 | _T_21566; // @[Mux.scala 27:72]
  wire [1:0] _T_21567 = _T_22201 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21822 = _T_21821 | _T_21567; // @[Mux.scala 27:72]
  wire [1:0] _T_21568 = _T_22203 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21823 = _T_21822 | _T_21568; // @[Mux.scala 27:72]
  wire [1:0] _T_21569 = _T_22205 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21824 = _T_21823 | _T_21569; // @[Mux.scala 27:72]
  wire [1:0] _T_21570 = _T_22207 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21825 = _T_21824 | _T_21570; // @[Mux.scala 27:72]
  wire [1:0] _T_21571 = _T_22209 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21826 = _T_21825 | _T_21571; // @[Mux.scala 27:72]
  wire [1:0] _T_21572 = _T_22211 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21827 = _T_21826 | _T_21572; // @[Mux.scala 27:72]
  wire [1:0] _T_21573 = _T_22213 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21828 = _T_21827 | _T_21573; // @[Mux.scala 27:72]
  wire [1:0] _T_21574 = _T_22215 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21829 = _T_21828 | _T_21574; // @[Mux.scala 27:72]
  wire [1:0] _T_21575 = _T_22217 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21830 = _T_21829 | _T_21575; // @[Mux.scala 27:72]
  wire [1:0] _T_21576 = _T_22219 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21831 = _T_21830 | _T_21576; // @[Mux.scala 27:72]
  wire [1:0] _T_21577 = _T_22221 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21832 = _T_21831 | _T_21577; // @[Mux.scala 27:72]
  wire [1:0] _T_21578 = _T_22223 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21833 = _T_21832 | _T_21578; // @[Mux.scala 27:72]
  wire [1:0] _T_21579 = _T_22225 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21834 = _T_21833 | _T_21579; // @[Mux.scala 27:72]
  wire [1:0] _T_21580 = _T_22227 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21835 = _T_21834 | _T_21580; // @[Mux.scala 27:72]
  wire [1:0] _T_21581 = _T_22229 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21836 = _T_21835 | _T_21581; // @[Mux.scala 27:72]
  wire [1:0] _T_21582 = _T_22231 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21837 = _T_21836 | _T_21582; // @[Mux.scala 27:72]
  wire [1:0] _T_21583 = _T_22233 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21838 = _T_21837 | _T_21583; // @[Mux.scala 27:72]
  wire [1:0] _T_21584 = _T_22235 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21839 = _T_21838 | _T_21584; // @[Mux.scala 27:72]
  wire [1:0] _T_21585 = _T_22237 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21840 = _T_21839 | _T_21585; // @[Mux.scala 27:72]
  wire [1:0] _T_21586 = _T_22239 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21841 = _T_21840 | _T_21586; // @[Mux.scala 27:72]
  wire [1:0] _T_21587 = _T_22241 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21842 = _T_21841 | _T_21587; // @[Mux.scala 27:72]
  wire [1:0] _T_21588 = _T_22243 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21843 = _T_21842 | _T_21588; // @[Mux.scala 27:72]
  wire [1:0] _T_21589 = _T_22245 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21844 = _T_21843 | _T_21589; // @[Mux.scala 27:72]
  wire [1:0] _T_21590 = _T_22247 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21845 = _T_21844 | _T_21590; // @[Mux.scala 27:72]
  wire [1:0] _T_21591 = _T_22249 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21846 = _T_21845 | _T_21591; // @[Mux.scala 27:72]
  wire [1:0] _T_21592 = _T_22251 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21847 = _T_21846 | _T_21592; // @[Mux.scala 27:72]
  wire [1:0] _T_21593 = _T_22253 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21848 = _T_21847 | _T_21593; // @[Mux.scala 27:72]
  wire [1:0] _T_21594 = _T_22255 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21849 = _T_21848 | _T_21594; // @[Mux.scala 27:72]
  wire [1:0] _T_21595 = _T_22257 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21850 = _T_21849 | _T_21595; // @[Mux.scala 27:72]
  wire [1:0] _T_21596 = _T_22259 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21851 = _T_21850 | _T_21596; // @[Mux.scala 27:72]
  wire [1:0] _T_21597 = _T_22261 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21852 = _T_21851 | _T_21597; // @[Mux.scala 27:72]
  wire [1:0] _T_21598 = _T_22263 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21853 = _T_21852 | _T_21598; // @[Mux.scala 27:72]
  wire [1:0] _T_21599 = _T_22265 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21854 = _T_21853 | _T_21599; // @[Mux.scala 27:72]
  wire [1:0] _T_21600 = _T_22267 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21855 = _T_21854 | _T_21600; // @[Mux.scala 27:72]
  wire [1:0] _T_21601 = _T_22269 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21856 = _T_21855 | _T_21601; // @[Mux.scala 27:72]
  wire [1:0] _T_21602 = _T_22271 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21857 = _T_21856 | _T_21602; // @[Mux.scala 27:72]
  wire [1:0] _T_21603 = _T_22273 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21858 = _T_21857 | _T_21603; // @[Mux.scala 27:72]
  wire [1:0] _T_21604 = _T_22275 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21859 = _T_21858 | _T_21604; // @[Mux.scala 27:72]
  wire [1:0] _T_21605 = _T_22277 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21860 = _T_21859 | _T_21605; // @[Mux.scala 27:72]
  wire [1:0] _T_21606 = _T_22279 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21861 = _T_21860 | _T_21606; // @[Mux.scala 27:72]
  wire [1:0] _T_21607 = _T_22281 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21862 = _T_21861 | _T_21607; // @[Mux.scala 27:72]
  wire [1:0] _T_21608 = _T_22283 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21863 = _T_21862 | _T_21608; // @[Mux.scala 27:72]
  wire [1:0] _T_21609 = _T_22285 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21864 = _T_21863 | _T_21609; // @[Mux.scala 27:72]
  wire [1:0] _T_21610 = _T_22287 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21865 = _T_21864 | _T_21610; // @[Mux.scala 27:72]
  wire [1:0] _T_21611 = _T_22289 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21866 = _T_21865 | _T_21611; // @[Mux.scala 27:72]
  wire [1:0] _T_21612 = _T_22291 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21867 = _T_21866 | _T_21612; // @[Mux.scala 27:72]
  wire [1:0] _T_21613 = _T_22293 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21868 = _T_21867 | _T_21613; // @[Mux.scala 27:72]
  wire [1:0] _T_21614 = _T_22295 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21869 = _T_21868 | _T_21614; // @[Mux.scala 27:72]
  wire [1:0] _T_21615 = _T_22297 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21870 = _T_21869 | _T_21615; // @[Mux.scala 27:72]
  wire [1:0] _T_21616 = _T_22299 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21871 = _T_21870 | _T_21616; // @[Mux.scala 27:72]
  wire [1:0] _T_21617 = _T_22301 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21872 = _T_21871 | _T_21617; // @[Mux.scala 27:72]
  wire [1:0] _T_21618 = _T_22303 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21873 = _T_21872 | _T_21618; // @[Mux.scala 27:72]
  wire [1:0] _T_21619 = _T_22305 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21874 = _T_21873 | _T_21619; // @[Mux.scala 27:72]
  wire [1:0] _T_21620 = _T_22307 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21875 = _T_21874 | _T_21620; // @[Mux.scala 27:72]
  wire [1:0] _T_21621 = _T_22309 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21876 = _T_21875 | _T_21621; // @[Mux.scala 27:72]
  wire [1:0] _T_21622 = _T_22311 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21877 = _T_21876 | _T_21622; // @[Mux.scala 27:72]
  wire [1:0] _T_21623 = _T_22313 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21878 = _T_21877 | _T_21623; // @[Mux.scala 27:72]
  wire [1:0] _T_21624 = _T_22315 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21879 = _T_21878 | _T_21624; // @[Mux.scala 27:72]
  wire [1:0] _T_21625 = _T_22317 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21880 = _T_21879 | _T_21625; // @[Mux.scala 27:72]
  wire [1:0] _T_21626 = _T_22319 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21881 = _T_21880 | _T_21626; // @[Mux.scala 27:72]
  wire [1:0] _T_21627 = _T_22321 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21882 = _T_21881 | _T_21627; // @[Mux.scala 27:72]
  wire [1:0] _T_21628 = _T_22323 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21883 = _T_21882 | _T_21628; // @[Mux.scala 27:72]
  wire [1:0] _T_21629 = _T_22325 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21884 = _T_21883 | _T_21629; // @[Mux.scala 27:72]
  wire [1:0] _T_21630 = _T_22327 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21885 = _T_21884 | _T_21630; // @[Mux.scala 27:72]
  wire [1:0] _T_21631 = _T_22329 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21886 = _T_21885 | _T_21631; // @[Mux.scala 27:72]
  wire [1:0] _T_21632 = _T_22331 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21887 = _T_21886 | _T_21632; // @[Mux.scala 27:72]
  wire [1:0] _T_21633 = _T_22333 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21888 = _T_21887 | _T_21633; // @[Mux.scala 27:72]
  wire [1:0] _T_21634 = _T_22335 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21889 = _T_21888 | _T_21634; // @[Mux.scala 27:72]
  wire [1:0] _T_21635 = _T_22337 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21890 = _T_21889 | _T_21635; // @[Mux.scala 27:72]
  wire [1:0] _T_21636 = _T_22339 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21891 = _T_21890 | _T_21636; // @[Mux.scala 27:72]
  wire [1:0] _T_21637 = _T_22341 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21892 = _T_21891 | _T_21637; // @[Mux.scala 27:72]
  wire [1:0] _T_21638 = _T_22343 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21893 = _T_21892 | _T_21638; // @[Mux.scala 27:72]
  wire [1:0] _T_21639 = _T_22345 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21894 = _T_21893 | _T_21639; // @[Mux.scala 27:72]
  wire [1:0] _T_21640 = _T_22347 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21895 = _T_21894 | _T_21640; // @[Mux.scala 27:72]
  wire [1:0] _T_21641 = _T_22349 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21896 = _T_21895 | _T_21641; // @[Mux.scala 27:72]
  wire [1:0] _T_21642 = _T_22351 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21897 = _T_21896 | _T_21642; // @[Mux.scala 27:72]
  wire [1:0] _T_21643 = _T_22353 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21898 = _T_21897 | _T_21643; // @[Mux.scala 27:72]
  wire [1:0] _T_21644 = _T_22355 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21899 = _T_21898 | _T_21644; // @[Mux.scala 27:72]
  wire [1:0] _T_21645 = _T_22357 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21900 = _T_21899 | _T_21645; // @[Mux.scala 27:72]
  wire [1:0] _T_21646 = _T_22359 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21901 = _T_21900 | _T_21646; // @[Mux.scala 27:72]
  wire [1:0] _T_21647 = _T_22361 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21902 = _T_21901 | _T_21647; // @[Mux.scala 27:72]
  wire [1:0] _T_21648 = _T_22363 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21903 = _T_21902 | _T_21648; // @[Mux.scala 27:72]
  wire [1:0] _T_21649 = _T_22365 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21904 = _T_21903 | _T_21649; // @[Mux.scala 27:72]
  wire [1:0] _T_21650 = _T_22367 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21905 = _T_21904 | _T_21650; // @[Mux.scala 27:72]
  wire [1:0] _T_21651 = _T_22369 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21906 = _T_21905 | _T_21651; // @[Mux.scala 27:72]
  wire [1:0] _T_21652 = _T_22371 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21907 = _T_21906 | _T_21652; // @[Mux.scala 27:72]
  wire [1:0] _T_21653 = _T_22373 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21908 = _T_21907 | _T_21653; // @[Mux.scala 27:72]
  wire [1:0] _T_21654 = _T_22375 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21909 = _T_21908 | _T_21654; // @[Mux.scala 27:72]
  wire [1:0] _T_21655 = _T_22377 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21910 = _T_21909 | _T_21655; // @[Mux.scala 27:72]
  wire [1:0] _T_21656 = _T_22379 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21911 = _T_21910 | _T_21656; // @[Mux.scala 27:72]
  wire [1:0] _T_21657 = _T_22381 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21912 = _T_21911 | _T_21657; // @[Mux.scala 27:72]
  wire [1:0] _T_21658 = _T_22383 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21913 = _T_21912 | _T_21658; // @[Mux.scala 27:72]
  wire [1:0] _T_21659 = _T_22385 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21914 = _T_21913 | _T_21659; // @[Mux.scala 27:72]
  wire [1:0] _T_21660 = _T_22387 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21915 = _T_21914 | _T_21660; // @[Mux.scala 27:72]
  wire [1:0] _T_21661 = _T_22389 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21916 = _T_21915 | _T_21661; // @[Mux.scala 27:72]
  wire [1:0] _T_21662 = _T_22391 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21917 = _T_21916 | _T_21662; // @[Mux.scala 27:72]
  wire [1:0] _T_21663 = _T_22393 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21918 = _T_21917 | _T_21663; // @[Mux.scala 27:72]
  wire [1:0] _T_21664 = _T_22395 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21919 = _T_21918 | _T_21664; // @[Mux.scala 27:72]
  wire [1:0] _T_21665 = _T_22397 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21920 = _T_21919 | _T_21665; // @[Mux.scala 27:72]
  wire [1:0] _T_21666 = _T_22399 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21921 = _T_21920 | _T_21666; // @[Mux.scala 27:72]
  wire [1:0] _T_21667 = _T_22401 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21922 = _T_21921 | _T_21667; // @[Mux.scala 27:72]
  wire [1:0] _T_21668 = _T_22403 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21923 = _T_21922 | _T_21668; // @[Mux.scala 27:72]
  wire [1:0] _T_21669 = _T_22405 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21924 = _T_21923 | _T_21669; // @[Mux.scala 27:72]
  wire [1:0] _T_21670 = _T_22407 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21925 = _T_21924 | _T_21670; // @[Mux.scala 27:72]
  wire [1:0] _T_21671 = _T_22409 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21926 = _T_21925 | _T_21671; // @[Mux.scala 27:72]
  wire [1:0] _T_21672 = _T_22411 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21927 = _T_21926 | _T_21672; // @[Mux.scala 27:72]
  wire [1:0] _T_21673 = _T_22413 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21928 = _T_21927 | _T_21673; // @[Mux.scala 27:72]
  wire [1:0] _T_21674 = _T_22415 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21929 = _T_21928 | _T_21674; // @[Mux.scala 27:72]
  wire [1:0] _T_21675 = _T_22417 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21930 = _T_21929 | _T_21675; // @[Mux.scala 27:72]
  wire [1:0] _T_21676 = _T_22419 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21931 = _T_21930 | _T_21676; // @[Mux.scala 27:72]
  wire [1:0] _T_21677 = _T_22421 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21932 = _T_21931 | _T_21677; // @[Mux.scala 27:72]
  wire [1:0] _T_21678 = _T_22423 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21933 = _T_21932 | _T_21678; // @[Mux.scala 27:72]
  wire [1:0] _T_21679 = _T_22425 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21934 = _T_21933 | _T_21679; // @[Mux.scala 27:72]
  wire [1:0] _T_21680 = _T_22427 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21935 = _T_21934 | _T_21680; // @[Mux.scala 27:72]
  wire [1:0] _T_21681 = _T_22429 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21936 = _T_21935 | _T_21681; // @[Mux.scala 27:72]
  wire [1:0] _T_21682 = _T_22431 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21937 = _T_21936 | _T_21682; // @[Mux.scala 27:72]
  wire [1:0] _T_21683 = _T_22433 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21938 = _T_21937 | _T_21683; // @[Mux.scala 27:72]
  wire [1:0] _T_21684 = _T_22435 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21939 = _T_21938 | _T_21684; // @[Mux.scala 27:72]
  wire [1:0] _T_21685 = _T_22437 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21940 = _T_21939 | _T_21685; // @[Mux.scala 27:72]
  wire [1:0] _T_21686 = _T_22439 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21941 = _T_21940 | _T_21686; // @[Mux.scala 27:72]
  wire [1:0] _T_21687 = _T_22441 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21942 = _T_21941 | _T_21687; // @[Mux.scala 27:72]
  wire [1:0] _T_21688 = _T_22443 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21943 = _T_21942 | _T_21688; // @[Mux.scala 27:72]
  wire [1:0] _T_21689 = _T_22445 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21944 = _T_21943 | _T_21689; // @[Mux.scala 27:72]
  wire [1:0] _T_21690 = _T_22447 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21945 = _T_21944 | _T_21690; // @[Mux.scala 27:72]
  wire [1:0] _T_21691 = _T_22449 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21946 = _T_21945 | _T_21691; // @[Mux.scala 27:72]
  wire [1:0] _T_21692 = _T_22451 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21947 = _T_21946 | _T_21692; // @[Mux.scala 27:72]
  wire [1:0] _T_21693 = _T_22453 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21948 = _T_21947 | _T_21693; // @[Mux.scala 27:72]
  wire [1:0] _T_21694 = _T_22455 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21949 = _T_21948 | _T_21694; // @[Mux.scala 27:72]
  wire [1:0] _T_21695 = _T_22457 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21950 = _T_21949 | _T_21695; // @[Mux.scala 27:72]
  wire [1:0] _T_21696 = _T_22459 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21951 = _T_21950 | _T_21696; // @[Mux.scala 27:72]
  wire [1:0] _T_21697 = _T_22461 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21952 = _T_21951 | _T_21697; // @[Mux.scala 27:72]
  wire [1:0] _T_21698 = _T_22463 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21953 = _T_21952 | _T_21698; // @[Mux.scala 27:72]
  wire [1:0] _T_21699 = _T_22465 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21954 = _T_21953 | _T_21699; // @[Mux.scala 27:72]
  wire [1:0] _T_21700 = _T_22467 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_21954 | _T_21700; // @[Mux.scala 27:72]
  wire [1:0] _T_245 = _T_147 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_246 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_245 | _T_246; // @[Mux.scala 27:72]
  wire  _T_263 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 299:45]
  wire  _T_265 = _T_263 & vwayhit_f[0]; // @[ifu_bp_ctl.scala 299:72]
  wire [1:0] bht_dir_f = {_T_260,_T_265}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[ifu_bp_ctl.scala 119:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_147}; // @[Cat.scala 29:58]
  wire  _T_36 = io_exu_bp_exu_mp_btag == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 140:53]
  wire  _T_37 = _T_36 & exu_mp_valid; // @[ifu_bp_ctl.scala 140:73]
  wire  _T_38 = _T_37 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 140:88]
  wire  _T_39 = io_exu_bp_exu_mp_index == btb_rd_addr_f; // @[ifu_bp_ctl.scala 140:124]
  wire  fetch_mp_collision_f = _T_38 & _T_39; // @[ifu_bp_ctl.scala 140:109]
  wire  _T_40 = io_exu_bp_exu_mp_btag == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 141:56]
  wire  _T_41 = _T_40 & exu_mp_valid; // @[ifu_bp_ctl.scala 141:79]
  wire  _T_42 = _T_41 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 141:94]
  wire  _T_43 = io_exu_bp_exu_mp_index == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 141:130]
  wire  fetch_mp_collision_p1_f = _T_42 & _T_43; // @[ifu_bp_ctl.scala 141:115]
  wire [1:0] _T_153 = ~vwayhit_f; // @[ifu_bp_ctl.scala 194:44]
  reg  exu_mp_way_f; // @[Reg.scala 27:20]
  wire [255:0] fetch_wrindex_dec = 256'h1 << btb_rd_addr_f; // @[ifu_bp_ctl.scala 213:31]
  reg [255:0] btb_lru_b0_f; // @[Reg.scala 27:20]
  wire [255:0] _T_181 = fetch_wrindex_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 239:78]
  wire  _T_182 = |_T_181; // @[ifu_bp_ctl.scala 239:94]
  wire  btb_lru_rd_f = fetch_mp_collision_f ? exu_mp_way_f : _T_182; // @[ifu_bp_ctl.scala 239:25]
  wire [1:0] _T_188 = {btb_lru_rd_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_192 = _T_147 ? _T_188 : 2'h0; // @[Mux.scala 27:72]
  wire [255:0] fetch_wrindex_p1_dec = 256'h1 << btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 216:34]
  wire [255:0] _T_184 = fetch_wrindex_p1_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 241:87]
  wire  _T_185 = |_T_184; // @[ifu_bp_ctl.scala 241:103]
  wire  btb_lru_rd_p1_f = fetch_mp_collision_p1_f ? exu_mp_way_f : _T_185; // @[ifu_bp_ctl.scala 241:28]
  wire [1:0] _T_191 = {btb_lru_rd_p1_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_193 = io_ifc_fetch_addr_f[0] ? _T_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_192 | _T_193; // @[Mux.scala 27:72]
  wire [1:0] _T_154 = _T_153 & btb_vlru_rd_f; // @[ifu_bp_ctl.scala 194:55]
  wire [1:0] _T_204 = _T_147 ? tag_match_way1_expanded_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_203 = {tag_match_way1_expanded_p1_f[0],tag_match_way1_expanded_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_205 = io_ifc_fetch_addr_f[0] ? _T_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_204 | _T_205; // @[Mux.scala 27:72]
  wire [255:0] mp_wrindex_dec = 256'h1 << io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 210:28]
  wire [255:0] _T_157 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] mp_wrlru_b0 = mp_wrindex_dec & _T_157; // @[ifu_bp_ctl.scala 219:36]
  wire  _T_160 = vwayhit_f[0] | vwayhit_f[1]; // @[ifu_bp_ctl.scala 222:42]
  wire  _T_161 = _T_160 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 222:58]
  wire  lru_update_valid_f = _T_161 & _T; // @[ifu_bp_ctl.scala 222:79]
  wire [255:0] _T_164 = lru_update_valid_f ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] fetch_wrlru_b0 = fetch_wrindex_dec & _T_164; // @[ifu_bp_ctl.scala 224:42]
  wire [255:0] fetch_wrlru_p1_b0 = fetch_wrindex_p1_dec & _T_164; // @[ifu_bp_ctl.scala 225:48]
  wire [255:0] _T_167 = ~mp_wrlru_b0; // @[ifu_bp_ctl.scala 227:25]
  wire [255:0] _T_168 = ~fetch_wrlru_b0; // @[ifu_bp_ctl.scala 227:40]
  wire [255:0] btb_lru_b0_hold = _T_167 & _T_168; // @[ifu_bp_ctl.scala 227:38]
  wire  _T_170 = ~io_exu_bp_exu_mp_pkt_bits_way; // @[ifu_bp_ctl.scala 234:39]
  wire [255:0] _T_173 = _T_170 ? mp_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_174 = tag_match_way0_f ? fetch_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_175 = tag_match_way0_p1_f ? fetch_wrlru_p1_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_176 = _T_173 | _T_174; // @[Mux.scala 27:72]
  wire [255:0] _T_177 = _T_176 | _T_175; // @[Mux.scala 27:72]
  wire [255:0] _T_179 = btb_lru_b0_hold & btb_lru_b0_f; // @[ifu_bp_ctl.scala 236:73]
  wire [255:0] btb_lru_b0_ns = _T_177 | _T_179; // @[ifu_bp_ctl.scala 236:55]
  wire  _T_208 = io_ifc_fetch_req_f | exu_mp_valid; // @[ifu_bp_ctl.scala 251:60]
  wire [15:0] _T_223 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_224 = btb_sel_f[0] ? btb_vbank0_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] btb_sel_data_f = _T_223 | _T_224; // @[Mux.scala 27:72]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 267:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[ifu_bp_ctl.scala 268:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[ifu_bp_ctl.scala 269:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[ifu_bp_ctl.scala 270:36]
  wire [1:0] _T_273 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_273; // @[ifu_bp_ctl.scala 305:34]
  wire [1:0] _T_227 = vwayhit_f & hist1_raw; // @[ifu_bp_ctl.scala 277:39]
  wire  _T_228 = |_T_227; // @[ifu_bp_ctl.scala 277:52]
  wire  _T_229 = _T_228 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 277:56]
  wire  _T_230 = ~leak_one_f_d1; // @[ifu_bp_ctl.scala 277:79]
  wire  _T_231 = _T_229 & _T_230; // @[ifu_bp_ctl.scala 277:77]
  wire  _T_232 = ~io_dec_bp_dec_tlu_bpred_disable; // @[ifu_bp_ctl.scala 277:96]
  wire  _T_268 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[ifu_bp_ctl.scala 302:51]
  wire  _T_269 = ~io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 302:69]
  wire  _T_279 = vwayhit_f[1] & btb_vbank1_rd_data_f[4]; // @[ifu_bp_ctl.scala 311:34]
  wire  _T_282 = vwayhit_f[0] & btb_vbank0_rd_data_f[4]; // @[ifu_bp_ctl.scala 312:34]
  wire  _T_285 = ~btb_vbank1_rd_data_f[2]; // @[ifu_bp_ctl.scala 315:37]
  wire  _T_286 = vwayhit_f[1] & _T_285; // @[ifu_bp_ctl.scala 315:35]
  wire  _T_288 = _T_286 & btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 315:65]
  wire  _T_291 = ~btb_vbank0_rd_data_f[2]; // @[ifu_bp_ctl.scala 316:37]
  wire  _T_292 = vwayhit_f[0] & _T_291; // @[ifu_bp_ctl.scala 316:35]
  wire  _T_294 = _T_292 & btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 316:65]
  wire [1:0] num_valids = vwayhit_f[1] + vwayhit_f[0]; // @[ifu_bp_ctl.scala 319:35]
  wire [1:0] _T_297 = btb_sel_f & bht_dir_f; // @[ifu_bp_ctl.scala 322:28]
  wire  final_h = |_T_297; // @[ifu_bp_ctl.scala 322:41]
  wire  _T_298 = num_valids == 2'h2; // @[ifu_bp_ctl.scala 326:41]
  wire [7:0] _T_302 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_303 = num_valids == 2'h1; // @[ifu_bp_ctl.scala 327:41]
  wire [7:0] _T_306 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_307 = num_valids == 2'h0; // @[ifu_bp_ctl.scala 328:41]
  wire [7:0] _T_310 = _T_298 ? _T_302 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_311 = _T_303 ? _T_306 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_312 = _T_307 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_313 = _T_310 | _T_311; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_313 | _T_312; // @[Mux.scala 27:72]
  reg  exu_flush_final_d1; // @[Reg.scala 27:20]
  wire  _T_316 = ~exu_flush_final_d1; // @[ifu_bp_ctl.scala 337:27]
  wire  _T_317 = _T_316 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 337:47]
  wire  _T_318 = _T_317 & io_ic_hit_f; // @[ifu_bp_ctl.scala 337:70]
  wire  _T_320 = _T_318 & _T_230; // @[ifu_bp_ctl.scala 337:84]
  wire  _T_323 = io_ifc_fetch_req_f & io_ic_hit_f; // @[ifu_bp_ctl.scala 338:70]
  wire  _T_325 = _T_323 & _T_230; // @[ifu_bp_ctl.scala 338:84]
  wire  _T_326 = ~_T_325; // @[ifu_bp_ctl.scala 338:49]
  wire  _T_327 = _T_316 & _T_326; // @[ifu_bp_ctl.scala 338:47]
  wire [7:0] _T_329 = exu_flush_final_d1 ? io_exu_bp_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_330 = _T_320 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_331 = _T_327 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_332 = _T_329 | _T_330; // @[Mux.scala 27:72]
  wire [7:0] fghr_ns = _T_332 | _T_331; // @[Mux.scala 27:72]
  wire  _T_336 = leak_one_f ^ leak_one_f_d1; // @[lib.scala 453:21]
  wire  _T_337 = |_T_336; // @[lib.scala 453:29]
  wire  _T_340 = io_exu_bp_exu_mp_pkt_bits_way ^ exu_mp_way_f; // @[lib.scala 453:21]
  wire  _T_341 = |_T_340; // @[lib.scala 453:29]
  wire  _T_344 = io_exu_flush_final ^ exu_flush_final_d1; // @[lib.scala 475:21]
  wire  _T_345 = |_T_344; // @[lib.scala 475:29]
  wire [7:0] _T_348 = fghr_ns ^ fghr; // @[lib.scala 453:21]
  wire  _T_349 = |_T_348; // @[lib.scala 453:29]
  wire [1:0] _T_352 = io_dec_bp_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_353 = ~_T_352; // @[ifu_bp_ctl.scala 350:36]
  wire  _T_357 = ~fetch_start_f[0]; // @[ifu_bp_ctl.scala 354:36]
  wire  _T_358 = bht_dir_f[0] & _T_357; // @[ifu_bp_ctl.scala 354:34]
  wire  _T_362 = _T_14 & fetch_start_f[0]; // @[ifu_bp_ctl.scala 354:72]
  wire  _T_363 = _T_358 | _T_362; // @[ifu_bp_ctl.scala 354:55]
  wire  _T_366 = bht_dir_f[0] & fetch_start_f[0]; // @[ifu_bp_ctl.scala 355:34]
  wire  _T_371 = _T_14 & _T_357; // @[ifu_bp_ctl.scala 355:71]
  wire  _T_372 = _T_366 | _T_371; // @[ifu_bp_ctl.scala 355:54]
  wire [1:0] bloc_f = {_T_363,_T_372}; // @[Cat.scala 29:58]
  wire  _T_376 = _T_14 & io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 357:35]
  wire  _T_377 = ~btb_rd_pc4_f; // @[ifu_bp_ctl.scala 357:62]
  wire  use_fa_plus = _T_376 & _T_377; // @[ifu_bp_ctl.scala 357:60]
  wire  _T_380 = fetch_start_f[0] & btb_sel_f[0]; // @[ifu_bp_ctl.scala 359:44]
  wire  btb_fg_crossing_f = _T_380 & btb_rd_pc4_f; // @[ifu_bp_ctl.scala 359:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[ifu_bp_ctl.scala 360:43]
  wire  _T_384 = io_ifc_fetch_req_f & _T_269; // @[ifu_bp_ctl.scala 361:117]
  wire  _T_385 = _T_384 & io_ic_hit_f; // @[ifu_bp_ctl.scala 361:142]
  reg [29:0] ifc_fetch_adder_prior; // @[Reg.scala 27:20]
  wire  _T_390 = ~btb_fg_crossing_f; // @[ifu_bp_ctl.scala 366:32]
  wire  _T_391 = ~use_fa_plus; // @[ifu_bp_ctl.scala 366:53]
  wire  _T_392 = _T_390 & _T_391; // @[ifu_bp_ctl.scala 366:51]
  wire [29:0] _T_395 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_396 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_397 = _T_392 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_398 = _T_395 | _T_396; // @[Mux.scala 27:72]
  wire [29:0] adder_pc_in_f = _T_398 | _T_397; // @[Mux.scala 27:72]
  wire [31:0] _T_402 = {adder_pc_in_f,bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_403 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_406 = _T_402[12:1] + _T_403[12:1]; // @[lib.scala 68:31]
  wire [18:0] _T_409 = _T_402[31:13] + 19'h1; // @[lib.scala 69:27]
  wire [18:0] _T_412 = _T_402[31:13] - 19'h1; // @[lib.scala 70:27]
  wire  _T_415 = ~_T_406[12]; // @[lib.scala 72:28]
  wire  _T_416 = _T_403[12] ^ _T_415; // @[lib.scala 72:26]
  wire  _T_419 = ~_T_403[12]; // @[lib.scala 73:20]
  wire  _T_421 = _T_419 & _T_406[12]; // @[lib.scala 73:26]
  wire  _T_425 = _T_403[12] & _T_415; // @[lib.scala 74:26]
  wire [18:0] _T_427 = _T_416 ? _T_402[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_428 = _T_421 ? _T_409 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_429 = _T_425 ? _T_412 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_430 = _T_427 | _T_428; // @[Mux.scala 27:72]
  wire [18:0] _T_431 = _T_430 | _T_429; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_431,_T_406[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_435 = ~btb_rd_call_f; // @[ifu_bp_ctl.scala 374:55]
  wire  _T_436 = btb_rd_ret_f & _T_435; // @[ifu_bp_ctl.scala 374:53]
  reg [31:0] rets_out_0; // @[Reg.scala 27:20]
  wire  _T_438 = _T_436 & rets_out_0[0]; // @[ifu_bp_ctl.scala 374:70]
  wire  _T_439 = _T_438 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 374:87]
  wire [30:0] _T_441 = _T_439 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_443 = _T_441 & rets_out_0[31:1]; // @[ifu_bp_ctl.scala 374:113]
  wire  _T_448 = ~_T_438; // @[ifu_bp_ctl.scala 375:15]
  wire  _T_449 = _T_448 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 375:65]
  wire [30:0] _T_451 = _T_449 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_453 = _T_451 & bp_btb_target_adder_f[31:1]; // @[ifu_bp_ctl.scala 375:91]
  wire [12:0] _T_461 = {11'h0,_T_377,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_464 = _T_402[12:1] + _T_461[12:1]; // @[lib.scala 68:31]
  wire  _T_473 = ~_T_464[12]; // @[lib.scala 72:28]
  wire  _T_474 = _T_461[12] ^ _T_473; // @[lib.scala 72:26]
  wire  _T_477 = ~_T_461[12]; // @[lib.scala 73:20]
  wire  _T_479 = _T_477 & _T_464[12]; // @[lib.scala 73:26]
  wire  _T_483 = _T_461[12] & _T_473; // @[lib.scala 74:26]
  wire [18:0] _T_485 = _T_474 ? _T_402[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_486 = _T_479 ? _T_409 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_487 = _T_483 ? _T_412 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_488 = _T_485 | _T_486; // @[Mux.scala 27:72]
  wire [18:0] _T_489 = _T_488 | _T_487; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_489,_T_464[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_493 = ~btb_rd_ret_f; // @[ifu_bp_ctl.scala 379:33]
  wire  _T_494 = btb_rd_call_f & _T_493; // @[ifu_bp_ctl.scala 379:31]
  wire  rs_push = _T_494 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 379:47]
  wire  rs_pop = _T_436 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 380:46]
  wire  _T_497 = ~rs_push; // @[ifu_bp_ctl.scala 381:17]
  wire  _T_498 = ~rs_pop; // @[ifu_bp_ctl.scala 381:28]
  wire  rs_hold = _T_497 & _T_498; // @[ifu_bp_ctl.scala 381:26]
  wire  rsenable_0 = ~rs_hold; // @[ifu_bp_ctl.scala 383:60]
  wire  rsenable_1 = rs_push | rs_pop; // @[ifu_bp_ctl.scala 383:119]
  wire [31:0] _T_501 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_503 = rs_push ? _T_501 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[Reg.scala 27:20]
  wire [31:0] _T_504 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_0 = _T_503 | _T_504; // @[Mux.scala 27:72]
  wire [31:0] _T_508 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[Reg.scala 27:20]
  wire [31:0] _T_509 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_1 = _T_508 | _T_509; // @[Mux.scala 27:72]
  wire [31:0] _T_513 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[Reg.scala 27:20]
  wire [31:0] _T_514 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_2 = _T_513 | _T_514; // @[Mux.scala 27:72]
  wire [31:0] _T_518 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[Reg.scala 27:20]
  wire [31:0] _T_519 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_3 = _T_518 | _T_519; // @[Mux.scala 27:72]
  wire [31:0] _T_523 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[Reg.scala 27:20]
  wire [31:0] _T_524 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_4 = _T_523 | _T_524; // @[Mux.scala 27:72]
  wire [31:0] _T_528 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[Reg.scala 27:20]
  wire [31:0] _T_529 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_5 = _T_528 | _T_529; // @[Mux.scala 27:72]
  wire [31:0] _T_533 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[Reg.scala 27:20]
  wire [31:0] _T_534 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_6 = _T_533 | _T_534; // @[Mux.scala 27:72]
  wire  _T_552 = ~dec_tlu_error_wb; // @[ifu_bp_ctl.scala 395:35]
  wire  btb_valid = exu_mp_valid & _T_552; // @[ifu_bp_ctl.scala 395:32]
  wire  _T_553 = io_exu_bp_exu_mp_pkt_bits_pcall | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 399:89]
  wire  _T_554 = io_exu_bp_exu_mp_pkt_bits_pret | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 399:113]
  wire [21:0] btb_wr_data = {io_exu_bp_exu_mp_btag,io_exu_bp_exu_mp_pkt_bits_toffset,io_exu_bp_exu_mp_pkt_bits_pc4,io_exu_bp_exu_mp_pkt_bits_boffset,_T_553,_T_554,btb_valid}; // @[Cat.scala 29:58]
  wire  _T_560 = exu_mp_valid & io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu_bp_ctl.scala 400:41]
  wire  _T_561 = ~io_exu_bp_exu_mp_pkt_valid; // @[ifu_bp_ctl.scala 400:59]
  wire  exu_mp_valid_write = _T_560 & _T_561; // @[ifu_bp_ctl.scala 400:57]
  wire  middle_of_bank = io_exu_bp_exu_mp_pkt_bits_pc4 ^ io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu_bp_ctl.scala 401:35]
  wire  _T_562 = ~io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu_bp_ctl.scala 404:43]
  wire  _T_563 = exu_mp_valid & _T_562; // @[ifu_bp_ctl.scala 404:41]
  wire  _T_564 = ~io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu_bp_ctl.scala 404:58]
  wire  _T_565 = _T_563 & _T_564; // @[ifu_bp_ctl.scala 404:56]
  wire  _T_566 = ~io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 404:72]
  wire  _T_567 = _T_565 & _T_566; // @[ifu_bp_ctl.scala 404:70]
  wire [1:0] _T_569 = _T_567 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_570 = ~middle_of_bank; // @[ifu_bp_ctl.scala 404:106]
  wire [1:0] _T_571 = {middle_of_bank,_T_570}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_569 & _T_571; // @[ifu_bp_ctl.scala 404:84]
  wire [1:0] _T_573 = io_dec_bp_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_574 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu_bp_ctl.scala 405:75]
  wire [1:0] _T_575 = {io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,_T_574}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_573 & _T_575; // @[ifu_bp_ctl.scala 405:46]
  wire [9:0] _T_576 = {io_exu_bp_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] mp_hashed = _T_576[9:2] ^ io_exu_bp_exu_mp_eghr; // @[lib.scala 56:35]
  wire [9:0] _T_579 = {io_exu_bp_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] br0_hashed_wb = _T_579[9:2] ^ io_exu_bp_exu_i0_br_fghr_r; // @[lib.scala 56:35]
  wire  _T_589 = _T_170 & exu_mp_valid_write; // @[ifu_bp_ctl.scala 424:39]
  wire  _T_591 = _T_589 & _T_552; // @[ifu_bp_ctl.scala 424:60]
  wire  _T_592 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu_bp_ctl.scala 424:87]
  wire  _T_593 = _T_592 & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 424:104]
  wire  btb_wr_en_way0 = _T_591 | _T_593; // @[ifu_bp_ctl.scala 424:83]
  wire  _T_594 = io_exu_bp_exu_mp_pkt_bits_way & exu_mp_valid_write; // @[ifu_bp_ctl.scala 425:36]
  wire  _T_596 = _T_594 & _T_552; // @[ifu_bp_ctl.scala 425:57]
  wire  _T_597 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 425:98]
  wire  btb_wr_en_way1 = _T_596 | _T_597; // @[ifu_bp_ctl.scala 425:80]
  wire [7:0] btb_wr_addr = dec_tlu_error_wb ? io_exu_bp_exu_i0_br_index_r : io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 428:24]
  wire  _T_613 = btb_wr_addr == 8'h0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_614 = _T_613 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_616 = btb_wr_addr == 8'h1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_617 = _T_616 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_619 = btb_wr_addr == 8'h2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_620 = _T_619 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_622 = btb_wr_addr == 8'h3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_623 = _T_622 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_625 = btb_wr_addr == 8'h4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_626 = _T_625 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_628 = btb_wr_addr == 8'h5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_629 = _T_628 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_631 = btb_wr_addr == 8'h6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_632 = _T_631 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_634 = btb_wr_addr == 8'h7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_635 = _T_634 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_637 = btb_wr_addr == 8'h8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_638 = _T_637 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_640 = btb_wr_addr == 8'h9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_641 = _T_640 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_643 = btb_wr_addr == 8'ha; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_644 = _T_643 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_646 = btb_wr_addr == 8'hb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_647 = _T_646 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_649 = btb_wr_addr == 8'hc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_650 = _T_649 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_652 = btb_wr_addr == 8'hd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_653 = _T_652 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_655 = btb_wr_addr == 8'he; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_656 = _T_655 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_658 = btb_wr_addr == 8'hf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_659 = _T_658 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_661 = btb_wr_addr == 8'h10; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_662 = _T_661 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_664 = btb_wr_addr == 8'h11; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_665 = _T_664 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_667 = btb_wr_addr == 8'h12; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_668 = _T_667 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_670 = btb_wr_addr == 8'h13; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_671 = _T_670 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_673 = btb_wr_addr == 8'h14; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_674 = _T_673 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_676 = btb_wr_addr == 8'h15; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_677 = _T_676 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_679 = btb_wr_addr == 8'h16; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_680 = _T_679 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_682 = btb_wr_addr == 8'h17; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_683 = _T_682 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_685 = btb_wr_addr == 8'h18; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_686 = _T_685 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_688 = btb_wr_addr == 8'h19; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_689 = _T_688 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_691 = btb_wr_addr == 8'h1a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_692 = _T_691 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_694 = btb_wr_addr == 8'h1b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_695 = _T_694 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_697 = btb_wr_addr == 8'h1c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_698 = _T_697 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_700 = btb_wr_addr == 8'h1d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_701 = _T_700 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_703 = btb_wr_addr == 8'h1e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_704 = _T_703 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_706 = btb_wr_addr == 8'h1f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_707 = _T_706 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_709 = btb_wr_addr == 8'h20; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_710 = _T_709 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_712 = btb_wr_addr == 8'h21; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_713 = _T_712 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_715 = btb_wr_addr == 8'h22; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_716 = _T_715 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_718 = btb_wr_addr == 8'h23; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_719 = _T_718 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_721 = btb_wr_addr == 8'h24; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_722 = _T_721 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_724 = btb_wr_addr == 8'h25; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_725 = _T_724 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_727 = btb_wr_addr == 8'h26; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_728 = _T_727 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_730 = btb_wr_addr == 8'h27; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_731 = _T_730 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_733 = btb_wr_addr == 8'h28; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_734 = _T_733 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_736 = btb_wr_addr == 8'h29; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_737 = _T_736 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_739 = btb_wr_addr == 8'h2a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_740 = _T_739 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_742 = btb_wr_addr == 8'h2b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_743 = _T_742 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_745 = btb_wr_addr == 8'h2c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_746 = _T_745 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_748 = btb_wr_addr == 8'h2d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_749 = _T_748 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_751 = btb_wr_addr == 8'h2e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_752 = _T_751 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_754 = btb_wr_addr == 8'h2f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_755 = _T_754 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_757 = btb_wr_addr == 8'h30; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_758 = _T_757 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_760 = btb_wr_addr == 8'h31; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_761 = _T_760 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_763 = btb_wr_addr == 8'h32; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_764 = _T_763 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_766 = btb_wr_addr == 8'h33; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_767 = _T_766 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_769 = btb_wr_addr == 8'h34; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_770 = _T_769 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_772 = btb_wr_addr == 8'h35; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_773 = _T_772 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_775 = btb_wr_addr == 8'h36; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_776 = _T_775 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_778 = btb_wr_addr == 8'h37; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_779 = _T_778 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_781 = btb_wr_addr == 8'h38; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_782 = _T_781 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_784 = btb_wr_addr == 8'h39; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_785 = _T_784 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_787 = btb_wr_addr == 8'h3a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_788 = _T_787 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_790 = btb_wr_addr == 8'h3b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_791 = _T_790 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_793 = btb_wr_addr == 8'h3c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_794 = _T_793 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_796 = btb_wr_addr == 8'h3d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_797 = _T_796 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_799 = btb_wr_addr == 8'h3e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_800 = _T_799 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_802 = btb_wr_addr == 8'h3f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_803 = _T_802 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_805 = btb_wr_addr == 8'h40; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_806 = _T_805 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_808 = btb_wr_addr == 8'h41; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_809 = _T_808 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_811 = btb_wr_addr == 8'h42; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_812 = _T_811 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_814 = btb_wr_addr == 8'h43; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_815 = _T_814 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_817 = btb_wr_addr == 8'h44; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_818 = _T_817 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_820 = btb_wr_addr == 8'h45; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_821 = _T_820 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_823 = btb_wr_addr == 8'h46; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_824 = _T_823 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_826 = btb_wr_addr == 8'h47; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_827 = _T_826 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_829 = btb_wr_addr == 8'h48; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_830 = _T_829 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_832 = btb_wr_addr == 8'h49; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_833 = _T_832 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_835 = btb_wr_addr == 8'h4a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_836 = _T_835 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_838 = btb_wr_addr == 8'h4b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_839 = _T_838 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_841 = btb_wr_addr == 8'h4c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_842 = _T_841 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_844 = btb_wr_addr == 8'h4d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_845 = _T_844 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_847 = btb_wr_addr == 8'h4e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_848 = _T_847 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_850 = btb_wr_addr == 8'h4f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_851 = _T_850 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_853 = btb_wr_addr == 8'h50; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_854 = _T_853 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_856 = btb_wr_addr == 8'h51; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_857 = _T_856 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_859 = btb_wr_addr == 8'h52; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_860 = _T_859 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_862 = btb_wr_addr == 8'h53; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_863 = _T_862 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_865 = btb_wr_addr == 8'h54; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_866 = _T_865 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_868 = btb_wr_addr == 8'h55; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_869 = _T_868 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_871 = btb_wr_addr == 8'h56; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_872 = _T_871 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_874 = btb_wr_addr == 8'h57; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_875 = _T_874 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_877 = btb_wr_addr == 8'h58; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_878 = _T_877 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_880 = btb_wr_addr == 8'h59; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_881 = _T_880 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_883 = btb_wr_addr == 8'h5a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_884 = _T_883 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_886 = btb_wr_addr == 8'h5b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_887 = _T_886 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_889 = btb_wr_addr == 8'h5c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_890 = _T_889 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_892 = btb_wr_addr == 8'h5d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_893 = _T_892 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_895 = btb_wr_addr == 8'h5e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_896 = _T_895 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_898 = btb_wr_addr == 8'h5f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_899 = _T_898 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_901 = btb_wr_addr == 8'h60; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_902 = _T_901 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_904 = btb_wr_addr == 8'h61; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_905 = _T_904 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_907 = btb_wr_addr == 8'h62; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_908 = _T_907 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_910 = btb_wr_addr == 8'h63; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_911 = _T_910 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_913 = btb_wr_addr == 8'h64; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_914 = _T_913 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_916 = btb_wr_addr == 8'h65; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_917 = _T_916 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_919 = btb_wr_addr == 8'h66; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_920 = _T_919 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_922 = btb_wr_addr == 8'h67; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_923 = _T_922 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_925 = btb_wr_addr == 8'h68; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_926 = _T_925 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_928 = btb_wr_addr == 8'h69; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_929 = _T_928 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_931 = btb_wr_addr == 8'h6a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_932 = _T_931 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_934 = btb_wr_addr == 8'h6b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_935 = _T_934 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_937 = btb_wr_addr == 8'h6c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_938 = _T_937 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_940 = btb_wr_addr == 8'h6d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_941 = _T_940 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_943 = btb_wr_addr == 8'h6e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_944 = _T_943 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_946 = btb_wr_addr == 8'h6f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_947 = _T_946 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_949 = btb_wr_addr == 8'h70; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_950 = _T_949 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_952 = btb_wr_addr == 8'h71; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_953 = _T_952 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_955 = btb_wr_addr == 8'h72; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_956 = _T_955 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_958 = btb_wr_addr == 8'h73; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_959 = _T_958 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_961 = btb_wr_addr == 8'h74; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_962 = _T_961 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_964 = btb_wr_addr == 8'h75; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_965 = _T_964 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_967 = btb_wr_addr == 8'h76; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_968 = _T_967 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_970 = btb_wr_addr == 8'h77; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_971 = _T_970 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_973 = btb_wr_addr == 8'h78; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_974 = _T_973 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_976 = btb_wr_addr == 8'h79; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_977 = _T_976 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_979 = btb_wr_addr == 8'h7a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_980 = _T_979 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_982 = btb_wr_addr == 8'h7b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_983 = _T_982 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_985 = btb_wr_addr == 8'h7c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_986 = _T_985 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_988 = btb_wr_addr == 8'h7d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_989 = _T_988 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_991 = btb_wr_addr == 8'h7e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_992 = _T_991 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_994 = btb_wr_addr == 8'h7f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_995 = _T_994 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_997 = btb_wr_addr == 8'h80; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_998 = _T_997 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1000 = btb_wr_addr == 8'h81; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1001 = _T_1000 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1003 = btb_wr_addr == 8'h82; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1004 = _T_1003 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1006 = btb_wr_addr == 8'h83; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1007 = _T_1006 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1009 = btb_wr_addr == 8'h84; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1010 = _T_1009 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1012 = btb_wr_addr == 8'h85; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1013 = _T_1012 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1015 = btb_wr_addr == 8'h86; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1016 = _T_1015 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1018 = btb_wr_addr == 8'h87; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1019 = _T_1018 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1021 = btb_wr_addr == 8'h88; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1022 = _T_1021 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1024 = btb_wr_addr == 8'h89; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1025 = _T_1024 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1027 = btb_wr_addr == 8'h8a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1028 = _T_1027 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1030 = btb_wr_addr == 8'h8b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1031 = _T_1030 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1033 = btb_wr_addr == 8'h8c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1034 = _T_1033 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1036 = btb_wr_addr == 8'h8d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1037 = _T_1036 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1039 = btb_wr_addr == 8'h8e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1040 = _T_1039 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1042 = btb_wr_addr == 8'h8f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1043 = _T_1042 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1045 = btb_wr_addr == 8'h90; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1046 = _T_1045 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1048 = btb_wr_addr == 8'h91; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1049 = _T_1048 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1051 = btb_wr_addr == 8'h92; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1052 = _T_1051 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1054 = btb_wr_addr == 8'h93; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1055 = _T_1054 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1057 = btb_wr_addr == 8'h94; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1058 = _T_1057 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1060 = btb_wr_addr == 8'h95; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1061 = _T_1060 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1063 = btb_wr_addr == 8'h96; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1064 = _T_1063 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1066 = btb_wr_addr == 8'h97; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1067 = _T_1066 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1069 = btb_wr_addr == 8'h98; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1070 = _T_1069 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1072 = btb_wr_addr == 8'h99; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1073 = _T_1072 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1075 = btb_wr_addr == 8'h9a; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1076 = _T_1075 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1078 = btb_wr_addr == 8'h9b; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1079 = _T_1078 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1081 = btb_wr_addr == 8'h9c; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1082 = _T_1081 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1084 = btb_wr_addr == 8'h9d; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1085 = _T_1084 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1087 = btb_wr_addr == 8'h9e; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1088 = _T_1087 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1090 = btb_wr_addr == 8'h9f; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1091 = _T_1090 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1093 = btb_wr_addr == 8'ha0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1094 = _T_1093 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1096 = btb_wr_addr == 8'ha1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1097 = _T_1096 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1099 = btb_wr_addr == 8'ha2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1100 = _T_1099 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1102 = btb_wr_addr == 8'ha3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1103 = _T_1102 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1105 = btb_wr_addr == 8'ha4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1106 = _T_1105 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1108 = btb_wr_addr == 8'ha5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1109 = _T_1108 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1111 = btb_wr_addr == 8'ha6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1112 = _T_1111 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1114 = btb_wr_addr == 8'ha7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1115 = _T_1114 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1117 = btb_wr_addr == 8'ha8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1118 = _T_1117 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1120 = btb_wr_addr == 8'ha9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1121 = _T_1120 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1123 = btb_wr_addr == 8'haa; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1124 = _T_1123 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1126 = btb_wr_addr == 8'hab; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1127 = _T_1126 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1129 = btb_wr_addr == 8'hac; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1130 = _T_1129 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1132 = btb_wr_addr == 8'had; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1133 = _T_1132 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1135 = btb_wr_addr == 8'hae; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1136 = _T_1135 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1138 = btb_wr_addr == 8'haf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1139 = _T_1138 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1141 = btb_wr_addr == 8'hb0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1142 = _T_1141 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1144 = btb_wr_addr == 8'hb1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1145 = _T_1144 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1147 = btb_wr_addr == 8'hb2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1148 = _T_1147 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1150 = btb_wr_addr == 8'hb3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1151 = _T_1150 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1153 = btb_wr_addr == 8'hb4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1154 = _T_1153 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1156 = btb_wr_addr == 8'hb5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1157 = _T_1156 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1159 = btb_wr_addr == 8'hb6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1160 = _T_1159 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1162 = btb_wr_addr == 8'hb7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1163 = _T_1162 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1165 = btb_wr_addr == 8'hb8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1166 = _T_1165 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1168 = btb_wr_addr == 8'hb9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1169 = _T_1168 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1171 = btb_wr_addr == 8'hba; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1172 = _T_1171 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1174 = btb_wr_addr == 8'hbb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1175 = _T_1174 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1177 = btb_wr_addr == 8'hbc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1178 = _T_1177 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1180 = btb_wr_addr == 8'hbd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1181 = _T_1180 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1183 = btb_wr_addr == 8'hbe; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1184 = _T_1183 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1186 = btb_wr_addr == 8'hbf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1187 = _T_1186 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1189 = btb_wr_addr == 8'hc0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1190 = _T_1189 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1192 = btb_wr_addr == 8'hc1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1193 = _T_1192 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1195 = btb_wr_addr == 8'hc2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1196 = _T_1195 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1198 = btb_wr_addr == 8'hc3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1199 = _T_1198 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1201 = btb_wr_addr == 8'hc4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1202 = _T_1201 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1204 = btb_wr_addr == 8'hc5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1205 = _T_1204 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1207 = btb_wr_addr == 8'hc6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1208 = _T_1207 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1210 = btb_wr_addr == 8'hc7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1211 = _T_1210 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1213 = btb_wr_addr == 8'hc8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1214 = _T_1213 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1216 = btb_wr_addr == 8'hc9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1217 = _T_1216 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1219 = btb_wr_addr == 8'hca; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1220 = _T_1219 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1222 = btb_wr_addr == 8'hcb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1223 = _T_1222 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1225 = btb_wr_addr == 8'hcc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1226 = _T_1225 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1228 = btb_wr_addr == 8'hcd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1229 = _T_1228 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1231 = btb_wr_addr == 8'hce; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1232 = _T_1231 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1234 = btb_wr_addr == 8'hcf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1235 = _T_1234 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1237 = btb_wr_addr == 8'hd0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1238 = _T_1237 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1240 = btb_wr_addr == 8'hd1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1241 = _T_1240 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1243 = btb_wr_addr == 8'hd2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1244 = _T_1243 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1246 = btb_wr_addr == 8'hd3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1247 = _T_1246 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1249 = btb_wr_addr == 8'hd4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1250 = _T_1249 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1252 = btb_wr_addr == 8'hd5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1253 = _T_1252 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1255 = btb_wr_addr == 8'hd6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1256 = _T_1255 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1258 = btb_wr_addr == 8'hd7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1259 = _T_1258 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1261 = btb_wr_addr == 8'hd8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1262 = _T_1261 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1264 = btb_wr_addr == 8'hd9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1265 = _T_1264 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1267 = btb_wr_addr == 8'hda; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1268 = _T_1267 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1270 = btb_wr_addr == 8'hdb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1271 = _T_1270 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1273 = btb_wr_addr == 8'hdc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1274 = _T_1273 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1276 = btb_wr_addr == 8'hdd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1277 = _T_1276 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1279 = btb_wr_addr == 8'hde; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1280 = _T_1279 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1282 = btb_wr_addr == 8'hdf; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1283 = _T_1282 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1285 = btb_wr_addr == 8'he0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1286 = _T_1285 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1288 = btb_wr_addr == 8'he1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1289 = _T_1288 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1291 = btb_wr_addr == 8'he2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1292 = _T_1291 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1294 = btb_wr_addr == 8'he3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1295 = _T_1294 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1297 = btb_wr_addr == 8'he4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1298 = _T_1297 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1300 = btb_wr_addr == 8'he5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1301 = _T_1300 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1303 = btb_wr_addr == 8'he6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1304 = _T_1303 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1306 = btb_wr_addr == 8'he7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1307 = _T_1306 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1309 = btb_wr_addr == 8'he8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1310 = _T_1309 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1312 = btb_wr_addr == 8'he9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1313 = _T_1312 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1315 = btb_wr_addr == 8'hea; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1316 = _T_1315 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1318 = btb_wr_addr == 8'heb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1319 = _T_1318 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1321 = btb_wr_addr == 8'hec; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1322 = _T_1321 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1324 = btb_wr_addr == 8'hed; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1325 = _T_1324 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1327 = btb_wr_addr == 8'hee; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1328 = _T_1327 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1330 = btb_wr_addr == 8'hef; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1331 = _T_1330 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1333 = btb_wr_addr == 8'hf0; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1334 = _T_1333 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1336 = btb_wr_addr == 8'hf1; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1337 = _T_1336 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1339 = btb_wr_addr == 8'hf2; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1340 = _T_1339 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1342 = btb_wr_addr == 8'hf3; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1343 = _T_1342 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1345 = btb_wr_addr == 8'hf4; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1346 = _T_1345 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1348 = btb_wr_addr == 8'hf5; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1349 = _T_1348 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1351 = btb_wr_addr == 8'hf6; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1352 = _T_1351 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1354 = btb_wr_addr == 8'hf7; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1355 = _T_1354 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1357 = btb_wr_addr == 8'hf8; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1358 = _T_1357 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1360 = btb_wr_addr == 8'hf9; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1361 = _T_1360 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1363 = btb_wr_addr == 8'hfa; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1364 = _T_1363 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1366 = btb_wr_addr == 8'hfb; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1367 = _T_1366 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1369 = btb_wr_addr == 8'hfc; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1370 = _T_1369 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1372 = btb_wr_addr == 8'hfd; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1373 = _T_1372 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1375 = btb_wr_addr == 8'hfe; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1376 = _T_1375 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1378 = btb_wr_addr == 8'hff; // @[ifu_bp_ctl.scala 432:98]
  wire  _T_1379 = _T_1378 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 432:107]
  wire  _T_1382 = _T_613 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1385 = _T_616 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1388 = _T_619 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1391 = _T_622 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1394 = _T_625 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1397 = _T_628 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1400 = _T_631 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1403 = _T_634 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1406 = _T_637 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1409 = _T_640 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1412 = _T_643 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1415 = _T_646 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1418 = _T_649 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1421 = _T_652 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1424 = _T_655 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1427 = _T_658 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1430 = _T_661 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1433 = _T_664 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1436 = _T_667 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1439 = _T_670 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1442 = _T_673 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1445 = _T_676 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1448 = _T_679 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1451 = _T_682 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1454 = _T_685 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1457 = _T_688 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1460 = _T_691 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1463 = _T_694 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1466 = _T_697 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1469 = _T_700 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1472 = _T_703 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1475 = _T_706 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1478 = _T_709 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1481 = _T_712 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1484 = _T_715 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1487 = _T_718 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1490 = _T_721 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1493 = _T_724 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1496 = _T_727 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1499 = _T_730 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1502 = _T_733 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1505 = _T_736 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1508 = _T_739 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1511 = _T_742 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1514 = _T_745 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1517 = _T_748 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1520 = _T_751 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1523 = _T_754 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1526 = _T_757 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1529 = _T_760 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1532 = _T_763 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1535 = _T_766 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1538 = _T_769 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1541 = _T_772 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1544 = _T_775 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1547 = _T_778 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1550 = _T_781 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1553 = _T_784 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1556 = _T_787 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1559 = _T_790 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1562 = _T_793 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1565 = _T_796 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1568 = _T_799 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1571 = _T_802 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1574 = _T_805 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1577 = _T_808 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1580 = _T_811 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1583 = _T_814 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1586 = _T_817 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1589 = _T_820 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1592 = _T_823 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1595 = _T_826 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1598 = _T_829 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1601 = _T_832 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1604 = _T_835 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1607 = _T_838 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1610 = _T_841 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1613 = _T_844 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1616 = _T_847 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1619 = _T_850 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1622 = _T_853 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1625 = _T_856 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1628 = _T_859 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1631 = _T_862 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1634 = _T_865 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1637 = _T_868 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1640 = _T_871 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1643 = _T_874 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1646 = _T_877 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1649 = _T_880 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1652 = _T_883 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1655 = _T_886 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1658 = _T_889 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1661 = _T_892 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1664 = _T_895 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1667 = _T_898 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1670 = _T_901 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1673 = _T_904 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1676 = _T_907 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1679 = _T_910 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1682 = _T_913 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1685 = _T_916 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1688 = _T_919 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1691 = _T_922 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1694 = _T_925 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1697 = _T_928 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1700 = _T_931 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1703 = _T_934 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1706 = _T_937 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1709 = _T_940 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1712 = _T_943 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1715 = _T_946 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1718 = _T_949 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1721 = _T_952 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1724 = _T_955 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1727 = _T_958 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1730 = _T_961 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1733 = _T_964 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1736 = _T_967 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1739 = _T_970 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1742 = _T_973 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1745 = _T_976 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1748 = _T_979 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1751 = _T_982 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1754 = _T_985 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1757 = _T_988 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1760 = _T_991 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1763 = _T_994 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1766 = _T_997 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1769 = _T_1000 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1772 = _T_1003 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1775 = _T_1006 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1778 = _T_1009 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1781 = _T_1012 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1784 = _T_1015 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1787 = _T_1018 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1790 = _T_1021 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1793 = _T_1024 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1796 = _T_1027 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1799 = _T_1030 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1802 = _T_1033 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1805 = _T_1036 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1808 = _T_1039 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1811 = _T_1042 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1814 = _T_1045 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1817 = _T_1048 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1820 = _T_1051 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1823 = _T_1054 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1826 = _T_1057 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1829 = _T_1060 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1832 = _T_1063 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1835 = _T_1066 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1838 = _T_1069 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1841 = _T_1072 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1844 = _T_1075 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1847 = _T_1078 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1850 = _T_1081 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1853 = _T_1084 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1856 = _T_1087 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1859 = _T_1090 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1862 = _T_1093 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1865 = _T_1096 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1868 = _T_1099 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1871 = _T_1102 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1874 = _T_1105 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1877 = _T_1108 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1880 = _T_1111 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1883 = _T_1114 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1886 = _T_1117 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1889 = _T_1120 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1892 = _T_1123 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1895 = _T_1126 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1898 = _T_1129 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1901 = _T_1132 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1904 = _T_1135 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1907 = _T_1138 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1910 = _T_1141 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1913 = _T_1144 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1916 = _T_1147 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1919 = _T_1150 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1922 = _T_1153 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1925 = _T_1156 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1928 = _T_1159 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1931 = _T_1162 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1934 = _T_1165 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1937 = _T_1168 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1940 = _T_1171 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1943 = _T_1174 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1946 = _T_1177 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1949 = _T_1180 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1952 = _T_1183 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1955 = _T_1186 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1958 = _T_1189 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1961 = _T_1192 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1964 = _T_1195 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1967 = _T_1198 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1970 = _T_1201 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1973 = _T_1204 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1976 = _T_1207 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1979 = _T_1210 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1982 = _T_1213 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1985 = _T_1216 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1988 = _T_1219 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1991 = _T_1222 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1994 = _T_1225 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_1997 = _T_1228 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2000 = _T_1231 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2003 = _T_1234 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2006 = _T_1237 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2009 = _T_1240 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2012 = _T_1243 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2015 = _T_1246 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2018 = _T_1249 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2021 = _T_1252 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2024 = _T_1255 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2027 = _T_1258 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2030 = _T_1261 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2033 = _T_1264 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2036 = _T_1267 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2039 = _T_1270 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2042 = _T_1273 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2045 = _T_1276 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2048 = _T_1279 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2051 = _T_1282 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2054 = _T_1285 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2057 = _T_1288 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2060 = _T_1291 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2063 = _T_1294 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2066 = _T_1297 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2069 = _T_1300 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2072 = _T_1303 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2075 = _T_1306 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2078 = _T_1309 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2081 = _T_1312 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2084 = _T_1315 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2087 = _T_1318 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2090 = _T_1321 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2093 = _T_1324 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2096 = _T_1327 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2099 = _T_1330 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2102 = _T_1333 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2105 = _T_1336 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2108 = _T_1339 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2111 = _T_1342 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2114 = _T_1345 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2117 = _T_1348 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2120 = _T_1351 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2123 = _T_1354 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2126 = _T_1357 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2129 = _T_1360 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2132 = _T_1363 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2135 = _T_1366 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2138 = _T_1369 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2141 = _T_1372 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2144 = _T_1375 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_2147 = _T_1378 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 433:107]
  wire  _T_6247 = mp_hashed[7:4] == 4'h0; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6249 = bht_wr_en0[0] & _T_6247; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6252 = br0_hashed_wb[7:4] == 4'h0; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6254 = bht_wr_en2[0] & _T_6252; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6258 = mp_hashed[7:4] == 4'h1; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6260 = bht_wr_en0[0] & _T_6258; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6263 = br0_hashed_wb[7:4] == 4'h1; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6265 = bht_wr_en2[0] & _T_6263; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6269 = mp_hashed[7:4] == 4'h2; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6271 = bht_wr_en0[0] & _T_6269; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6274 = br0_hashed_wb[7:4] == 4'h2; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6276 = bht_wr_en2[0] & _T_6274; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6280 = mp_hashed[7:4] == 4'h3; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6282 = bht_wr_en0[0] & _T_6280; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6285 = br0_hashed_wb[7:4] == 4'h3; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6287 = bht_wr_en2[0] & _T_6285; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6291 = mp_hashed[7:4] == 4'h4; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6293 = bht_wr_en0[0] & _T_6291; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6296 = br0_hashed_wb[7:4] == 4'h4; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6298 = bht_wr_en2[0] & _T_6296; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6302 = mp_hashed[7:4] == 4'h5; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6304 = bht_wr_en0[0] & _T_6302; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6307 = br0_hashed_wb[7:4] == 4'h5; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6309 = bht_wr_en2[0] & _T_6307; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6313 = mp_hashed[7:4] == 4'h6; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6315 = bht_wr_en0[0] & _T_6313; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6318 = br0_hashed_wb[7:4] == 4'h6; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6320 = bht_wr_en2[0] & _T_6318; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6324 = mp_hashed[7:4] == 4'h7; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6326 = bht_wr_en0[0] & _T_6324; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6329 = br0_hashed_wb[7:4] == 4'h7; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6331 = bht_wr_en2[0] & _T_6329; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6335 = mp_hashed[7:4] == 4'h8; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6337 = bht_wr_en0[0] & _T_6335; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6340 = br0_hashed_wb[7:4] == 4'h8; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6342 = bht_wr_en2[0] & _T_6340; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6346 = mp_hashed[7:4] == 4'h9; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6348 = bht_wr_en0[0] & _T_6346; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6351 = br0_hashed_wb[7:4] == 4'h9; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6353 = bht_wr_en2[0] & _T_6351; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6357 = mp_hashed[7:4] == 4'ha; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6359 = bht_wr_en0[0] & _T_6357; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6362 = br0_hashed_wb[7:4] == 4'ha; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6364 = bht_wr_en2[0] & _T_6362; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6368 = mp_hashed[7:4] == 4'hb; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6370 = bht_wr_en0[0] & _T_6368; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6373 = br0_hashed_wb[7:4] == 4'hb; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6375 = bht_wr_en2[0] & _T_6373; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6379 = mp_hashed[7:4] == 4'hc; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6381 = bht_wr_en0[0] & _T_6379; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6384 = br0_hashed_wb[7:4] == 4'hc; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6386 = bht_wr_en2[0] & _T_6384; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6390 = mp_hashed[7:4] == 4'hd; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6392 = bht_wr_en0[0] & _T_6390; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6395 = br0_hashed_wb[7:4] == 4'hd; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6397 = bht_wr_en2[0] & _T_6395; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6401 = mp_hashed[7:4] == 4'he; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6403 = bht_wr_en0[0] & _T_6401; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6406 = br0_hashed_wb[7:4] == 4'he; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6408 = bht_wr_en2[0] & _T_6406; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6412 = mp_hashed[7:4] == 4'hf; // @[ifu_bp_ctl.scala 512:109]
  wire  _T_6414 = bht_wr_en0[0] & _T_6412; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6417 = br0_hashed_wb[7:4] == 4'hf; // @[ifu_bp_ctl.scala 513:109]
  wire  _T_6419 = bht_wr_en2[0] & _T_6417; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6425 = bht_wr_en0[1] & _T_6247; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6430 = bht_wr_en2[1] & _T_6252; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6436 = bht_wr_en0[1] & _T_6258; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6441 = bht_wr_en2[1] & _T_6263; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6447 = bht_wr_en0[1] & _T_6269; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6452 = bht_wr_en2[1] & _T_6274; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6458 = bht_wr_en0[1] & _T_6280; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6463 = bht_wr_en2[1] & _T_6285; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6469 = bht_wr_en0[1] & _T_6291; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6474 = bht_wr_en2[1] & _T_6296; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6480 = bht_wr_en0[1] & _T_6302; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6485 = bht_wr_en2[1] & _T_6307; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6491 = bht_wr_en0[1] & _T_6313; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6496 = bht_wr_en2[1] & _T_6318; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6502 = bht_wr_en0[1] & _T_6324; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6507 = bht_wr_en2[1] & _T_6329; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6513 = bht_wr_en0[1] & _T_6335; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6518 = bht_wr_en2[1] & _T_6340; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6524 = bht_wr_en0[1] & _T_6346; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6529 = bht_wr_en2[1] & _T_6351; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6535 = bht_wr_en0[1] & _T_6357; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6540 = bht_wr_en2[1] & _T_6362; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6546 = bht_wr_en0[1] & _T_6368; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6551 = bht_wr_en2[1] & _T_6373; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6557 = bht_wr_en0[1] & _T_6379; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6562 = bht_wr_en2[1] & _T_6384; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6568 = bht_wr_en0[1] & _T_6390; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6573 = bht_wr_en2[1] & _T_6395; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6579 = bht_wr_en0[1] & _T_6401; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6584 = bht_wr_en2[1] & _T_6406; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6590 = bht_wr_en0[1] & _T_6412; // @[ifu_bp_ctl.scala 512:44]
  wire  _T_6595 = bht_wr_en2[1] & _T_6417; // @[ifu_bp_ctl.scala 513:44]
  wire  _T_6599 = br0_hashed_wb[3:0] == 4'h0; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6600 = bht_wr_en2[0] & _T_6599; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6604 = _T_6600 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6608 = br0_hashed_wb[3:0] == 4'h1; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6609 = bht_wr_en2[0] & _T_6608; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6613 = _T_6609 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6617 = br0_hashed_wb[3:0] == 4'h2; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6618 = bht_wr_en2[0] & _T_6617; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6622 = _T_6618 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6626 = br0_hashed_wb[3:0] == 4'h3; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6627 = bht_wr_en2[0] & _T_6626; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6631 = _T_6627 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6635 = br0_hashed_wb[3:0] == 4'h4; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6636 = bht_wr_en2[0] & _T_6635; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6640 = _T_6636 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6644 = br0_hashed_wb[3:0] == 4'h5; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6645 = bht_wr_en2[0] & _T_6644; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6649 = _T_6645 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6653 = br0_hashed_wb[3:0] == 4'h6; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6654 = bht_wr_en2[0] & _T_6653; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6658 = _T_6654 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6662 = br0_hashed_wb[3:0] == 4'h7; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6663 = bht_wr_en2[0] & _T_6662; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6667 = _T_6663 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6671 = br0_hashed_wb[3:0] == 4'h8; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6672 = bht_wr_en2[0] & _T_6671; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6676 = _T_6672 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6680 = br0_hashed_wb[3:0] == 4'h9; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6681 = bht_wr_en2[0] & _T_6680; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6685 = _T_6681 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6689 = br0_hashed_wb[3:0] == 4'ha; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6690 = bht_wr_en2[0] & _T_6689; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6694 = _T_6690 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6698 = br0_hashed_wb[3:0] == 4'hb; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6699 = bht_wr_en2[0] & _T_6698; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6703 = _T_6699 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6707 = br0_hashed_wb[3:0] == 4'hc; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6708 = bht_wr_en2[0] & _T_6707; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6712 = _T_6708 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6716 = br0_hashed_wb[3:0] == 4'hd; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6717 = bht_wr_en2[0] & _T_6716; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6721 = _T_6717 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6725 = br0_hashed_wb[3:0] == 4'he; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6726 = bht_wr_en2[0] & _T_6725; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6730 = _T_6726 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6734 = br0_hashed_wb[3:0] == 4'hf; // @[ifu_bp_ctl.scala 517:74]
  wire  _T_6735 = bht_wr_en2[0] & _T_6734; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_6739 = _T_6735 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6748 = _T_6600 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6757 = _T_6609 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6766 = _T_6618 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6775 = _T_6627 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6784 = _T_6636 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6793 = _T_6645 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6802 = _T_6654 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6811 = _T_6663 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6820 = _T_6672 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6829 = _T_6681 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6838 = _T_6690 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6847 = _T_6699 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6856 = _T_6708 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6865 = _T_6717 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6874 = _T_6726 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6883 = _T_6735 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6892 = _T_6600 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6901 = _T_6609 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6910 = _T_6618 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6919 = _T_6627 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6928 = _T_6636 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6937 = _T_6645 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6946 = _T_6654 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6955 = _T_6663 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6964 = _T_6672 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6973 = _T_6681 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6982 = _T_6690 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_6991 = _T_6699 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7000 = _T_6708 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7009 = _T_6717 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7018 = _T_6726 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7027 = _T_6735 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7036 = _T_6600 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7045 = _T_6609 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7054 = _T_6618 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7063 = _T_6627 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7072 = _T_6636 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7081 = _T_6645 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7090 = _T_6654 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7099 = _T_6663 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7108 = _T_6672 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7117 = _T_6681 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7126 = _T_6690 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7135 = _T_6699 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7144 = _T_6708 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7153 = _T_6717 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7162 = _T_6726 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7171 = _T_6735 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7180 = _T_6600 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7189 = _T_6609 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7198 = _T_6618 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7207 = _T_6627 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7216 = _T_6636 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7225 = _T_6645 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7234 = _T_6654 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7243 = _T_6663 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7252 = _T_6672 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7261 = _T_6681 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7270 = _T_6690 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7279 = _T_6699 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7288 = _T_6708 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7297 = _T_6717 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7306 = _T_6726 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7315 = _T_6735 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7324 = _T_6600 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7333 = _T_6609 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7342 = _T_6618 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7351 = _T_6627 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7360 = _T_6636 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7369 = _T_6645 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7378 = _T_6654 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7387 = _T_6663 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7396 = _T_6672 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7405 = _T_6681 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7414 = _T_6690 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7423 = _T_6699 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7432 = _T_6708 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7441 = _T_6717 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7450 = _T_6726 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7459 = _T_6735 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7468 = _T_6600 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7477 = _T_6609 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7486 = _T_6618 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7495 = _T_6627 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7504 = _T_6636 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7513 = _T_6645 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7522 = _T_6654 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7531 = _T_6663 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7540 = _T_6672 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7549 = _T_6681 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7558 = _T_6690 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7567 = _T_6699 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7576 = _T_6708 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7585 = _T_6717 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7594 = _T_6726 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7603 = _T_6735 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7612 = _T_6600 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7621 = _T_6609 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7630 = _T_6618 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7639 = _T_6627 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7648 = _T_6636 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7657 = _T_6645 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7666 = _T_6654 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7675 = _T_6663 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7684 = _T_6672 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7693 = _T_6681 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7702 = _T_6690 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7711 = _T_6699 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7720 = _T_6708 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7729 = _T_6717 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7738 = _T_6726 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7747 = _T_6735 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7756 = _T_6600 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7765 = _T_6609 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7774 = _T_6618 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7783 = _T_6627 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7792 = _T_6636 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7801 = _T_6645 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7810 = _T_6654 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7819 = _T_6663 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7828 = _T_6672 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7837 = _T_6681 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7846 = _T_6690 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7855 = _T_6699 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7864 = _T_6708 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7873 = _T_6717 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7882 = _T_6726 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7891 = _T_6735 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7900 = _T_6600 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7909 = _T_6609 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7918 = _T_6618 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7927 = _T_6627 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7936 = _T_6636 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7945 = _T_6645 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7954 = _T_6654 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7963 = _T_6663 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7972 = _T_6672 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7981 = _T_6681 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7990 = _T_6690 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_7999 = _T_6699 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8008 = _T_6708 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8017 = _T_6717 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8026 = _T_6726 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8035 = _T_6735 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8044 = _T_6600 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8053 = _T_6609 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8062 = _T_6618 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8071 = _T_6627 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8080 = _T_6636 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8089 = _T_6645 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8098 = _T_6654 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8107 = _T_6663 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8116 = _T_6672 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8125 = _T_6681 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8134 = _T_6690 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8143 = _T_6699 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8152 = _T_6708 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8161 = _T_6717 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8170 = _T_6726 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8179 = _T_6735 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8188 = _T_6600 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8197 = _T_6609 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8206 = _T_6618 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8215 = _T_6627 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8224 = _T_6636 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8233 = _T_6645 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8242 = _T_6654 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8251 = _T_6663 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8260 = _T_6672 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8269 = _T_6681 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8278 = _T_6690 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8287 = _T_6699 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8296 = _T_6708 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8305 = _T_6717 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8314 = _T_6726 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8323 = _T_6735 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8332 = _T_6600 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8341 = _T_6609 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8350 = _T_6618 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8359 = _T_6627 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8368 = _T_6636 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8377 = _T_6645 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8386 = _T_6654 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8395 = _T_6663 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8404 = _T_6672 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8413 = _T_6681 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8422 = _T_6690 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8431 = _T_6699 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8440 = _T_6708 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8449 = _T_6717 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8458 = _T_6726 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8467 = _T_6735 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8476 = _T_6600 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8485 = _T_6609 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8494 = _T_6618 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8503 = _T_6627 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8512 = _T_6636 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8521 = _T_6645 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8530 = _T_6654 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8539 = _T_6663 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8548 = _T_6672 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8557 = _T_6681 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8566 = _T_6690 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8575 = _T_6699 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8584 = _T_6708 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8593 = _T_6717 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8602 = _T_6726 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8611 = _T_6735 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8620 = _T_6600 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8629 = _T_6609 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8638 = _T_6618 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8647 = _T_6627 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8656 = _T_6636 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8665 = _T_6645 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8674 = _T_6654 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8683 = _T_6663 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8692 = _T_6672 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8701 = _T_6681 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8710 = _T_6690 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8719 = _T_6699 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8728 = _T_6708 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8737 = _T_6717 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8746 = _T_6726 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8755 = _T_6735 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8764 = _T_6600 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8773 = _T_6609 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8782 = _T_6618 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8791 = _T_6627 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8800 = _T_6636 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8809 = _T_6645 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8818 = _T_6654 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8827 = _T_6663 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8836 = _T_6672 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8845 = _T_6681 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8854 = _T_6690 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8863 = _T_6699 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8872 = _T_6708 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8881 = _T_6717 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8890 = _T_6726 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8899 = _T_6735 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8904 = bht_wr_en2[1] & _T_6599; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8908 = _T_8904 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8913 = bht_wr_en2[1] & _T_6608; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8917 = _T_8913 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8922 = bht_wr_en2[1] & _T_6617; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8926 = _T_8922 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8931 = bht_wr_en2[1] & _T_6626; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8935 = _T_8931 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8940 = bht_wr_en2[1] & _T_6635; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8944 = _T_8940 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8949 = bht_wr_en2[1] & _T_6644; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8953 = _T_8949 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8958 = bht_wr_en2[1] & _T_6653; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8962 = _T_8958 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8967 = bht_wr_en2[1] & _T_6662; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8971 = _T_8967 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8976 = bht_wr_en2[1] & _T_6671; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8980 = _T_8976 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8985 = bht_wr_en2[1] & _T_6680; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8989 = _T_8985 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_8994 = bht_wr_en2[1] & _T_6689; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_8998 = _T_8994 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9003 = bht_wr_en2[1] & _T_6698; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9007 = _T_9003 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9012 = bht_wr_en2[1] & _T_6707; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9016 = _T_9012 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9021 = bht_wr_en2[1] & _T_6716; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9025 = _T_9021 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9030 = bht_wr_en2[1] & _T_6725; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9034 = _T_9030 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9039 = bht_wr_en2[1] & _T_6734; // @[ifu_bp_ctl.scala 517:23]
  wire  _T_9043 = _T_9039 & _T_6252; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9052 = _T_8904 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9061 = _T_8913 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9070 = _T_8922 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9079 = _T_8931 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9088 = _T_8940 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9097 = _T_8949 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9106 = _T_8958 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9115 = _T_8967 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9124 = _T_8976 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9133 = _T_8985 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9142 = _T_8994 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9151 = _T_9003 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9160 = _T_9012 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9169 = _T_9021 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9178 = _T_9030 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9187 = _T_9039 & _T_6263; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9196 = _T_8904 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9205 = _T_8913 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9214 = _T_8922 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9223 = _T_8931 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9232 = _T_8940 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9241 = _T_8949 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9250 = _T_8958 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9259 = _T_8967 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9268 = _T_8976 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9277 = _T_8985 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9286 = _T_8994 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9295 = _T_9003 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9304 = _T_9012 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9313 = _T_9021 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9322 = _T_9030 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9331 = _T_9039 & _T_6274; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9340 = _T_8904 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9349 = _T_8913 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9358 = _T_8922 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9367 = _T_8931 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9376 = _T_8940 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9385 = _T_8949 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9394 = _T_8958 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9403 = _T_8967 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9412 = _T_8976 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9421 = _T_8985 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9430 = _T_8994 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9439 = _T_9003 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9448 = _T_9012 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9457 = _T_9021 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9466 = _T_9030 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9475 = _T_9039 & _T_6285; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9484 = _T_8904 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9493 = _T_8913 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9502 = _T_8922 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9511 = _T_8931 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9520 = _T_8940 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9529 = _T_8949 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9538 = _T_8958 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9547 = _T_8967 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9556 = _T_8976 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9565 = _T_8985 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9574 = _T_8994 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9583 = _T_9003 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9592 = _T_9012 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9601 = _T_9021 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9610 = _T_9030 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9619 = _T_9039 & _T_6296; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9628 = _T_8904 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9637 = _T_8913 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9646 = _T_8922 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9655 = _T_8931 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9664 = _T_8940 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9673 = _T_8949 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9682 = _T_8958 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9691 = _T_8967 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9700 = _T_8976 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9709 = _T_8985 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9718 = _T_8994 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9727 = _T_9003 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9736 = _T_9012 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9745 = _T_9021 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9754 = _T_9030 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9763 = _T_9039 & _T_6307; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9772 = _T_8904 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9781 = _T_8913 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9790 = _T_8922 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9799 = _T_8931 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9808 = _T_8940 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9817 = _T_8949 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9826 = _T_8958 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9835 = _T_8967 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9844 = _T_8976 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9853 = _T_8985 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9862 = _T_8994 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9871 = _T_9003 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9880 = _T_9012 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9889 = _T_9021 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9898 = _T_9030 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9907 = _T_9039 & _T_6318; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9916 = _T_8904 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9925 = _T_8913 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9934 = _T_8922 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9943 = _T_8931 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9952 = _T_8940 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9961 = _T_8949 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9970 = _T_8958 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9979 = _T_8967 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9988 = _T_8976 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_9997 = _T_8985 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10006 = _T_8994 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10015 = _T_9003 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10024 = _T_9012 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10033 = _T_9021 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10042 = _T_9030 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10051 = _T_9039 & _T_6329; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10060 = _T_8904 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10069 = _T_8913 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10078 = _T_8922 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10087 = _T_8931 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10096 = _T_8940 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10105 = _T_8949 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10114 = _T_8958 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10123 = _T_8967 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10132 = _T_8976 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10141 = _T_8985 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10150 = _T_8994 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10159 = _T_9003 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10168 = _T_9012 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10177 = _T_9021 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10186 = _T_9030 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10195 = _T_9039 & _T_6340; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10204 = _T_8904 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10213 = _T_8913 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10222 = _T_8922 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10231 = _T_8931 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10240 = _T_8940 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10249 = _T_8949 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10258 = _T_8958 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10267 = _T_8967 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10276 = _T_8976 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10285 = _T_8985 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10294 = _T_8994 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10303 = _T_9003 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10312 = _T_9012 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10321 = _T_9021 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10330 = _T_9030 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10339 = _T_9039 & _T_6351; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10348 = _T_8904 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10357 = _T_8913 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10366 = _T_8922 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10375 = _T_8931 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10384 = _T_8940 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10393 = _T_8949 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10402 = _T_8958 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10411 = _T_8967 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10420 = _T_8976 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10429 = _T_8985 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10438 = _T_8994 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10447 = _T_9003 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10456 = _T_9012 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10465 = _T_9021 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10474 = _T_9030 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10483 = _T_9039 & _T_6362; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10492 = _T_8904 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10501 = _T_8913 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10510 = _T_8922 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10519 = _T_8931 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10528 = _T_8940 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10537 = _T_8949 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10546 = _T_8958 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10555 = _T_8967 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10564 = _T_8976 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10573 = _T_8985 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10582 = _T_8994 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10591 = _T_9003 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10600 = _T_9012 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10609 = _T_9021 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10618 = _T_9030 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10627 = _T_9039 & _T_6373; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10636 = _T_8904 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10645 = _T_8913 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10654 = _T_8922 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10663 = _T_8931 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10672 = _T_8940 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10681 = _T_8949 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10690 = _T_8958 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10699 = _T_8967 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10708 = _T_8976 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10717 = _T_8985 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10726 = _T_8994 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10735 = _T_9003 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10744 = _T_9012 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10753 = _T_9021 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10762 = _T_9030 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10771 = _T_9039 & _T_6384; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10780 = _T_8904 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10789 = _T_8913 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10798 = _T_8922 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10807 = _T_8931 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10816 = _T_8940 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10825 = _T_8949 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10834 = _T_8958 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10843 = _T_8967 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10852 = _T_8976 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10861 = _T_8985 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10870 = _T_8994 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10879 = _T_9003 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10888 = _T_9012 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10897 = _T_9021 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10906 = _T_9030 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10915 = _T_9039 & _T_6395; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10924 = _T_8904 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10933 = _T_8913 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10942 = _T_8922 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10951 = _T_8931 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10960 = _T_8940 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10969 = _T_8949 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10978 = _T_8958 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10987 = _T_8967 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_10996 = _T_8976 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11005 = _T_8985 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11014 = _T_8994 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11023 = _T_9003 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11032 = _T_9012 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11041 = _T_9021 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11050 = _T_9030 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11059 = _T_9039 & _T_6406; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11068 = _T_8904 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11077 = _T_8913 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11086 = _T_8922 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11095 = _T_8931 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11104 = _T_8940 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11113 = _T_8949 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11122 = _T_8958 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11131 = _T_8967 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11140 = _T_8976 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11149 = _T_8985 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11158 = _T_8994 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11167 = _T_9003 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11176 = _T_9012 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11185 = _T_9021 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11194 = _T_9030 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11203 = _T_9039 & _T_6417; // @[ifu_bp_ctl.scala 517:81]
  wire  _T_11207 = mp_hashed[3:0] == 4'h0; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11208 = bht_wr_en0[0] & _T_11207; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11212 = _T_11208 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_0 = _T_11212 | _T_6604; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11224 = mp_hashed[3:0] == 4'h1; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11225 = bht_wr_en0[0] & _T_11224; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11229 = _T_11225 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_1 = _T_11229 | _T_6613; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11241 = mp_hashed[3:0] == 4'h2; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11242 = bht_wr_en0[0] & _T_11241; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11246 = _T_11242 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_2 = _T_11246 | _T_6622; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11258 = mp_hashed[3:0] == 4'h3; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11259 = bht_wr_en0[0] & _T_11258; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11263 = _T_11259 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_3 = _T_11263 | _T_6631; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11275 = mp_hashed[3:0] == 4'h4; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11276 = bht_wr_en0[0] & _T_11275; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11280 = _T_11276 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_4 = _T_11280 | _T_6640; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11292 = mp_hashed[3:0] == 4'h5; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11293 = bht_wr_en0[0] & _T_11292; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11297 = _T_11293 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_5 = _T_11297 | _T_6649; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11309 = mp_hashed[3:0] == 4'h6; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11310 = bht_wr_en0[0] & _T_11309; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11314 = _T_11310 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_6 = _T_11314 | _T_6658; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11326 = mp_hashed[3:0] == 4'h7; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11327 = bht_wr_en0[0] & _T_11326; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11331 = _T_11327 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_7 = _T_11331 | _T_6667; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11343 = mp_hashed[3:0] == 4'h8; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11344 = bht_wr_en0[0] & _T_11343; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11348 = _T_11344 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_8 = _T_11348 | _T_6676; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11360 = mp_hashed[3:0] == 4'h9; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11361 = bht_wr_en0[0] & _T_11360; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11365 = _T_11361 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_9 = _T_11365 | _T_6685; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11377 = mp_hashed[3:0] == 4'ha; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11378 = bht_wr_en0[0] & _T_11377; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11382 = _T_11378 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_10 = _T_11382 | _T_6694; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11394 = mp_hashed[3:0] == 4'hb; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11395 = bht_wr_en0[0] & _T_11394; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11399 = _T_11395 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_11 = _T_11399 | _T_6703; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11411 = mp_hashed[3:0] == 4'hc; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11412 = bht_wr_en0[0] & _T_11411; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11416 = _T_11412 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_12 = _T_11416 | _T_6712; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11428 = mp_hashed[3:0] == 4'hd; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11429 = bht_wr_en0[0] & _T_11428; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11433 = _T_11429 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_13 = _T_11433 | _T_6721; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11445 = mp_hashed[3:0] == 4'he; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11446 = bht_wr_en0[0] & _T_11445; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11450 = _T_11446 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_14 = _T_11450 | _T_6730; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11462 = mp_hashed[3:0] == 4'hf; // @[ifu_bp_ctl.scala 526:97]
  wire  _T_11463 = bht_wr_en0[0] & _T_11462; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_11467 = _T_11463 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_0_15 = _T_11467 | _T_6739; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11484 = _T_11208 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_0 = _T_11484 | _T_6748; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11501 = _T_11225 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_1 = _T_11501 | _T_6757; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11518 = _T_11242 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_2 = _T_11518 | _T_6766; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11535 = _T_11259 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_3 = _T_11535 | _T_6775; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11552 = _T_11276 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_4 = _T_11552 | _T_6784; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11569 = _T_11293 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_5 = _T_11569 | _T_6793; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11586 = _T_11310 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_6 = _T_11586 | _T_6802; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11603 = _T_11327 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_7 = _T_11603 | _T_6811; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11620 = _T_11344 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_8 = _T_11620 | _T_6820; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11637 = _T_11361 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_9 = _T_11637 | _T_6829; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11654 = _T_11378 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_10 = _T_11654 | _T_6838; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11671 = _T_11395 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_11 = _T_11671 | _T_6847; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11688 = _T_11412 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_12 = _T_11688 | _T_6856; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11705 = _T_11429 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_13 = _T_11705 | _T_6865; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11722 = _T_11446 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_14 = _T_11722 | _T_6874; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11739 = _T_11463 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_1_15 = _T_11739 | _T_6883; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11756 = _T_11208 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_0 = _T_11756 | _T_6892; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11773 = _T_11225 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_1 = _T_11773 | _T_6901; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11790 = _T_11242 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_2 = _T_11790 | _T_6910; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11807 = _T_11259 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_3 = _T_11807 | _T_6919; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11824 = _T_11276 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_4 = _T_11824 | _T_6928; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11841 = _T_11293 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_5 = _T_11841 | _T_6937; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11858 = _T_11310 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_6 = _T_11858 | _T_6946; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11875 = _T_11327 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_7 = _T_11875 | _T_6955; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11892 = _T_11344 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_8 = _T_11892 | _T_6964; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11909 = _T_11361 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_9 = _T_11909 | _T_6973; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11926 = _T_11378 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_10 = _T_11926 | _T_6982; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11943 = _T_11395 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_11 = _T_11943 | _T_6991; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11960 = _T_11412 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_12 = _T_11960 | _T_7000; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11977 = _T_11429 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_13 = _T_11977 | _T_7009; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_11994 = _T_11446 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_14 = _T_11994 | _T_7018; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12011 = _T_11463 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_2_15 = _T_12011 | _T_7027; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12028 = _T_11208 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_0 = _T_12028 | _T_7036; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12045 = _T_11225 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_1 = _T_12045 | _T_7045; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12062 = _T_11242 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_2 = _T_12062 | _T_7054; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12079 = _T_11259 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_3 = _T_12079 | _T_7063; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12096 = _T_11276 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_4 = _T_12096 | _T_7072; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12113 = _T_11293 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_5 = _T_12113 | _T_7081; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12130 = _T_11310 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_6 = _T_12130 | _T_7090; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12147 = _T_11327 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_7 = _T_12147 | _T_7099; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12164 = _T_11344 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_8 = _T_12164 | _T_7108; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12181 = _T_11361 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_9 = _T_12181 | _T_7117; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12198 = _T_11378 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_10 = _T_12198 | _T_7126; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12215 = _T_11395 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_11 = _T_12215 | _T_7135; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12232 = _T_11412 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_12 = _T_12232 | _T_7144; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12249 = _T_11429 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_13 = _T_12249 | _T_7153; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12266 = _T_11446 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_14 = _T_12266 | _T_7162; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12283 = _T_11463 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_3_15 = _T_12283 | _T_7171; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12300 = _T_11208 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_0 = _T_12300 | _T_7180; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12317 = _T_11225 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_1 = _T_12317 | _T_7189; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12334 = _T_11242 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_2 = _T_12334 | _T_7198; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12351 = _T_11259 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_3 = _T_12351 | _T_7207; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12368 = _T_11276 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_4 = _T_12368 | _T_7216; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12385 = _T_11293 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_5 = _T_12385 | _T_7225; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12402 = _T_11310 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_6 = _T_12402 | _T_7234; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12419 = _T_11327 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_7 = _T_12419 | _T_7243; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12436 = _T_11344 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_8 = _T_12436 | _T_7252; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12453 = _T_11361 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_9 = _T_12453 | _T_7261; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12470 = _T_11378 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_10 = _T_12470 | _T_7270; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12487 = _T_11395 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_11 = _T_12487 | _T_7279; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12504 = _T_11412 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_12 = _T_12504 | _T_7288; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12521 = _T_11429 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_13 = _T_12521 | _T_7297; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12538 = _T_11446 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_14 = _T_12538 | _T_7306; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12555 = _T_11463 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_4_15 = _T_12555 | _T_7315; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12572 = _T_11208 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_0 = _T_12572 | _T_7324; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12589 = _T_11225 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_1 = _T_12589 | _T_7333; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12606 = _T_11242 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_2 = _T_12606 | _T_7342; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12623 = _T_11259 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_3 = _T_12623 | _T_7351; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12640 = _T_11276 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_4 = _T_12640 | _T_7360; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12657 = _T_11293 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_5 = _T_12657 | _T_7369; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12674 = _T_11310 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_6 = _T_12674 | _T_7378; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12691 = _T_11327 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_7 = _T_12691 | _T_7387; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12708 = _T_11344 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_8 = _T_12708 | _T_7396; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12725 = _T_11361 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_9 = _T_12725 | _T_7405; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12742 = _T_11378 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_10 = _T_12742 | _T_7414; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12759 = _T_11395 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_11 = _T_12759 | _T_7423; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12776 = _T_11412 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_12 = _T_12776 | _T_7432; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12793 = _T_11429 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_13 = _T_12793 | _T_7441; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12810 = _T_11446 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_14 = _T_12810 | _T_7450; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12827 = _T_11463 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_5_15 = _T_12827 | _T_7459; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12844 = _T_11208 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_0 = _T_12844 | _T_7468; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12861 = _T_11225 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_1 = _T_12861 | _T_7477; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12878 = _T_11242 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_2 = _T_12878 | _T_7486; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12895 = _T_11259 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_3 = _T_12895 | _T_7495; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12912 = _T_11276 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_4 = _T_12912 | _T_7504; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12929 = _T_11293 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_5 = _T_12929 | _T_7513; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12946 = _T_11310 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_6 = _T_12946 | _T_7522; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12963 = _T_11327 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_7 = _T_12963 | _T_7531; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12980 = _T_11344 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_8 = _T_12980 | _T_7540; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_12997 = _T_11361 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_9 = _T_12997 | _T_7549; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13014 = _T_11378 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_10 = _T_13014 | _T_7558; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13031 = _T_11395 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_11 = _T_13031 | _T_7567; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13048 = _T_11412 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_12 = _T_13048 | _T_7576; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13065 = _T_11429 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_13 = _T_13065 | _T_7585; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13082 = _T_11446 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_14 = _T_13082 | _T_7594; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13099 = _T_11463 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_6_15 = _T_13099 | _T_7603; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13116 = _T_11208 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_0 = _T_13116 | _T_7612; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13133 = _T_11225 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_1 = _T_13133 | _T_7621; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13150 = _T_11242 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_2 = _T_13150 | _T_7630; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13167 = _T_11259 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_3 = _T_13167 | _T_7639; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13184 = _T_11276 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_4 = _T_13184 | _T_7648; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13201 = _T_11293 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_5 = _T_13201 | _T_7657; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13218 = _T_11310 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_6 = _T_13218 | _T_7666; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13235 = _T_11327 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_7 = _T_13235 | _T_7675; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13252 = _T_11344 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_8 = _T_13252 | _T_7684; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13269 = _T_11361 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_9 = _T_13269 | _T_7693; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13286 = _T_11378 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_10 = _T_13286 | _T_7702; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13303 = _T_11395 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_11 = _T_13303 | _T_7711; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13320 = _T_11412 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_12 = _T_13320 | _T_7720; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13337 = _T_11429 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_13 = _T_13337 | _T_7729; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13354 = _T_11446 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_14 = _T_13354 | _T_7738; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13371 = _T_11463 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_7_15 = _T_13371 | _T_7747; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13388 = _T_11208 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_0 = _T_13388 | _T_7756; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13405 = _T_11225 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_1 = _T_13405 | _T_7765; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13422 = _T_11242 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_2 = _T_13422 | _T_7774; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13439 = _T_11259 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_3 = _T_13439 | _T_7783; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13456 = _T_11276 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_4 = _T_13456 | _T_7792; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13473 = _T_11293 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_5 = _T_13473 | _T_7801; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13490 = _T_11310 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_6 = _T_13490 | _T_7810; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13507 = _T_11327 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_7 = _T_13507 | _T_7819; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13524 = _T_11344 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_8 = _T_13524 | _T_7828; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13541 = _T_11361 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_9 = _T_13541 | _T_7837; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13558 = _T_11378 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_10 = _T_13558 | _T_7846; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13575 = _T_11395 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_11 = _T_13575 | _T_7855; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13592 = _T_11412 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_12 = _T_13592 | _T_7864; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13609 = _T_11429 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_13 = _T_13609 | _T_7873; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13626 = _T_11446 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_14 = _T_13626 | _T_7882; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13643 = _T_11463 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_8_15 = _T_13643 | _T_7891; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13660 = _T_11208 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_0 = _T_13660 | _T_7900; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13677 = _T_11225 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_1 = _T_13677 | _T_7909; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13694 = _T_11242 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_2 = _T_13694 | _T_7918; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13711 = _T_11259 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_3 = _T_13711 | _T_7927; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13728 = _T_11276 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_4 = _T_13728 | _T_7936; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13745 = _T_11293 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_5 = _T_13745 | _T_7945; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13762 = _T_11310 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_6 = _T_13762 | _T_7954; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13779 = _T_11327 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_7 = _T_13779 | _T_7963; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13796 = _T_11344 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_8 = _T_13796 | _T_7972; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13813 = _T_11361 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_9 = _T_13813 | _T_7981; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13830 = _T_11378 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_10 = _T_13830 | _T_7990; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13847 = _T_11395 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_11 = _T_13847 | _T_7999; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13864 = _T_11412 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_12 = _T_13864 | _T_8008; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13881 = _T_11429 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_13 = _T_13881 | _T_8017; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13898 = _T_11446 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_14 = _T_13898 | _T_8026; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13915 = _T_11463 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_9_15 = _T_13915 | _T_8035; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13932 = _T_11208 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_0 = _T_13932 | _T_8044; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13949 = _T_11225 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_1 = _T_13949 | _T_8053; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13966 = _T_11242 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_2 = _T_13966 | _T_8062; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_13983 = _T_11259 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_3 = _T_13983 | _T_8071; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14000 = _T_11276 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_4 = _T_14000 | _T_8080; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14017 = _T_11293 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_5 = _T_14017 | _T_8089; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14034 = _T_11310 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_6 = _T_14034 | _T_8098; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14051 = _T_11327 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_7 = _T_14051 | _T_8107; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14068 = _T_11344 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_8 = _T_14068 | _T_8116; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14085 = _T_11361 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_9 = _T_14085 | _T_8125; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14102 = _T_11378 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_10 = _T_14102 | _T_8134; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14119 = _T_11395 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_11 = _T_14119 | _T_8143; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14136 = _T_11412 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_12 = _T_14136 | _T_8152; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14153 = _T_11429 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_13 = _T_14153 | _T_8161; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14170 = _T_11446 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_14 = _T_14170 | _T_8170; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14187 = _T_11463 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_10_15 = _T_14187 | _T_8179; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14204 = _T_11208 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_0 = _T_14204 | _T_8188; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14221 = _T_11225 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_1 = _T_14221 | _T_8197; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14238 = _T_11242 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_2 = _T_14238 | _T_8206; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14255 = _T_11259 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_3 = _T_14255 | _T_8215; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14272 = _T_11276 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_4 = _T_14272 | _T_8224; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14289 = _T_11293 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_5 = _T_14289 | _T_8233; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14306 = _T_11310 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_6 = _T_14306 | _T_8242; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14323 = _T_11327 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_7 = _T_14323 | _T_8251; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14340 = _T_11344 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_8 = _T_14340 | _T_8260; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14357 = _T_11361 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_9 = _T_14357 | _T_8269; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14374 = _T_11378 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_10 = _T_14374 | _T_8278; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14391 = _T_11395 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_11 = _T_14391 | _T_8287; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14408 = _T_11412 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_12 = _T_14408 | _T_8296; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14425 = _T_11429 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_13 = _T_14425 | _T_8305; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14442 = _T_11446 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_14 = _T_14442 | _T_8314; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14459 = _T_11463 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_11_15 = _T_14459 | _T_8323; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14476 = _T_11208 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_0 = _T_14476 | _T_8332; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14493 = _T_11225 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_1 = _T_14493 | _T_8341; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14510 = _T_11242 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_2 = _T_14510 | _T_8350; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14527 = _T_11259 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_3 = _T_14527 | _T_8359; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14544 = _T_11276 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_4 = _T_14544 | _T_8368; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14561 = _T_11293 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_5 = _T_14561 | _T_8377; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14578 = _T_11310 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_6 = _T_14578 | _T_8386; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14595 = _T_11327 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_7 = _T_14595 | _T_8395; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14612 = _T_11344 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_8 = _T_14612 | _T_8404; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14629 = _T_11361 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_9 = _T_14629 | _T_8413; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14646 = _T_11378 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_10 = _T_14646 | _T_8422; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14663 = _T_11395 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_11 = _T_14663 | _T_8431; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14680 = _T_11412 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_12 = _T_14680 | _T_8440; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14697 = _T_11429 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_13 = _T_14697 | _T_8449; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14714 = _T_11446 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_14 = _T_14714 | _T_8458; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14731 = _T_11463 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_12_15 = _T_14731 | _T_8467; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14748 = _T_11208 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_0 = _T_14748 | _T_8476; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14765 = _T_11225 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_1 = _T_14765 | _T_8485; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14782 = _T_11242 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_2 = _T_14782 | _T_8494; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14799 = _T_11259 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_3 = _T_14799 | _T_8503; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14816 = _T_11276 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_4 = _T_14816 | _T_8512; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14833 = _T_11293 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_5 = _T_14833 | _T_8521; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14850 = _T_11310 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_6 = _T_14850 | _T_8530; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14867 = _T_11327 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_7 = _T_14867 | _T_8539; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14884 = _T_11344 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_8 = _T_14884 | _T_8548; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14901 = _T_11361 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_9 = _T_14901 | _T_8557; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14918 = _T_11378 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_10 = _T_14918 | _T_8566; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14935 = _T_11395 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_11 = _T_14935 | _T_8575; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14952 = _T_11412 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_12 = _T_14952 | _T_8584; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14969 = _T_11429 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_13 = _T_14969 | _T_8593; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_14986 = _T_11446 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_14 = _T_14986 | _T_8602; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15003 = _T_11463 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_13_15 = _T_15003 | _T_8611; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15020 = _T_11208 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_0 = _T_15020 | _T_8620; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15037 = _T_11225 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_1 = _T_15037 | _T_8629; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15054 = _T_11242 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_2 = _T_15054 | _T_8638; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15071 = _T_11259 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_3 = _T_15071 | _T_8647; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15088 = _T_11276 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_4 = _T_15088 | _T_8656; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15105 = _T_11293 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_5 = _T_15105 | _T_8665; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15122 = _T_11310 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_6 = _T_15122 | _T_8674; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15139 = _T_11327 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_7 = _T_15139 | _T_8683; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15156 = _T_11344 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_8 = _T_15156 | _T_8692; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15173 = _T_11361 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_9 = _T_15173 | _T_8701; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15190 = _T_11378 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_10 = _T_15190 | _T_8710; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15207 = _T_11395 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_11 = _T_15207 | _T_8719; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15224 = _T_11412 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_12 = _T_15224 | _T_8728; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15241 = _T_11429 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_13 = _T_15241 | _T_8737; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15258 = _T_11446 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_14 = _T_15258 | _T_8746; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15275 = _T_11463 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_14_15 = _T_15275 | _T_8755; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15292 = _T_11208 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_0 = _T_15292 | _T_8764; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15309 = _T_11225 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_1 = _T_15309 | _T_8773; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15326 = _T_11242 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_2 = _T_15326 | _T_8782; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15343 = _T_11259 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_3 = _T_15343 | _T_8791; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15360 = _T_11276 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_4 = _T_15360 | _T_8800; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15377 = _T_11293 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_5 = _T_15377 | _T_8809; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15394 = _T_11310 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_6 = _T_15394 | _T_8818; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15411 = _T_11327 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_7 = _T_15411 | _T_8827; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15428 = _T_11344 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_8 = _T_15428 | _T_8836; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15445 = _T_11361 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_9 = _T_15445 | _T_8845; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15462 = _T_11378 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_10 = _T_15462 | _T_8854; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15479 = _T_11395 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_11 = _T_15479 | _T_8863; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15496 = _T_11412 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_12 = _T_15496 | _T_8872; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15513 = _T_11429 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_13 = _T_15513 | _T_8881; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15530 = _T_11446 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_14 = _T_15530 | _T_8890; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15547 = _T_11463 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_0_15_15 = _T_15547 | _T_8899; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15560 = bht_wr_en0[1] & _T_11207; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15564 = _T_15560 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_0 = _T_15564 | _T_8908; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15577 = bht_wr_en0[1] & _T_11224; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15581 = _T_15577 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_1 = _T_15581 | _T_8917; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15594 = bht_wr_en0[1] & _T_11241; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15598 = _T_15594 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_2 = _T_15598 | _T_8926; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15611 = bht_wr_en0[1] & _T_11258; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15615 = _T_15611 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_3 = _T_15615 | _T_8935; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15628 = bht_wr_en0[1] & _T_11275; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15632 = _T_15628 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_4 = _T_15632 | _T_8944; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15645 = bht_wr_en0[1] & _T_11292; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15649 = _T_15645 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_5 = _T_15649 | _T_8953; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15662 = bht_wr_en0[1] & _T_11309; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15666 = _T_15662 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_6 = _T_15666 | _T_8962; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15679 = bht_wr_en0[1] & _T_11326; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15683 = _T_15679 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_7 = _T_15683 | _T_8971; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15696 = bht_wr_en0[1] & _T_11343; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15700 = _T_15696 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_8 = _T_15700 | _T_8980; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15713 = bht_wr_en0[1] & _T_11360; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15717 = _T_15713 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_9 = _T_15717 | _T_8989; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15730 = bht_wr_en0[1] & _T_11377; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15734 = _T_15730 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_10 = _T_15734 | _T_8998; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15747 = bht_wr_en0[1] & _T_11394; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15751 = _T_15747 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_11 = _T_15751 | _T_9007; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15764 = bht_wr_en0[1] & _T_11411; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15768 = _T_15764 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_12 = _T_15768 | _T_9016; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15781 = bht_wr_en0[1] & _T_11428; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15785 = _T_15781 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_13 = _T_15785 | _T_9025; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15798 = bht_wr_en0[1] & _T_11445; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15802 = _T_15798 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_14 = _T_15802 | _T_9034; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15815 = bht_wr_en0[1] & _T_11462; // @[ifu_bp_ctl.scala 526:45]
  wire  _T_15819 = _T_15815 & _T_6247; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_0_15 = _T_15819 | _T_9043; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15836 = _T_15560 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_0 = _T_15836 | _T_9052; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15853 = _T_15577 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_1 = _T_15853 | _T_9061; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15870 = _T_15594 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_2 = _T_15870 | _T_9070; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15887 = _T_15611 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_3 = _T_15887 | _T_9079; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15904 = _T_15628 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_4 = _T_15904 | _T_9088; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15921 = _T_15645 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_5 = _T_15921 | _T_9097; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15938 = _T_15662 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_6 = _T_15938 | _T_9106; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15955 = _T_15679 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_7 = _T_15955 | _T_9115; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15972 = _T_15696 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_8 = _T_15972 | _T_9124; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_15989 = _T_15713 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_9 = _T_15989 | _T_9133; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16006 = _T_15730 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_10 = _T_16006 | _T_9142; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16023 = _T_15747 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_11 = _T_16023 | _T_9151; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16040 = _T_15764 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_12 = _T_16040 | _T_9160; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16057 = _T_15781 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_13 = _T_16057 | _T_9169; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16074 = _T_15798 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_14 = _T_16074 | _T_9178; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16091 = _T_15815 & _T_6258; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_1_15 = _T_16091 | _T_9187; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16108 = _T_15560 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_0 = _T_16108 | _T_9196; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16125 = _T_15577 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_1 = _T_16125 | _T_9205; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16142 = _T_15594 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_2 = _T_16142 | _T_9214; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16159 = _T_15611 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_3 = _T_16159 | _T_9223; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16176 = _T_15628 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_4 = _T_16176 | _T_9232; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16193 = _T_15645 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_5 = _T_16193 | _T_9241; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16210 = _T_15662 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_6 = _T_16210 | _T_9250; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16227 = _T_15679 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_7 = _T_16227 | _T_9259; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16244 = _T_15696 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_8 = _T_16244 | _T_9268; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16261 = _T_15713 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_9 = _T_16261 | _T_9277; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16278 = _T_15730 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_10 = _T_16278 | _T_9286; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16295 = _T_15747 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_11 = _T_16295 | _T_9295; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16312 = _T_15764 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_12 = _T_16312 | _T_9304; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16329 = _T_15781 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_13 = _T_16329 | _T_9313; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16346 = _T_15798 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_14 = _T_16346 | _T_9322; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16363 = _T_15815 & _T_6269; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_2_15 = _T_16363 | _T_9331; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16380 = _T_15560 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_0 = _T_16380 | _T_9340; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16397 = _T_15577 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_1 = _T_16397 | _T_9349; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16414 = _T_15594 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_2 = _T_16414 | _T_9358; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16431 = _T_15611 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_3 = _T_16431 | _T_9367; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16448 = _T_15628 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_4 = _T_16448 | _T_9376; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16465 = _T_15645 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_5 = _T_16465 | _T_9385; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16482 = _T_15662 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_6 = _T_16482 | _T_9394; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16499 = _T_15679 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_7 = _T_16499 | _T_9403; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16516 = _T_15696 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_8 = _T_16516 | _T_9412; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16533 = _T_15713 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_9 = _T_16533 | _T_9421; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16550 = _T_15730 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_10 = _T_16550 | _T_9430; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16567 = _T_15747 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_11 = _T_16567 | _T_9439; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16584 = _T_15764 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_12 = _T_16584 | _T_9448; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16601 = _T_15781 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_13 = _T_16601 | _T_9457; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16618 = _T_15798 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_14 = _T_16618 | _T_9466; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16635 = _T_15815 & _T_6280; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_3_15 = _T_16635 | _T_9475; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16652 = _T_15560 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_0 = _T_16652 | _T_9484; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16669 = _T_15577 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_1 = _T_16669 | _T_9493; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16686 = _T_15594 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_2 = _T_16686 | _T_9502; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16703 = _T_15611 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_3 = _T_16703 | _T_9511; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16720 = _T_15628 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_4 = _T_16720 | _T_9520; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16737 = _T_15645 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_5 = _T_16737 | _T_9529; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16754 = _T_15662 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_6 = _T_16754 | _T_9538; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16771 = _T_15679 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_7 = _T_16771 | _T_9547; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16788 = _T_15696 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_8 = _T_16788 | _T_9556; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16805 = _T_15713 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_9 = _T_16805 | _T_9565; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16822 = _T_15730 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_10 = _T_16822 | _T_9574; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16839 = _T_15747 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_11 = _T_16839 | _T_9583; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16856 = _T_15764 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_12 = _T_16856 | _T_9592; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16873 = _T_15781 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_13 = _T_16873 | _T_9601; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16890 = _T_15798 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_14 = _T_16890 | _T_9610; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16907 = _T_15815 & _T_6291; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_4_15 = _T_16907 | _T_9619; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16924 = _T_15560 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_0 = _T_16924 | _T_9628; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16941 = _T_15577 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_1 = _T_16941 | _T_9637; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16958 = _T_15594 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_2 = _T_16958 | _T_9646; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16975 = _T_15611 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_3 = _T_16975 | _T_9655; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_16992 = _T_15628 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_4 = _T_16992 | _T_9664; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17009 = _T_15645 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_5 = _T_17009 | _T_9673; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17026 = _T_15662 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_6 = _T_17026 | _T_9682; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17043 = _T_15679 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_7 = _T_17043 | _T_9691; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17060 = _T_15696 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_8 = _T_17060 | _T_9700; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17077 = _T_15713 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_9 = _T_17077 | _T_9709; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17094 = _T_15730 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_10 = _T_17094 | _T_9718; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17111 = _T_15747 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_11 = _T_17111 | _T_9727; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17128 = _T_15764 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_12 = _T_17128 | _T_9736; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17145 = _T_15781 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_13 = _T_17145 | _T_9745; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17162 = _T_15798 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_14 = _T_17162 | _T_9754; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17179 = _T_15815 & _T_6302; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_5_15 = _T_17179 | _T_9763; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17196 = _T_15560 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_0 = _T_17196 | _T_9772; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17213 = _T_15577 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_1 = _T_17213 | _T_9781; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17230 = _T_15594 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_2 = _T_17230 | _T_9790; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17247 = _T_15611 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_3 = _T_17247 | _T_9799; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17264 = _T_15628 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_4 = _T_17264 | _T_9808; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17281 = _T_15645 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_5 = _T_17281 | _T_9817; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17298 = _T_15662 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_6 = _T_17298 | _T_9826; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17315 = _T_15679 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_7 = _T_17315 | _T_9835; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17332 = _T_15696 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_8 = _T_17332 | _T_9844; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17349 = _T_15713 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_9 = _T_17349 | _T_9853; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17366 = _T_15730 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_10 = _T_17366 | _T_9862; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17383 = _T_15747 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_11 = _T_17383 | _T_9871; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17400 = _T_15764 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_12 = _T_17400 | _T_9880; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17417 = _T_15781 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_13 = _T_17417 | _T_9889; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17434 = _T_15798 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_14 = _T_17434 | _T_9898; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17451 = _T_15815 & _T_6313; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_6_15 = _T_17451 | _T_9907; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17468 = _T_15560 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_0 = _T_17468 | _T_9916; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17485 = _T_15577 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_1 = _T_17485 | _T_9925; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17502 = _T_15594 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_2 = _T_17502 | _T_9934; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17519 = _T_15611 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_3 = _T_17519 | _T_9943; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17536 = _T_15628 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_4 = _T_17536 | _T_9952; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17553 = _T_15645 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_5 = _T_17553 | _T_9961; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17570 = _T_15662 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_6 = _T_17570 | _T_9970; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17587 = _T_15679 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_7 = _T_17587 | _T_9979; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17604 = _T_15696 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_8 = _T_17604 | _T_9988; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17621 = _T_15713 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_9 = _T_17621 | _T_9997; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17638 = _T_15730 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_10 = _T_17638 | _T_10006; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17655 = _T_15747 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_11 = _T_17655 | _T_10015; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17672 = _T_15764 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_12 = _T_17672 | _T_10024; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17689 = _T_15781 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_13 = _T_17689 | _T_10033; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17706 = _T_15798 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_14 = _T_17706 | _T_10042; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17723 = _T_15815 & _T_6324; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_7_15 = _T_17723 | _T_10051; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17740 = _T_15560 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_0 = _T_17740 | _T_10060; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17757 = _T_15577 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_1 = _T_17757 | _T_10069; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17774 = _T_15594 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_2 = _T_17774 | _T_10078; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17791 = _T_15611 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_3 = _T_17791 | _T_10087; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17808 = _T_15628 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_4 = _T_17808 | _T_10096; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17825 = _T_15645 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_5 = _T_17825 | _T_10105; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17842 = _T_15662 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_6 = _T_17842 | _T_10114; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17859 = _T_15679 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_7 = _T_17859 | _T_10123; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17876 = _T_15696 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_8 = _T_17876 | _T_10132; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17893 = _T_15713 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_9 = _T_17893 | _T_10141; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17910 = _T_15730 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_10 = _T_17910 | _T_10150; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17927 = _T_15747 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_11 = _T_17927 | _T_10159; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17944 = _T_15764 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_12 = _T_17944 | _T_10168; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17961 = _T_15781 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_13 = _T_17961 | _T_10177; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17978 = _T_15798 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_14 = _T_17978 | _T_10186; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_17995 = _T_15815 & _T_6335; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_8_15 = _T_17995 | _T_10195; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18012 = _T_15560 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_0 = _T_18012 | _T_10204; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18029 = _T_15577 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_1 = _T_18029 | _T_10213; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18046 = _T_15594 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_2 = _T_18046 | _T_10222; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18063 = _T_15611 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_3 = _T_18063 | _T_10231; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18080 = _T_15628 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_4 = _T_18080 | _T_10240; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18097 = _T_15645 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_5 = _T_18097 | _T_10249; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18114 = _T_15662 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_6 = _T_18114 | _T_10258; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18131 = _T_15679 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_7 = _T_18131 | _T_10267; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18148 = _T_15696 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_8 = _T_18148 | _T_10276; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18165 = _T_15713 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_9 = _T_18165 | _T_10285; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18182 = _T_15730 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_10 = _T_18182 | _T_10294; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18199 = _T_15747 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_11 = _T_18199 | _T_10303; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18216 = _T_15764 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_12 = _T_18216 | _T_10312; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18233 = _T_15781 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_13 = _T_18233 | _T_10321; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18250 = _T_15798 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_14 = _T_18250 | _T_10330; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18267 = _T_15815 & _T_6346; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_9_15 = _T_18267 | _T_10339; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18284 = _T_15560 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_0 = _T_18284 | _T_10348; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18301 = _T_15577 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_1 = _T_18301 | _T_10357; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18318 = _T_15594 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_2 = _T_18318 | _T_10366; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18335 = _T_15611 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_3 = _T_18335 | _T_10375; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18352 = _T_15628 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_4 = _T_18352 | _T_10384; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18369 = _T_15645 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_5 = _T_18369 | _T_10393; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18386 = _T_15662 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_6 = _T_18386 | _T_10402; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18403 = _T_15679 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_7 = _T_18403 | _T_10411; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18420 = _T_15696 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_8 = _T_18420 | _T_10420; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18437 = _T_15713 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_9 = _T_18437 | _T_10429; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18454 = _T_15730 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_10 = _T_18454 | _T_10438; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18471 = _T_15747 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_11 = _T_18471 | _T_10447; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18488 = _T_15764 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_12 = _T_18488 | _T_10456; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18505 = _T_15781 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_13 = _T_18505 | _T_10465; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18522 = _T_15798 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_14 = _T_18522 | _T_10474; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18539 = _T_15815 & _T_6357; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_10_15 = _T_18539 | _T_10483; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18556 = _T_15560 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_0 = _T_18556 | _T_10492; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18573 = _T_15577 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_1 = _T_18573 | _T_10501; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18590 = _T_15594 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_2 = _T_18590 | _T_10510; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18607 = _T_15611 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_3 = _T_18607 | _T_10519; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18624 = _T_15628 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_4 = _T_18624 | _T_10528; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18641 = _T_15645 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_5 = _T_18641 | _T_10537; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18658 = _T_15662 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_6 = _T_18658 | _T_10546; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18675 = _T_15679 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_7 = _T_18675 | _T_10555; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18692 = _T_15696 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_8 = _T_18692 | _T_10564; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18709 = _T_15713 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_9 = _T_18709 | _T_10573; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18726 = _T_15730 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_10 = _T_18726 | _T_10582; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18743 = _T_15747 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_11 = _T_18743 | _T_10591; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18760 = _T_15764 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_12 = _T_18760 | _T_10600; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18777 = _T_15781 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_13 = _T_18777 | _T_10609; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18794 = _T_15798 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_14 = _T_18794 | _T_10618; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18811 = _T_15815 & _T_6368; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_11_15 = _T_18811 | _T_10627; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18828 = _T_15560 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_0 = _T_18828 | _T_10636; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18845 = _T_15577 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_1 = _T_18845 | _T_10645; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18862 = _T_15594 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_2 = _T_18862 | _T_10654; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18879 = _T_15611 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_3 = _T_18879 | _T_10663; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18896 = _T_15628 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_4 = _T_18896 | _T_10672; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18913 = _T_15645 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_5 = _T_18913 | _T_10681; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18930 = _T_15662 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_6 = _T_18930 | _T_10690; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18947 = _T_15679 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_7 = _T_18947 | _T_10699; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18964 = _T_15696 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_8 = _T_18964 | _T_10708; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18981 = _T_15713 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_9 = _T_18981 | _T_10717; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_18998 = _T_15730 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_10 = _T_18998 | _T_10726; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19015 = _T_15747 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_11 = _T_19015 | _T_10735; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19032 = _T_15764 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_12 = _T_19032 | _T_10744; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19049 = _T_15781 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_13 = _T_19049 | _T_10753; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19066 = _T_15798 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_14 = _T_19066 | _T_10762; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19083 = _T_15815 & _T_6379; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_12_15 = _T_19083 | _T_10771; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19100 = _T_15560 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_0 = _T_19100 | _T_10780; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19117 = _T_15577 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_1 = _T_19117 | _T_10789; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19134 = _T_15594 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_2 = _T_19134 | _T_10798; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19151 = _T_15611 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_3 = _T_19151 | _T_10807; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19168 = _T_15628 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_4 = _T_19168 | _T_10816; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19185 = _T_15645 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_5 = _T_19185 | _T_10825; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19202 = _T_15662 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_6 = _T_19202 | _T_10834; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19219 = _T_15679 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_7 = _T_19219 | _T_10843; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19236 = _T_15696 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_8 = _T_19236 | _T_10852; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19253 = _T_15713 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_9 = _T_19253 | _T_10861; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19270 = _T_15730 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_10 = _T_19270 | _T_10870; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19287 = _T_15747 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_11 = _T_19287 | _T_10879; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19304 = _T_15764 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_12 = _T_19304 | _T_10888; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19321 = _T_15781 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_13 = _T_19321 | _T_10897; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19338 = _T_15798 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_14 = _T_19338 | _T_10906; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19355 = _T_15815 & _T_6390; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_13_15 = _T_19355 | _T_10915; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19372 = _T_15560 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_0 = _T_19372 | _T_10924; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19389 = _T_15577 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_1 = _T_19389 | _T_10933; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19406 = _T_15594 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_2 = _T_19406 | _T_10942; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19423 = _T_15611 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_3 = _T_19423 | _T_10951; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19440 = _T_15628 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_4 = _T_19440 | _T_10960; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19457 = _T_15645 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_5 = _T_19457 | _T_10969; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19474 = _T_15662 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_6 = _T_19474 | _T_10978; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19491 = _T_15679 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_7 = _T_19491 | _T_10987; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19508 = _T_15696 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_8 = _T_19508 | _T_10996; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19525 = _T_15713 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_9 = _T_19525 | _T_11005; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19542 = _T_15730 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_10 = _T_19542 | _T_11014; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19559 = _T_15747 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_11 = _T_19559 | _T_11023; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19576 = _T_15764 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_12 = _T_19576 | _T_11032; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19593 = _T_15781 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_13 = _T_19593 | _T_11041; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19610 = _T_15798 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_14 = _T_19610 | _T_11050; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19627 = _T_15815 & _T_6401; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_14_15 = _T_19627 | _T_11059; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19644 = _T_15560 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_0 = _T_19644 | _T_11068; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19661 = _T_15577 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_1 = _T_19661 | _T_11077; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19678 = _T_15594 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_2 = _T_19678 | _T_11086; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19695 = _T_15611 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_3 = _T_19695 | _T_11095; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19712 = _T_15628 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_4 = _T_19712 | _T_11104; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19729 = _T_15645 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_5 = _T_19729 | _T_11113; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19746 = _T_15662 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_6 = _T_19746 | _T_11122; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19763 = _T_15679 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_7 = _T_19763 | _T_11131; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19780 = _T_15696 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_8 = _T_19780 | _T_11140; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19797 = _T_15713 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_9 = _T_19797 | _T_11149; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19814 = _T_15730 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_10 = _T_19814 | _T_11158; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19831 = _T_15747 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_11 = _T_19831 | _T_11167; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19848 = _T_15764 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_12 = _T_19848 | _T_11176; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19865 = _T_15781 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_13 = _T_19865 | _T_11185; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19882 = _T_15798 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_14 = _T_19882 | _T_11194; // @[ifu_bp_ctl.scala 526:223]
  wire  _T_19899 = _T_15815 & _T_6412; // @[ifu_bp_ctl.scala 526:110]
  wire  bht_bank_sel_1_15_15 = _T_19899 | _T_11203; // @[ifu_bp_ctl.scala 526:223]
  rvclkhdr rvclkhdr ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en)
  );
  rvclkhdr rvclkhdr_47 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en)
  );
  rvclkhdr rvclkhdr_48 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en)
  );
  rvclkhdr rvclkhdr_49 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en)
  );
  rvclkhdr rvclkhdr_50 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en)
  );
  rvclkhdr rvclkhdr_51 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en)
  );
  rvclkhdr rvclkhdr_52 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en)
  );
  rvclkhdr rvclkhdr_53 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en)
  );
  rvclkhdr rvclkhdr_54 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en)
  );
  rvclkhdr rvclkhdr_55 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en)
  );
  rvclkhdr rvclkhdr_56 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en)
  );
  rvclkhdr rvclkhdr_57 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en)
  );
  rvclkhdr rvclkhdr_58 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en)
  );
  rvclkhdr rvclkhdr_59 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en)
  );
  rvclkhdr rvclkhdr_60 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en)
  );
  rvclkhdr rvclkhdr_61 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en)
  );
  rvclkhdr rvclkhdr_62 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en)
  );
  rvclkhdr rvclkhdr_63 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en)
  );
  rvclkhdr rvclkhdr_64 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en)
  );
  rvclkhdr rvclkhdr_65 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en)
  );
  rvclkhdr rvclkhdr_66 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en)
  );
  rvclkhdr rvclkhdr_67 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en)
  );
  rvclkhdr rvclkhdr_68 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en)
  );
  rvclkhdr rvclkhdr_69 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en)
  );
  rvclkhdr rvclkhdr_70 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en)
  );
  rvclkhdr rvclkhdr_71 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en)
  );
  rvclkhdr rvclkhdr_72 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en)
  );
  rvclkhdr rvclkhdr_73 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en)
  );
  rvclkhdr rvclkhdr_74 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en)
  );
  rvclkhdr rvclkhdr_75 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en)
  );
  rvclkhdr rvclkhdr_76 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en)
  );
  rvclkhdr rvclkhdr_77 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en)
  );
  rvclkhdr rvclkhdr_78 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en)
  );
  rvclkhdr rvclkhdr_79 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en)
  );
  rvclkhdr rvclkhdr_80 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en)
  );
  rvclkhdr rvclkhdr_81 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en)
  );
  rvclkhdr rvclkhdr_82 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en)
  );
  rvclkhdr rvclkhdr_83 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en)
  );
  rvclkhdr rvclkhdr_84 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en)
  );
  rvclkhdr rvclkhdr_85 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en)
  );
  rvclkhdr rvclkhdr_86 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en)
  );
  rvclkhdr rvclkhdr_87 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en)
  );
  rvclkhdr rvclkhdr_88 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en)
  );
  rvclkhdr rvclkhdr_89 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en)
  );
  rvclkhdr rvclkhdr_90 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en)
  );
  rvclkhdr rvclkhdr_91 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en)
  );
  rvclkhdr rvclkhdr_92 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en)
  );
  rvclkhdr rvclkhdr_93 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en)
  );
  rvclkhdr rvclkhdr_94 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_94_io_clk),
    .io_en(rvclkhdr_94_io_en)
  );
  rvclkhdr rvclkhdr_95 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_95_io_clk),
    .io_en(rvclkhdr_95_io_en)
  );
  rvclkhdr rvclkhdr_96 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_96_io_clk),
    .io_en(rvclkhdr_96_io_en)
  );
  rvclkhdr rvclkhdr_97 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_97_io_clk),
    .io_en(rvclkhdr_97_io_en)
  );
  rvclkhdr rvclkhdr_98 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_98_io_clk),
    .io_en(rvclkhdr_98_io_en)
  );
  rvclkhdr rvclkhdr_99 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_99_io_clk),
    .io_en(rvclkhdr_99_io_en)
  );
  rvclkhdr rvclkhdr_100 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_100_io_clk),
    .io_en(rvclkhdr_100_io_en)
  );
  rvclkhdr rvclkhdr_101 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_101_io_clk),
    .io_en(rvclkhdr_101_io_en)
  );
  rvclkhdr rvclkhdr_102 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_102_io_clk),
    .io_en(rvclkhdr_102_io_en)
  );
  rvclkhdr rvclkhdr_103 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_103_io_clk),
    .io_en(rvclkhdr_103_io_en)
  );
  rvclkhdr rvclkhdr_104 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_104_io_clk),
    .io_en(rvclkhdr_104_io_en)
  );
  rvclkhdr rvclkhdr_105 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_105_io_clk),
    .io_en(rvclkhdr_105_io_en)
  );
  rvclkhdr rvclkhdr_106 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_106_io_clk),
    .io_en(rvclkhdr_106_io_en)
  );
  rvclkhdr rvclkhdr_107 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_107_io_clk),
    .io_en(rvclkhdr_107_io_en)
  );
  rvclkhdr rvclkhdr_108 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_108_io_clk),
    .io_en(rvclkhdr_108_io_en)
  );
  rvclkhdr rvclkhdr_109 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_109_io_clk),
    .io_en(rvclkhdr_109_io_en)
  );
  rvclkhdr rvclkhdr_110 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_110_io_clk),
    .io_en(rvclkhdr_110_io_en)
  );
  rvclkhdr rvclkhdr_111 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_111_io_clk),
    .io_en(rvclkhdr_111_io_en)
  );
  rvclkhdr rvclkhdr_112 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_112_io_clk),
    .io_en(rvclkhdr_112_io_en)
  );
  rvclkhdr rvclkhdr_113 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_113_io_clk),
    .io_en(rvclkhdr_113_io_en)
  );
  rvclkhdr rvclkhdr_114 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_114_io_clk),
    .io_en(rvclkhdr_114_io_en)
  );
  rvclkhdr rvclkhdr_115 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_115_io_clk),
    .io_en(rvclkhdr_115_io_en)
  );
  rvclkhdr rvclkhdr_116 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_116_io_clk),
    .io_en(rvclkhdr_116_io_en)
  );
  rvclkhdr rvclkhdr_117 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_117_io_clk),
    .io_en(rvclkhdr_117_io_en)
  );
  rvclkhdr rvclkhdr_118 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_118_io_clk),
    .io_en(rvclkhdr_118_io_en)
  );
  rvclkhdr rvclkhdr_119 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_119_io_clk),
    .io_en(rvclkhdr_119_io_en)
  );
  rvclkhdr rvclkhdr_120 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_120_io_clk),
    .io_en(rvclkhdr_120_io_en)
  );
  rvclkhdr rvclkhdr_121 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_121_io_clk),
    .io_en(rvclkhdr_121_io_en)
  );
  rvclkhdr rvclkhdr_122 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_122_io_clk),
    .io_en(rvclkhdr_122_io_en)
  );
  rvclkhdr rvclkhdr_123 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_123_io_clk),
    .io_en(rvclkhdr_123_io_en)
  );
  rvclkhdr rvclkhdr_124 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_124_io_clk),
    .io_en(rvclkhdr_124_io_en)
  );
  rvclkhdr rvclkhdr_125 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_125_io_clk),
    .io_en(rvclkhdr_125_io_en)
  );
  rvclkhdr rvclkhdr_126 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_126_io_clk),
    .io_en(rvclkhdr_126_io_en)
  );
  rvclkhdr rvclkhdr_127 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_127_io_clk),
    .io_en(rvclkhdr_127_io_en)
  );
  rvclkhdr rvclkhdr_128 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_128_io_clk),
    .io_en(rvclkhdr_128_io_en)
  );
  rvclkhdr rvclkhdr_129 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_129_io_clk),
    .io_en(rvclkhdr_129_io_en)
  );
  rvclkhdr rvclkhdr_130 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_130_io_clk),
    .io_en(rvclkhdr_130_io_en)
  );
  rvclkhdr rvclkhdr_131 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_131_io_clk),
    .io_en(rvclkhdr_131_io_en)
  );
  rvclkhdr rvclkhdr_132 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_132_io_clk),
    .io_en(rvclkhdr_132_io_en)
  );
  rvclkhdr rvclkhdr_133 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_133_io_clk),
    .io_en(rvclkhdr_133_io_en)
  );
  rvclkhdr rvclkhdr_134 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_134_io_clk),
    .io_en(rvclkhdr_134_io_en)
  );
  rvclkhdr rvclkhdr_135 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_135_io_clk),
    .io_en(rvclkhdr_135_io_en)
  );
  rvclkhdr rvclkhdr_136 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_136_io_clk),
    .io_en(rvclkhdr_136_io_en)
  );
  rvclkhdr rvclkhdr_137 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_137_io_clk),
    .io_en(rvclkhdr_137_io_en)
  );
  rvclkhdr rvclkhdr_138 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_138_io_clk),
    .io_en(rvclkhdr_138_io_en)
  );
  rvclkhdr rvclkhdr_139 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_139_io_clk),
    .io_en(rvclkhdr_139_io_en)
  );
  rvclkhdr rvclkhdr_140 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_140_io_clk),
    .io_en(rvclkhdr_140_io_en)
  );
  rvclkhdr rvclkhdr_141 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_141_io_clk),
    .io_en(rvclkhdr_141_io_en)
  );
  rvclkhdr rvclkhdr_142 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_142_io_clk),
    .io_en(rvclkhdr_142_io_en)
  );
  rvclkhdr rvclkhdr_143 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_143_io_clk),
    .io_en(rvclkhdr_143_io_en)
  );
  rvclkhdr rvclkhdr_144 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_144_io_clk),
    .io_en(rvclkhdr_144_io_en)
  );
  rvclkhdr rvclkhdr_145 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_145_io_clk),
    .io_en(rvclkhdr_145_io_en)
  );
  rvclkhdr rvclkhdr_146 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_146_io_clk),
    .io_en(rvclkhdr_146_io_en)
  );
  rvclkhdr rvclkhdr_147 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_147_io_clk),
    .io_en(rvclkhdr_147_io_en)
  );
  rvclkhdr rvclkhdr_148 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_148_io_clk),
    .io_en(rvclkhdr_148_io_en)
  );
  rvclkhdr rvclkhdr_149 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_149_io_clk),
    .io_en(rvclkhdr_149_io_en)
  );
  rvclkhdr rvclkhdr_150 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_150_io_clk),
    .io_en(rvclkhdr_150_io_en)
  );
  rvclkhdr rvclkhdr_151 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_151_io_clk),
    .io_en(rvclkhdr_151_io_en)
  );
  rvclkhdr rvclkhdr_152 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_152_io_clk),
    .io_en(rvclkhdr_152_io_en)
  );
  rvclkhdr rvclkhdr_153 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_153_io_clk),
    .io_en(rvclkhdr_153_io_en)
  );
  rvclkhdr rvclkhdr_154 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_154_io_clk),
    .io_en(rvclkhdr_154_io_en)
  );
  rvclkhdr rvclkhdr_155 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_155_io_clk),
    .io_en(rvclkhdr_155_io_en)
  );
  rvclkhdr rvclkhdr_156 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_156_io_clk),
    .io_en(rvclkhdr_156_io_en)
  );
  rvclkhdr rvclkhdr_157 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_157_io_clk),
    .io_en(rvclkhdr_157_io_en)
  );
  rvclkhdr rvclkhdr_158 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_158_io_clk),
    .io_en(rvclkhdr_158_io_en)
  );
  rvclkhdr rvclkhdr_159 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_159_io_clk),
    .io_en(rvclkhdr_159_io_en)
  );
  rvclkhdr rvclkhdr_160 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_160_io_clk),
    .io_en(rvclkhdr_160_io_en)
  );
  rvclkhdr rvclkhdr_161 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_161_io_clk),
    .io_en(rvclkhdr_161_io_en)
  );
  rvclkhdr rvclkhdr_162 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_162_io_clk),
    .io_en(rvclkhdr_162_io_en)
  );
  rvclkhdr rvclkhdr_163 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_163_io_clk),
    .io_en(rvclkhdr_163_io_en)
  );
  rvclkhdr rvclkhdr_164 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_164_io_clk),
    .io_en(rvclkhdr_164_io_en)
  );
  rvclkhdr rvclkhdr_165 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_165_io_clk),
    .io_en(rvclkhdr_165_io_en)
  );
  rvclkhdr rvclkhdr_166 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_166_io_clk),
    .io_en(rvclkhdr_166_io_en)
  );
  rvclkhdr rvclkhdr_167 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_167_io_clk),
    .io_en(rvclkhdr_167_io_en)
  );
  rvclkhdr rvclkhdr_168 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_168_io_clk),
    .io_en(rvclkhdr_168_io_en)
  );
  rvclkhdr rvclkhdr_169 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_169_io_clk),
    .io_en(rvclkhdr_169_io_en)
  );
  rvclkhdr rvclkhdr_170 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_170_io_clk),
    .io_en(rvclkhdr_170_io_en)
  );
  rvclkhdr rvclkhdr_171 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_171_io_clk),
    .io_en(rvclkhdr_171_io_en)
  );
  rvclkhdr rvclkhdr_172 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_172_io_clk),
    .io_en(rvclkhdr_172_io_en)
  );
  rvclkhdr rvclkhdr_173 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_173_io_clk),
    .io_en(rvclkhdr_173_io_en)
  );
  rvclkhdr rvclkhdr_174 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_174_io_clk),
    .io_en(rvclkhdr_174_io_en)
  );
  rvclkhdr rvclkhdr_175 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_175_io_clk),
    .io_en(rvclkhdr_175_io_en)
  );
  rvclkhdr rvclkhdr_176 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_176_io_clk),
    .io_en(rvclkhdr_176_io_en)
  );
  rvclkhdr rvclkhdr_177 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_177_io_clk),
    .io_en(rvclkhdr_177_io_en)
  );
  rvclkhdr rvclkhdr_178 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_178_io_clk),
    .io_en(rvclkhdr_178_io_en)
  );
  rvclkhdr rvclkhdr_179 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_179_io_clk),
    .io_en(rvclkhdr_179_io_en)
  );
  rvclkhdr rvclkhdr_180 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_180_io_clk),
    .io_en(rvclkhdr_180_io_en)
  );
  rvclkhdr rvclkhdr_181 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_181_io_clk),
    .io_en(rvclkhdr_181_io_en)
  );
  rvclkhdr rvclkhdr_182 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_182_io_clk),
    .io_en(rvclkhdr_182_io_en)
  );
  rvclkhdr rvclkhdr_183 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_183_io_clk),
    .io_en(rvclkhdr_183_io_en)
  );
  rvclkhdr rvclkhdr_184 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_184_io_clk),
    .io_en(rvclkhdr_184_io_en)
  );
  rvclkhdr rvclkhdr_185 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_185_io_clk),
    .io_en(rvclkhdr_185_io_en)
  );
  rvclkhdr rvclkhdr_186 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_186_io_clk),
    .io_en(rvclkhdr_186_io_en)
  );
  rvclkhdr rvclkhdr_187 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_187_io_clk),
    .io_en(rvclkhdr_187_io_en)
  );
  rvclkhdr rvclkhdr_188 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_188_io_clk),
    .io_en(rvclkhdr_188_io_en)
  );
  rvclkhdr rvclkhdr_189 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_189_io_clk),
    .io_en(rvclkhdr_189_io_en)
  );
  rvclkhdr rvclkhdr_190 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_190_io_clk),
    .io_en(rvclkhdr_190_io_en)
  );
  rvclkhdr rvclkhdr_191 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_191_io_clk),
    .io_en(rvclkhdr_191_io_en)
  );
  rvclkhdr rvclkhdr_192 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_192_io_clk),
    .io_en(rvclkhdr_192_io_en)
  );
  rvclkhdr rvclkhdr_193 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_193_io_clk),
    .io_en(rvclkhdr_193_io_en)
  );
  rvclkhdr rvclkhdr_194 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_194_io_clk),
    .io_en(rvclkhdr_194_io_en)
  );
  rvclkhdr rvclkhdr_195 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_195_io_clk),
    .io_en(rvclkhdr_195_io_en)
  );
  rvclkhdr rvclkhdr_196 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_196_io_clk),
    .io_en(rvclkhdr_196_io_en)
  );
  rvclkhdr rvclkhdr_197 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_197_io_clk),
    .io_en(rvclkhdr_197_io_en)
  );
  rvclkhdr rvclkhdr_198 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_198_io_clk),
    .io_en(rvclkhdr_198_io_en)
  );
  rvclkhdr rvclkhdr_199 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_199_io_clk),
    .io_en(rvclkhdr_199_io_en)
  );
  rvclkhdr rvclkhdr_200 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_200_io_clk),
    .io_en(rvclkhdr_200_io_en)
  );
  rvclkhdr rvclkhdr_201 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_201_io_clk),
    .io_en(rvclkhdr_201_io_en)
  );
  rvclkhdr rvclkhdr_202 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_202_io_clk),
    .io_en(rvclkhdr_202_io_en)
  );
  rvclkhdr rvclkhdr_203 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_203_io_clk),
    .io_en(rvclkhdr_203_io_en)
  );
  rvclkhdr rvclkhdr_204 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_204_io_clk),
    .io_en(rvclkhdr_204_io_en)
  );
  rvclkhdr rvclkhdr_205 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_205_io_clk),
    .io_en(rvclkhdr_205_io_en)
  );
  rvclkhdr rvclkhdr_206 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_206_io_clk),
    .io_en(rvclkhdr_206_io_en)
  );
  rvclkhdr rvclkhdr_207 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_207_io_clk),
    .io_en(rvclkhdr_207_io_en)
  );
  rvclkhdr rvclkhdr_208 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_208_io_clk),
    .io_en(rvclkhdr_208_io_en)
  );
  rvclkhdr rvclkhdr_209 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_209_io_clk),
    .io_en(rvclkhdr_209_io_en)
  );
  rvclkhdr rvclkhdr_210 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_210_io_clk),
    .io_en(rvclkhdr_210_io_en)
  );
  rvclkhdr rvclkhdr_211 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_211_io_clk),
    .io_en(rvclkhdr_211_io_en)
  );
  rvclkhdr rvclkhdr_212 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_212_io_clk),
    .io_en(rvclkhdr_212_io_en)
  );
  rvclkhdr rvclkhdr_213 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_213_io_clk),
    .io_en(rvclkhdr_213_io_en)
  );
  rvclkhdr rvclkhdr_214 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_214_io_clk),
    .io_en(rvclkhdr_214_io_en)
  );
  rvclkhdr rvclkhdr_215 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_215_io_clk),
    .io_en(rvclkhdr_215_io_en)
  );
  rvclkhdr rvclkhdr_216 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_216_io_clk),
    .io_en(rvclkhdr_216_io_en)
  );
  rvclkhdr rvclkhdr_217 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_217_io_clk),
    .io_en(rvclkhdr_217_io_en)
  );
  rvclkhdr rvclkhdr_218 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_218_io_clk),
    .io_en(rvclkhdr_218_io_en)
  );
  rvclkhdr rvclkhdr_219 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_219_io_clk),
    .io_en(rvclkhdr_219_io_en)
  );
  rvclkhdr rvclkhdr_220 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_220_io_clk),
    .io_en(rvclkhdr_220_io_en)
  );
  rvclkhdr rvclkhdr_221 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_221_io_clk),
    .io_en(rvclkhdr_221_io_en)
  );
  rvclkhdr rvclkhdr_222 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_222_io_clk),
    .io_en(rvclkhdr_222_io_en)
  );
  rvclkhdr rvclkhdr_223 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_223_io_clk),
    .io_en(rvclkhdr_223_io_en)
  );
  rvclkhdr rvclkhdr_224 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_224_io_clk),
    .io_en(rvclkhdr_224_io_en)
  );
  rvclkhdr rvclkhdr_225 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_225_io_clk),
    .io_en(rvclkhdr_225_io_en)
  );
  rvclkhdr rvclkhdr_226 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_226_io_clk),
    .io_en(rvclkhdr_226_io_en)
  );
  rvclkhdr rvclkhdr_227 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_227_io_clk),
    .io_en(rvclkhdr_227_io_en)
  );
  rvclkhdr rvclkhdr_228 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_228_io_clk),
    .io_en(rvclkhdr_228_io_en)
  );
  rvclkhdr rvclkhdr_229 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_229_io_clk),
    .io_en(rvclkhdr_229_io_en)
  );
  rvclkhdr rvclkhdr_230 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_230_io_clk),
    .io_en(rvclkhdr_230_io_en)
  );
  rvclkhdr rvclkhdr_231 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_231_io_clk),
    .io_en(rvclkhdr_231_io_en)
  );
  rvclkhdr rvclkhdr_232 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_232_io_clk),
    .io_en(rvclkhdr_232_io_en)
  );
  rvclkhdr rvclkhdr_233 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_233_io_clk),
    .io_en(rvclkhdr_233_io_en)
  );
  rvclkhdr rvclkhdr_234 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_234_io_clk),
    .io_en(rvclkhdr_234_io_en)
  );
  rvclkhdr rvclkhdr_235 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_235_io_clk),
    .io_en(rvclkhdr_235_io_en)
  );
  rvclkhdr rvclkhdr_236 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_236_io_clk),
    .io_en(rvclkhdr_236_io_en)
  );
  rvclkhdr rvclkhdr_237 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_237_io_clk),
    .io_en(rvclkhdr_237_io_en)
  );
  rvclkhdr rvclkhdr_238 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_238_io_clk),
    .io_en(rvclkhdr_238_io_en)
  );
  rvclkhdr rvclkhdr_239 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_239_io_clk),
    .io_en(rvclkhdr_239_io_en)
  );
  rvclkhdr rvclkhdr_240 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_240_io_clk),
    .io_en(rvclkhdr_240_io_en)
  );
  rvclkhdr rvclkhdr_241 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_241_io_clk),
    .io_en(rvclkhdr_241_io_en)
  );
  rvclkhdr rvclkhdr_242 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_242_io_clk),
    .io_en(rvclkhdr_242_io_en)
  );
  rvclkhdr rvclkhdr_243 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_243_io_clk),
    .io_en(rvclkhdr_243_io_en)
  );
  rvclkhdr rvclkhdr_244 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_244_io_clk),
    .io_en(rvclkhdr_244_io_en)
  );
  rvclkhdr rvclkhdr_245 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_245_io_clk),
    .io_en(rvclkhdr_245_io_en)
  );
  rvclkhdr rvclkhdr_246 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_246_io_clk),
    .io_en(rvclkhdr_246_io_en)
  );
  rvclkhdr rvclkhdr_247 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_247_io_clk),
    .io_en(rvclkhdr_247_io_en)
  );
  rvclkhdr rvclkhdr_248 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_248_io_clk),
    .io_en(rvclkhdr_248_io_en)
  );
  rvclkhdr rvclkhdr_249 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_249_io_clk),
    .io_en(rvclkhdr_249_io_en)
  );
  rvclkhdr rvclkhdr_250 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_250_io_clk),
    .io_en(rvclkhdr_250_io_en)
  );
  rvclkhdr rvclkhdr_251 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_251_io_clk),
    .io_en(rvclkhdr_251_io_en)
  );
  rvclkhdr rvclkhdr_252 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_252_io_clk),
    .io_en(rvclkhdr_252_io_en)
  );
  rvclkhdr rvclkhdr_253 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_253_io_clk),
    .io_en(rvclkhdr_253_io_en)
  );
  rvclkhdr rvclkhdr_254 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_254_io_clk),
    .io_en(rvclkhdr_254_io_en)
  );
  rvclkhdr rvclkhdr_255 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_255_io_clk),
    .io_en(rvclkhdr_255_io_en)
  );
  rvclkhdr rvclkhdr_256 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_256_io_clk),
    .io_en(rvclkhdr_256_io_en)
  );
  rvclkhdr rvclkhdr_257 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_257_io_clk),
    .io_en(rvclkhdr_257_io_en)
  );
  rvclkhdr rvclkhdr_258 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_258_io_clk),
    .io_en(rvclkhdr_258_io_en)
  );
  rvclkhdr rvclkhdr_259 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_259_io_clk),
    .io_en(rvclkhdr_259_io_en)
  );
  rvclkhdr rvclkhdr_260 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_260_io_clk),
    .io_en(rvclkhdr_260_io_en)
  );
  rvclkhdr rvclkhdr_261 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_261_io_clk),
    .io_en(rvclkhdr_261_io_en)
  );
  rvclkhdr rvclkhdr_262 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_262_io_clk),
    .io_en(rvclkhdr_262_io_en)
  );
  rvclkhdr rvclkhdr_263 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_263_io_clk),
    .io_en(rvclkhdr_263_io_en)
  );
  rvclkhdr rvclkhdr_264 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_264_io_clk),
    .io_en(rvclkhdr_264_io_en)
  );
  rvclkhdr rvclkhdr_265 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_265_io_clk),
    .io_en(rvclkhdr_265_io_en)
  );
  rvclkhdr rvclkhdr_266 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_266_io_clk),
    .io_en(rvclkhdr_266_io_en)
  );
  rvclkhdr rvclkhdr_267 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_267_io_clk),
    .io_en(rvclkhdr_267_io_en)
  );
  rvclkhdr rvclkhdr_268 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_268_io_clk),
    .io_en(rvclkhdr_268_io_en)
  );
  rvclkhdr rvclkhdr_269 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_269_io_clk),
    .io_en(rvclkhdr_269_io_en)
  );
  rvclkhdr rvclkhdr_270 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_270_io_clk),
    .io_en(rvclkhdr_270_io_en)
  );
  rvclkhdr rvclkhdr_271 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_271_io_clk),
    .io_en(rvclkhdr_271_io_en)
  );
  rvclkhdr rvclkhdr_272 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_272_io_clk),
    .io_en(rvclkhdr_272_io_en)
  );
  rvclkhdr rvclkhdr_273 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_273_io_clk),
    .io_en(rvclkhdr_273_io_en)
  );
  rvclkhdr rvclkhdr_274 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_274_io_clk),
    .io_en(rvclkhdr_274_io_en)
  );
  rvclkhdr rvclkhdr_275 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_275_io_clk),
    .io_en(rvclkhdr_275_io_en)
  );
  rvclkhdr rvclkhdr_276 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_276_io_clk),
    .io_en(rvclkhdr_276_io_en)
  );
  rvclkhdr rvclkhdr_277 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_277_io_clk),
    .io_en(rvclkhdr_277_io_en)
  );
  rvclkhdr rvclkhdr_278 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_278_io_clk),
    .io_en(rvclkhdr_278_io_en)
  );
  rvclkhdr rvclkhdr_279 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_279_io_clk),
    .io_en(rvclkhdr_279_io_en)
  );
  rvclkhdr rvclkhdr_280 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_280_io_clk),
    .io_en(rvclkhdr_280_io_en)
  );
  rvclkhdr rvclkhdr_281 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_281_io_clk),
    .io_en(rvclkhdr_281_io_en)
  );
  rvclkhdr rvclkhdr_282 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_282_io_clk),
    .io_en(rvclkhdr_282_io_en)
  );
  rvclkhdr rvclkhdr_283 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_283_io_clk),
    .io_en(rvclkhdr_283_io_en)
  );
  rvclkhdr rvclkhdr_284 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_284_io_clk),
    .io_en(rvclkhdr_284_io_en)
  );
  rvclkhdr rvclkhdr_285 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_285_io_clk),
    .io_en(rvclkhdr_285_io_en)
  );
  rvclkhdr rvclkhdr_286 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_286_io_clk),
    .io_en(rvclkhdr_286_io_en)
  );
  rvclkhdr rvclkhdr_287 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_287_io_clk),
    .io_en(rvclkhdr_287_io_en)
  );
  rvclkhdr rvclkhdr_288 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_288_io_clk),
    .io_en(rvclkhdr_288_io_en)
  );
  rvclkhdr rvclkhdr_289 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_289_io_clk),
    .io_en(rvclkhdr_289_io_en)
  );
  rvclkhdr rvclkhdr_290 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_290_io_clk),
    .io_en(rvclkhdr_290_io_en)
  );
  rvclkhdr rvclkhdr_291 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_291_io_clk),
    .io_en(rvclkhdr_291_io_en)
  );
  rvclkhdr rvclkhdr_292 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_292_io_clk),
    .io_en(rvclkhdr_292_io_en)
  );
  rvclkhdr rvclkhdr_293 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_293_io_clk),
    .io_en(rvclkhdr_293_io_en)
  );
  rvclkhdr rvclkhdr_294 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_294_io_clk),
    .io_en(rvclkhdr_294_io_en)
  );
  rvclkhdr rvclkhdr_295 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_295_io_clk),
    .io_en(rvclkhdr_295_io_en)
  );
  rvclkhdr rvclkhdr_296 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_296_io_clk),
    .io_en(rvclkhdr_296_io_en)
  );
  rvclkhdr rvclkhdr_297 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_297_io_clk),
    .io_en(rvclkhdr_297_io_en)
  );
  rvclkhdr rvclkhdr_298 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_298_io_clk),
    .io_en(rvclkhdr_298_io_en)
  );
  rvclkhdr rvclkhdr_299 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_299_io_clk),
    .io_en(rvclkhdr_299_io_en)
  );
  rvclkhdr rvclkhdr_300 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_300_io_clk),
    .io_en(rvclkhdr_300_io_en)
  );
  rvclkhdr rvclkhdr_301 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_301_io_clk),
    .io_en(rvclkhdr_301_io_en)
  );
  rvclkhdr rvclkhdr_302 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_302_io_clk),
    .io_en(rvclkhdr_302_io_en)
  );
  rvclkhdr rvclkhdr_303 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_303_io_clk),
    .io_en(rvclkhdr_303_io_en)
  );
  rvclkhdr rvclkhdr_304 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_304_io_clk),
    .io_en(rvclkhdr_304_io_en)
  );
  rvclkhdr rvclkhdr_305 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_305_io_clk),
    .io_en(rvclkhdr_305_io_en)
  );
  rvclkhdr rvclkhdr_306 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_306_io_clk),
    .io_en(rvclkhdr_306_io_en)
  );
  rvclkhdr rvclkhdr_307 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_307_io_clk),
    .io_en(rvclkhdr_307_io_en)
  );
  rvclkhdr rvclkhdr_308 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_308_io_clk),
    .io_en(rvclkhdr_308_io_en)
  );
  rvclkhdr rvclkhdr_309 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_309_io_clk),
    .io_en(rvclkhdr_309_io_en)
  );
  rvclkhdr rvclkhdr_310 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_310_io_clk),
    .io_en(rvclkhdr_310_io_en)
  );
  rvclkhdr rvclkhdr_311 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_311_io_clk),
    .io_en(rvclkhdr_311_io_en)
  );
  rvclkhdr rvclkhdr_312 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_312_io_clk),
    .io_en(rvclkhdr_312_io_en)
  );
  rvclkhdr rvclkhdr_313 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_313_io_clk),
    .io_en(rvclkhdr_313_io_en)
  );
  rvclkhdr rvclkhdr_314 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_314_io_clk),
    .io_en(rvclkhdr_314_io_en)
  );
  rvclkhdr rvclkhdr_315 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_315_io_clk),
    .io_en(rvclkhdr_315_io_en)
  );
  rvclkhdr rvclkhdr_316 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_316_io_clk),
    .io_en(rvclkhdr_316_io_en)
  );
  rvclkhdr rvclkhdr_317 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_317_io_clk),
    .io_en(rvclkhdr_317_io_en)
  );
  rvclkhdr rvclkhdr_318 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_318_io_clk),
    .io_en(rvclkhdr_318_io_en)
  );
  rvclkhdr rvclkhdr_319 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_319_io_clk),
    .io_en(rvclkhdr_319_io_en)
  );
  rvclkhdr rvclkhdr_320 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_320_io_clk),
    .io_en(rvclkhdr_320_io_en)
  );
  rvclkhdr rvclkhdr_321 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_321_io_clk),
    .io_en(rvclkhdr_321_io_en)
  );
  rvclkhdr rvclkhdr_322 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_322_io_clk),
    .io_en(rvclkhdr_322_io_en)
  );
  rvclkhdr rvclkhdr_323 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_323_io_clk),
    .io_en(rvclkhdr_323_io_en)
  );
  rvclkhdr rvclkhdr_324 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_324_io_clk),
    .io_en(rvclkhdr_324_io_en)
  );
  rvclkhdr rvclkhdr_325 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_325_io_clk),
    .io_en(rvclkhdr_325_io_en)
  );
  rvclkhdr rvclkhdr_326 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_326_io_clk),
    .io_en(rvclkhdr_326_io_en)
  );
  rvclkhdr rvclkhdr_327 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_327_io_clk),
    .io_en(rvclkhdr_327_io_en)
  );
  rvclkhdr rvclkhdr_328 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_328_io_clk),
    .io_en(rvclkhdr_328_io_en)
  );
  rvclkhdr rvclkhdr_329 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_329_io_clk),
    .io_en(rvclkhdr_329_io_en)
  );
  rvclkhdr rvclkhdr_330 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_330_io_clk),
    .io_en(rvclkhdr_330_io_en)
  );
  rvclkhdr rvclkhdr_331 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_331_io_clk),
    .io_en(rvclkhdr_331_io_en)
  );
  rvclkhdr rvclkhdr_332 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_332_io_clk),
    .io_en(rvclkhdr_332_io_en)
  );
  rvclkhdr rvclkhdr_333 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_333_io_clk),
    .io_en(rvclkhdr_333_io_en)
  );
  rvclkhdr rvclkhdr_334 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_334_io_clk),
    .io_en(rvclkhdr_334_io_en)
  );
  rvclkhdr rvclkhdr_335 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_335_io_clk),
    .io_en(rvclkhdr_335_io_en)
  );
  rvclkhdr rvclkhdr_336 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_336_io_clk),
    .io_en(rvclkhdr_336_io_en)
  );
  rvclkhdr rvclkhdr_337 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_337_io_clk),
    .io_en(rvclkhdr_337_io_en)
  );
  rvclkhdr rvclkhdr_338 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_338_io_clk),
    .io_en(rvclkhdr_338_io_en)
  );
  rvclkhdr rvclkhdr_339 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_339_io_clk),
    .io_en(rvclkhdr_339_io_en)
  );
  rvclkhdr rvclkhdr_340 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_340_io_clk),
    .io_en(rvclkhdr_340_io_en)
  );
  rvclkhdr rvclkhdr_341 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_341_io_clk),
    .io_en(rvclkhdr_341_io_en)
  );
  rvclkhdr rvclkhdr_342 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_342_io_clk),
    .io_en(rvclkhdr_342_io_en)
  );
  rvclkhdr rvclkhdr_343 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_343_io_clk),
    .io_en(rvclkhdr_343_io_en)
  );
  rvclkhdr rvclkhdr_344 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_344_io_clk),
    .io_en(rvclkhdr_344_io_en)
  );
  rvclkhdr rvclkhdr_345 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_345_io_clk),
    .io_en(rvclkhdr_345_io_en)
  );
  rvclkhdr rvclkhdr_346 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_346_io_clk),
    .io_en(rvclkhdr_346_io_en)
  );
  rvclkhdr rvclkhdr_347 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_347_io_clk),
    .io_en(rvclkhdr_347_io_en)
  );
  rvclkhdr rvclkhdr_348 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_348_io_clk),
    .io_en(rvclkhdr_348_io_en)
  );
  rvclkhdr rvclkhdr_349 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_349_io_clk),
    .io_en(rvclkhdr_349_io_en)
  );
  rvclkhdr rvclkhdr_350 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_350_io_clk),
    .io_en(rvclkhdr_350_io_en)
  );
  rvclkhdr rvclkhdr_351 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_351_io_clk),
    .io_en(rvclkhdr_351_io_en)
  );
  rvclkhdr rvclkhdr_352 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_352_io_clk),
    .io_en(rvclkhdr_352_io_en)
  );
  rvclkhdr rvclkhdr_353 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_353_io_clk),
    .io_en(rvclkhdr_353_io_en)
  );
  rvclkhdr rvclkhdr_354 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_354_io_clk),
    .io_en(rvclkhdr_354_io_en)
  );
  rvclkhdr rvclkhdr_355 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_355_io_clk),
    .io_en(rvclkhdr_355_io_en)
  );
  rvclkhdr rvclkhdr_356 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_356_io_clk),
    .io_en(rvclkhdr_356_io_en)
  );
  rvclkhdr rvclkhdr_357 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_357_io_clk),
    .io_en(rvclkhdr_357_io_en)
  );
  rvclkhdr rvclkhdr_358 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_358_io_clk),
    .io_en(rvclkhdr_358_io_en)
  );
  rvclkhdr rvclkhdr_359 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_359_io_clk),
    .io_en(rvclkhdr_359_io_en)
  );
  rvclkhdr rvclkhdr_360 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_360_io_clk),
    .io_en(rvclkhdr_360_io_en)
  );
  rvclkhdr rvclkhdr_361 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_361_io_clk),
    .io_en(rvclkhdr_361_io_en)
  );
  rvclkhdr rvclkhdr_362 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_362_io_clk),
    .io_en(rvclkhdr_362_io_en)
  );
  rvclkhdr rvclkhdr_363 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_363_io_clk),
    .io_en(rvclkhdr_363_io_en)
  );
  rvclkhdr rvclkhdr_364 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_364_io_clk),
    .io_en(rvclkhdr_364_io_en)
  );
  rvclkhdr rvclkhdr_365 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_365_io_clk),
    .io_en(rvclkhdr_365_io_en)
  );
  rvclkhdr rvclkhdr_366 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_366_io_clk),
    .io_en(rvclkhdr_366_io_en)
  );
  rvclkhdr rvclkhdr_367 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_367_io_clk),
    .io_en(rvclkhdr_367_io_en)
  );
  rvclkhdr rvclkhdr_368 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_368_io_clk),
    .io_en(rvclkhdr_368_io_en)
  );
  rvclkhdr rvclkhdr_369 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_369_io_clk),
    .io_en(rvclkhdr_369_io_en)
  );
  rvclkhdr rvclkhdr_370 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_370_io_clk),
    .io_en(rvclkhdr_370_io_en)
  );
  rvclkhdr rvclkhdr_371 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_371_io_clk),
    .io_en(rvclkhdr_371_io_en)
  );
  rvclkhdr rvclkhdr_372 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_372_io_clk),
    .io_en(rvclkhdr_372_io_en)
  );
  rvclkhdr rvclkhdr_373 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_373_io_clk),
    .io_en(rvclkhdr_373_io_en)
  );
  rvclkhdr rvclkhdr_374 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_374_io_clk),
    .io_en(rvclkhdr_374_io_en)
  );
  rvclkhdr rvclkhdr_375 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_375_io_clk),
    .io_en(rvclkhdr_375_io_en)
  );
  rvclkhdr rvclkhdr_376 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_376_io_clk),
    .io_en(rvclkhdr_376_io_en)
  );
  rvclkhdr rvclkhdr_377 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_377_io_clk),
    .io_en(rvclkhdr_377_io_en)
  );
  rvclkhdr rvclkhdr_378 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_378_io_clk),
    .io_en(rvclkhdr_378_io_en)
  );
  rvclkhdr rvclkhdr_379 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_379_io_clk),
    .io_en(rvclkhdr_379_io_en)
  );
  rvclkhdr rvclkhdr_380 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_380_io_clk),
    .io_en(rvclkhdr_380_io_en)
  );
  rvclkhdr rvclkhdr_381 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_381_io_clk),
    .io_en(rvclkhdr_381_io_en)
  );
  rvclkhdr rvclkhdr_382 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_382_io_clk),
    .io_en(rvclkhdr_382_io_en)
  );
  rvclkhdr rvclkhdr_383 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_383_io_clk),
    .io_en(rvclkhdr_383_io_en)
  );
  rvclkhdr rvclkhdr_384 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_384_io_clk),
    .io_en(rvclkhdr_384_io_en)
  );
  rvclkhdr rvclkhdr_385 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_385_io_clk),
    .io_en(rvclkhdr_385_io_en)
  );
  rvclkhdr rvclkhdr_386 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_386_io_clk),
    .io_en(rvclkhdr_386_io_en)
  );
  rvclkhdr rvclkhdr_387 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_387_io_clk),
    .io_en(rvclkhdr_387_io_en)
  );
  rvclkhdr rvclkhdr_388 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_388_io_clk),
    .io_en(rvclkhdr_388_io_en)
  );
  rvclkhdr rvclkhdr_389 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_389_io_clk),
    .io_en(rvclkhdr_389_io_en)
  );
  rvclkhdr rvclkhdr_390 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_390_io_clk),
    .io_en(rvclkhdr_390_io_en)
  );
  rvclkhdr rvclkhdr_391 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_391_io_clk),
    .io_en(rvclkhdr_391_io_en)
  );
  rvclkhdr rvclkhdr_392 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_392_io_clk),
    .io_en(rvclkhdr_392_io_en)
  );
  rvclkhdr rvclkhdr_393 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_393_io_clk),
    .io_en(rvclkhdr_393_io_en)
  );
  rvclkhdr rvclkhdr_394 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_394_io_clk),
    .io_en(rvclkhdr_394_io_en)
  );
  rvclkhdr rvclkhdr_395 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_395_io_clk),
    .io_en(rvclkhdr_395_io_en)
  );
  rvclkhdr rvclkhdr_396 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_396_io_clk),
    .io_en(rvclkhdr_396_io_en)
  );
  rvclkhdr rvclkhdr_397 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_397_io_clk),
    .io_en(rvclkhdr_397_io_en)
  );
  rvclkhdr rvclkhdr_398 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_398_io_clk),
    .io_en(rvclkhdr_398_io_en)
  );
  rvclkhdr rvclkhdr_399 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_399_io_clk),
    .io_en(rvclkhdr_399_io_en)
  );
  rvclkhdr rvclkhdr_400 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_400_io_clk),
    .io_en(rvclkhdr_400_io_en)
  );
  rvclkhdr rvclkhdr_401 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_401_io_clk),
    .io_en(rvclkhdr_401_io_en)
  );
  rvclkhdr rvclkhdr_402 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_402_io_clk),
    .io_en(rvclkhdr_402_io_en)
  );
  rvclkhdr rvclkhdr_403 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_403_io_clk),
    .io_en(rvclkhdr_403_io_en)
  );
  rvclkhdr rvclkhdr_404 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_404_io_clk),
    .io_en(rvclkhdr_404_io_en)
  );
  rvclkhdr rvclkhdr_405 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_405_io_clk),
    .io_en(rvclkhdr_405_io_en)
  );
  rvclkhdr rvclkhdr_406 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_406_io_clk),
    .io_en(rvclkhdr_406_io_en)
  );
  rvclkhdr rvclkhdr_407 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_407_io_clk),
    .io_en(rvclkhdr_407_io_en)
  );
  rvclkhdr rvclkhdr_408 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_408_io_clk),
    .io_en(rvclkhdr_408_io_en)
  );
  rvclkhdr rvclkhdr_409 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_409_io_clk),
    .io_en(rvclkhdr_409_io_en)
  );
  rvclkhdr rvclkhdr_410 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_410_io_clk),
    .io_en(rvclkhdr_410_io_en)
  );
  rvclkhdr rvclkhdr_411 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_411_io_clk),
    .io_en(rvclkhdr_411_io_en)
  );
  rvclkhdr rvclkhdr_412 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_412_io_clk),
    .io_en(rvclkhdr_412_io_en)
  );
  rvclkhdr rvclkhdr_413 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_413_io_clk),
    .io_en(rvclkhdr_413_io_en)
  );
  rvclkhdr rvclkhdr_414 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_414_io_clk),
    .io_en(rvclkhdr_414_io_en)
  );
  rvclkhdr rvclkhdr_415 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_415_io_clk),
    .io_en(rvclkhdr_415_io_en)
  );
  rvclkhdr rvclkhdr_416 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_416_io_clk),
    .io_en(rvclkhdr_416_io_en)
  );
  rvclkhdr rvclkhdr_417 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_417_io_clk),
    .io_en(rvclkhdr_417_io_en)
  );
  rvclkhdr rvclkhdr_418 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_418_io_clk),
    .io_en(rvclkhdr_418_io_en)
  );
  rvclkhdr rvclkhdr_419 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_419_io_clk),
    .io_en(rvclkhdr_419_io_en)
  );
  rvclkhdr rvclkhdr_420 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_420_io_clk),
    .io_en(rvclkhdr_420_io_en)
  );
  rvclkhdr rvclkhdr_421 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_421_io_clk),
    .io_en(rvclkhdr_421_io_en)
  );
  rvclkhdr rvclkhdr_422 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_422_io_clk),
    .io_en(rvclkhdr_422_io_en)
  );
  rvclkhdr rvclkhdr_423 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_423_io_clk),
    .io_en(rvclkhdr_423_io_en)
  );
  rvclkhdr rvclkhdr_424 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_424_io_clk),
    .io_en(rvclkhdr_424_io_en)
  );
  rvclkhdr rvclkhdr_425 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_425_io_clk),
    .io_en(rvclkhdr_425_io_en)
  );
  rvclkhdr rvclkhdr_426 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_426_io_clk),
    .io_en(rvclkhdr_426_io_en)
  );
  rvclkhdr rvclkhdr_427 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_427_io_clk),
    .io_en(rvclkhdr_427_io_en)
  );
  rvclkhdr rvclkhdr_428 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_428_io_clk),
    .io_en(rvclkhdr_428_io_en)
  );
  rvclkhdr rvclkhdr_429 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_429_io_clk),
    .io_en(rvclkhdr_429_io_en)
  );
  rvclkhdr rvclkhdr_430 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_430_io_clk),
    .io_en(rvclkhdr_430_io_en)
  );
  rvclkhdr rvclkhdr_431 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_431_io_clk),
    .io_en(rvclkhdr_431_io_en)
  );
  rvclkhdr rvclkhdr_432 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_432_io_clk),
    .io_en(rvclkhdr_432_io_en)
  );
  rvclkhdr rvclkhdr_433 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_433_io_clk),
    .io_en(rvclkhdr_433_io_en)
  );
  rvclkhdr rvclkhdr_434 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_434_io_clk),
    .io_en(rvclkhdr_434_io_en)
  );
  rvclkhdr rvclkhdr_435 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_435_io_clk),
    .io_en(rvclkhdr_435_io_en)
  );
  rvclkhdr rvclkhdr_436 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_436_io_clk),
    .io_en(rvclkhdr_436_io_en)
  );
  rvclkhdr rvclkhdr_437 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_437_io_clk),
    .io_en(rvclkhdr_437_io_en)
  );
  rvclkhdr rvclkhdr_438 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_438_io_clk),
    .io_en(rvclkhdr_438_io_en)
  );
  rvclkhdr rvclkhdr_439 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_439_io_clk),
    .io_en(rvclkhdr_439_io_en)
  );
  rvclkhdr rvclkhdr_440 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_440_io_clk),
    .io_en(rvclkhdr_440_io_en)
  );
  rvclkhdr rvclkhdr_441 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_441_io_clk),
    .io_en(rvclkhdr_441_io_en)
  );
  rvclkhdr rvclkhdr_442 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_442_io_clk),
    .io_en(rvclkhdr_442_io_en)
  );
  rvclkhdr rvclkhdr_443 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_443_io_clk),
    .io_en(rvclkhdr_443_io_en)
  );
  rvclkhdr rvclkhdr_444 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_444_io_clk),
    .io_en(rvclkhdr_444_io_en)
  );
  rvclkhdr rvclkhdr_445 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_445_io_clk),
    .io_en(rvclkhdr_445_io_en)
  );
  rvclkhdr rvclkhdr_446 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_446_io_clk),
    .io_en(rvclkhdr_446_io_en)
  );
  rvclkhdr rvclkhdr_447 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_447_io_clk),
    .io_en(rvclkhdr_447_io_en)
  );
  rvclkhdr rvclkhdr_448 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_448_io_clk),
    .io_en(rvclkhdr_448_io_en)
  );
  rvclkhdr rvclkhdr_449 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_449_io_clk),
    .io_en(rvclkhdr_449_io_en)
  );
  rvclkhdr rvclkhdr_450 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_450_io_clk),
    .io_en(rvclkhdr_450_io_en)
  );
  rvclkhdr rvclkhdr_451 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_451_io_clk),
    .io_en(rvclkhdr_451_io_en)
  );
  rvclkhdr rvclkhdr_452 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_452_io_clk),
    .io_en(rvclkhdr_452_io_en)
  );
  rvclkhdr rvclkhdr_453 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_453_io_clk),
    .io_en(rvclkhdr_453_io_en)
  );
  rvclkhdr rvclkhdr_454 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_454_io_clk),
    .io_en(rvclkhdr_454_io_en)
  );
  rvclkhdr rvclkhdr_455 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_455_io_clk),
    .io_en(rvclkhdr_455_io_en)
  );
  rvclkhdr rvclkhdr_456 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_456_io_clk),
    .io_en(rvclkhdr_456_io_en)
  );
  rvclkhdr rvclkhdr_457 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_457_io_clk),
    .io_en(rvclkhdr_457_io_en)
  );
  rvclkhdr rvclkhdr_458 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_458_io_clk),
    .io_en(rvclkhdr_458_io_en)
  );
  rvclkhdr rvclkhdr_459 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_459_io_clk),
    .io_en(rvclkhdr_459_io_en)
  );
  rvclkhdr rvclkhdr_460 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_460_io_clk),
    .io_en(rvclkhdr_460_io_en)
  );
  rvclkhdr rvclkhdr_461 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_461_io_clk),
    .io_en(rvclkhdr_461_io_en)
  );
  rvclkhdr rvclkhdr_462 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_462_io_clk),
    .io_en(rvclkhdr_462_io_en)
  );
  rvclkhdr rvclkhdr_463 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_463_io_clk),
    .io_en(rvclkhdr_463_io_en)
  );
  rvclkhdr rvclkhdr_464 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_464_io_clk),
    .io_en(rvclkhdr_464_io_en)
  );
  rvclkhdr rvclkhdr_465 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_465_io_clk),
    .io_en(rvclkhdr_465_io_en)
  );
  rvclkhdr rvclkhdr_466 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_466_io_clk),
    .io_en(rvclkhdr_466_io_en)
  );
  rvclkhdr rvclkhdr_467 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_467_io_clk),
    .io_en(rvclkhdr_467_io_en)
  );
  rvclkhdr rvclkhdr_468 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_468_io_clk),
    .io_en(rvclkhdr_468_io_en)
  );
  rvclkhdr rvclkhdr_469 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_469_io_clk),
    .io_en(rvclkhdr_469_io_en)
  );
  rvclkhdr rvclkhdr_470 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_470_io_clk),
    .io_en(rvclkhdr_470_io_en)
  );
  rvclkhdr rvclkhdr_471 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_471_io_clk),
    .io_en(rvclkhdr_471_io_en)
  );
  rvclkhdr rvclkhdr_472 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_472_io_clk),
    .io_en(rvclkhdr_472_io_en)
  );
  rvclkhdr rvclkhdr_473 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_473_io_clk),
    .io_en(rvclkhdr_473_io_en)
  );
  rvclkhdr rvclkhdr_474 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_474_io_clk),
    .io_en(rvclkhdr_474_io_en)
  );
  rvclkhdr rvclkhdr_475 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_475_io_clk),
    .io_en(rvclkhdr_475_io_en)
  );
  rvclkhdr rvclkhdr_476 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_476_io_clk),
    .io_en(rvclkhdr_476_io_en)
  );
  rvclkhdr rvclkhdr_477 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_477_io_clk),
    .io_en(rvclkhdr_477_io_en)
  );
  rvclkhdr rvclkhdr_478 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_478_io_clk),
    .io_en(rvclkhdr_478_io_en)
  );
  rvclkhdr rvclkhdr_479 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_479_io_clk),
    .io_en(rvclkhdr_479_io_en)
  );
  rvclkhdr rvclkhdr_480 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_480_io_clk),
    .io_en(rvclkhdr_480_io_en)
  );
  rvclkhdr rvclkhdr_481 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_481_io_clk),
    .io_en(rvclkhdr_481_io_en)
  );
  rvclkhdr rvclkhdr_482 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_482_io_clk),
    .io_en(rvclkhdr_482_io_en)
  );
  rvclkhdr rvclkhdr_483 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_483_io_clk),
    .io_en(rvclkhdr_483_io_en)
  );
  rvclkhdr rvclkhdr_484 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_484_io_clk),
    .io_en(rvclkhdr_484_io_en)
  );
  rvclkhdr rvclkhdr_485 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_485_io_clk),
    .io_en(rvclkhdr_485_io_en)
  );
  rvclkhdr rvclkhdr_486 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_486_io_clk),
    .io_en(rvclkhdr_486_io_en)
  );
  rvclkhdr rvclkhdr_487 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_487_io_clk),
    .io_en(rvclkhdr_487_io_en)
  );
  rvclkhdr rvclkhdr_488 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_488_io_clk),
    .io_en(rvclkhdr_488_io_en)
  );
  rvclkhdr rvclkhdr_489 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_489_io_clk),
    .io_en(rvclkhdr_489_io_en)
  );
  rvclkhdr rvclkhdr_490 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_490_io_clk),
    .io_en(rvclkhdr_490_io_en)
  );
  rvclkhdr rvclkhdr_491 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_491_io_clk),
    .io_en(rvclkhdr_491_io_en)
  );
  rvclkhdr rvclkhdr_492 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_492_io_clk),
    .io_en(rvclkhdr_492_io_en)
  );
  rvclkhdr rvclkhdr_493 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_493_io_clk),
    .io_en(rvclkhdr_493_io_en)
  );
  rvclkhdr rvclkhdr_494 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_494_io_clk),
    .io_en(rvclkhdr_494_io_en)
  );
  rvclkhdr rvclkhdr_495 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_495_io_clk),
    .io_en(rvclkhdr_495_io_en)
  );
  rvclkhdr rvclkhdr_496 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_496_io_clk),
    .io_en(rvclkhdr_496_io_en)
  );
  rvclkhdr rvclkhdr_497 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_497_io_clk),
    .io_en(rvclkhdr_497_io_en)
  );
  rvclkhdr rvclkhdr_498 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_498_io_clk),
    .io_en(rvclkhdr_498_io_en)
  );
  rvclkhdr rvclkhdr_499 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_499_io_clk),
    .io_en(rvclkhdr_499_io_en)
  );
  rvclkhdr rvclkhdr_500 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_500_io_clk),
    .io_en(rvclkhdr_500_io_en)
  );
  rvclkhdr rvclkhdr_501 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_501_io_clk),
    .io_en(rvclkhdr_501_io_en)
  );
  rvclkhdr rvclkhdr_502 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_502_io_clk),
    .io_en(rvclkhdr_502_io_en)
  );
  rvclkhdr rvclkhdr_503 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_503_io_clk),
    .io_en(rvclkhdr_503_io_en)
  );
  rvclkhdr rvclkhdr_504 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_504_io_clk),
    .io_en(rvclkhdr_504_io_en)
  );
  rvclkhdr rvclkhdr_505 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_505_io_clk),
    .io_en(rvclkhdr_505_io_en)
  );
  rvclkhdr rvclkhdr_506 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_506_io_clk),
    .io_en(rvclkhdr_506_io_en)
  );
  rvclkhdr rvclkhdr_507 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_507_io_clk),
    .io_en(rvclkhdr_507_io_en)
  );
  rvclkhdr rvclkhdr_508 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_508_io_clk),
    .io_en(rvclkhdr_508_io_en)
  );
  rvclkhdr rvclkhdr_509 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_509_io_clk),
    .io_en(rvclkhdr_509_io_en)
  );
  rvclkhdr rvclkhdr_510 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_510_io_clk),
    .io_en(rvclkhdr_510_io_en)
  );
  rvclkhdr rvclkhdr_511 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_511_io_clk),
    .io_en(rvclkhdr_511_io_en)
  );
  rvclkhdr rvclkhdr_512 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_512_io_clk),
    .io_en(rvclkhdr_512_io_en)
  );
  rvclkhdr rvclkhdr_513 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_513_io_clk),
    .io_en(rvclkhdr_513_io_en)
  );
  rvclkhdr rvclkhdr_514 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_514_io_clk),
    .io_en(rvclkhdr_514_io_en)
  );
  rvclkhdr rvclkhdr_515 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_515_io_clk),
    .io_en(rvclkhdr_515_io_en)
  );
  rvclkhdr rvclkhdr_516 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_516_io_clk),
    .io_en(rvclkhdr_516_io_en)
  );
  rvclkhdr rvclkhdr_517 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_517_io_clk),
    .io_en(rvclkhdr_517_io_en)
  );
  rvclkhdr rvclkhdr_518 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_518_io_clk),
    .io_en(rvclkhdr_518_io_en)
  );
  rvclkhdr rvclkhdr_519 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_519_io_clk),
    .io_en(rvclkhdr_519_io_en)
  );
  rvclkhdr rvclkhdr_520 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_520_io_clk),
    .io_en(rvclkhdr_520_io_en)
  );
  rvclkhdr rvclkhdr_521 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_521_io_clk),
    .io_en(rvclkhdr_521_io_en)
  );
  rvclkhdr rvclkhdr_522 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_522_io_clk),
    .io_en(rvclkhdr_522_io_en)
  );
  rvclkhdr rvclkhdr_523 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_523_io_clk),
    .io_en(rvclkhdr_523_io_en)
  );
  rvclkhdr rvclkhdr_524 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_524_io_clk),
    .io_en(rvclkhdr_524_io_en)
  );
  rvclkhdr rvclkhdr_525 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_525_io_clk),
    .io_en(rvclkhdr_525_io_en)
  );
  rvclkhdr rvclkhdr_526 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_526_io_clk),
    .io_en(rvclkhdr_526_io_en)
  );
  rvclkhdr rvclkhdr_527 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_527_io_clk),
    .io_en(rvclkhdr_527_io_en)
  );
  rvclkhdr rvclkhdr_528 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_528_io_clk),
    .io_en(rvclkhdr_528_io_en)
  );
  rvclkhdr rvclkhdr_529 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_529_io_clk),
    .io_en(rvclkhdr_529_io_en)
  );
  rvclkhdr rvclkhdr_530 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_530_io_clk),
    .io_en(rvclkhdr_530_io_en)
  );
  rvclkhdr rvclkhdr_531 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_531_io_clk),
    .io_en(rvclkhdr_531_io_en)
  );
  rvclkhdr rvclkhdr_532 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_532_io_clk),
    .io_en(rvclkhdr_532_io_en)
  );
  rvclkhdr rvclkhdr_533 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_533_io_clk),
    .io_en(rvclkhdr_533_io_en)
  );
  rvclkhdr rvclkhdr_534 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_534_io_clk),
    .io_en(rvclkhdr_534_io_en)
  );
  rvclkhdr rvclkhdr_535 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_535_io_clk),
    .io_en(rvclkhdr_535_io_en)
  );
  rvclkhdr rvclkhdr_536 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_536_io_clk),
    .io_en(rvclkhdr_536_io_en)
  );
  rvclkhdr rvclkhdr_537 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_537_io_clk),
    .io_en(rvclkhdr_537_io_en)
  );
  rvclkhdr rvclkhdr_538 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_538_io_clk),
    .io_en(rvclkhdr_538_io_en)
  );
  rvclkhdr rvclkhdr_539 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_539_io_clk),
    .io_en(rvclkhdr_539_io_en)
  );
  rvclkhdr rvclkhdr_540 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_540_io_clk),
    .io_en(rvclkhdr_540_io_en)
  );
  rvclkhdr rvclkhdr_541 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_541_io_clk),
    .io_en(rvclkhdr_541_io_en)
  );
  rvclkhdr rvclkhdr_542 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_542_io_clk),
    .io_en(rvclkhdr_542_io_en)
  );
  rvclkhdr rvclkhdr_543 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_543_io_clk),
    .io_en(rvclkhdr_543_io_en)
  );
  rvclkhdr rvclkhdr_544 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_544_io_clk),
    .io_en(rvclkhdr_544_io_en)
  );
  rvclkhdr rvclkhdr_545 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_545_io_clk),
    .io_en(rvclkhdr_545_io_en)
  );
  rvclkhdr rvclkhdr_546 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_546_io_clk),
    .io_en(rvclkhdr_546_io_en)
  );
  rvclkhdr rvclkhdr_547 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_547_io_clk),
    .io_en(rvclkhdr_547_io_en)
  );
  rvclkhdr rvclkhdr_548 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_548_io_clk),
    .io_en(rvclkhdr_548_io_en)
  );
  rvclkhdr rvclkhdr_549 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_549_io_clk),
    .io_en(rvclkhdr_549_io_en)
  );
  rvclkhdr rvclkhdr_550 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_550_io_clk),
    .io_en(rvclkhdr_550_io_en)
  );
  rvclkhdr rvclkhdr_551 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_551_io_clk),
    .io_en(rvclkhdr_551_io_en)
  );
  rvclkhdr rvclkhdr_552 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_552_io_clk),
    .io_en(rvclkhdr_552_io_en)
  );
  assign io_ifu_bp_hit_taken_f = _T_231 & _T_232; // @[ifu_bp_ctl.scala 277:25]
  assign io_ifu_bp_btb_target_f = _T_443 | _T_453; // @[ifu_bp_ctl.scala 374:26]
  assign io_ifu_bp_inst_mask_f = _T_268 | _T_269; // @[ifu_bp_ctl.scala 302:25]
  assign io_ifu_bp_fghr_f = fghr; // @[ifu_bp_ctl.scala 345:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_154; // @[ifu_bp_ctl.scala 254:19]
  assign io_ifu_bp_ret_f = {_T_288,_T_294}; // @[ifu_bp_ctl.scala 351:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_273; // @[ifu_bp_ctl.scala 346:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[ifu_bp_ctl.scala 347:21]
  assign io_ifu_bp_pc4_f = {_T_279,_T_282}; // @[ifu_bp_ctl.scala 348:19]
  assign io_ifu_bp_valid_f = vwayhit_f & _T_353; // @[ifu_bp_ctl.scala 350:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 362:23]
  assign io_ifu_bp_fa_index_f_0 = 9'h0; // @[ifu_bp_ctl.scala 35:24]
  assign io_ifu_bp_fa_index_f_1 = 9'h0; // @[ifu_bp_ctl.scala 35:24]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_io_en = io_ifc_fetch_req_f | exu_mp_valid; // @[lib.scala 412:17]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_1_io_en = ~rs_hold; // @[lib.scala 412:17]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_2_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_3_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_4_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_5_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_6_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_7_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_8_io_en = _T_494 & io_ifu_bp_hit_taken_f; // @[lib.scala 412:17]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_9_io_en = _T_613 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_10_io_en = _T_616 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_11_io_en = _T_619 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_12_io_en = _T_622 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_13_io_en = _T_625 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_14_io_en = _T_628 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_15_io_en = _T_631 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_16_io_en = _T_634 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_17_io_en = _T_637 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_18_io_en = _T_640 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_19_io_en = _T_643 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_20_io_en = _T_646 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_21_io_en = _T_649 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_22_io_en = _T_652 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_23_io_en = _T_655 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_24_io_en = _T_658 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_25_io_en = _T_661 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_26_io_en = _T_664 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_27_io_en = _T_667 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_28_io_en = _T_670 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_29_io_en = _T_673 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_30_io_en = _T_676 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_31_io_en = _T_679 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_32_io_en = _T_682 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_33_io_en = _T_685 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_34_io_en = _T_688 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_35_io_en = _T_691 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_36_io_en = _T_694 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_37_io_en = _T_697 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_38_io_en = _T_700 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_39_io_en = _T_703 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_40_io_en = _T_706 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_41_io_en = _T_709 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_42_io_en = _T_712 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_43_io_en = _T_715 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_44_io_en = _T_718 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_45_io_en = _T_721 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_46_io_en = _T_724 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_47_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_47_io_en = _T_727 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_48_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_48_io_en = _T_730 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_49_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_49_io_en = _T_733 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_50_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_50_io_en = _T_736 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_51_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_51_io_en = _T_739 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_52_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_52_io_en = _T_742 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_53_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_53_io_en = _T_745 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_54_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_54_io_en = _T_748 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_55_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_55_io_en = _T_751 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_56_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_56_io_en = _T_754 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_57_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_57_io_en = _T_757 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_58_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_58_io_en = _T_760 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_59_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_59_io_en = _T_763 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_60_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_60_io_en = _T_766 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_61_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_61_io_en = _T_769 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_62_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_62_io_en = _T_772 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_63_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_63_io_en = _T_775 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_64_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_64_io_en = _T_778 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_65_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_65_io_en = _T_781 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_66_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_66_io_en = _T_784 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_67_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_67_io_en = _T_787 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_68_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_68_io_en = _T_790 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_69_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_69_io_en = _T_793 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_70_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_70_io_en = _T_796 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_71_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_71_io_en = _T_799 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_72_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_72_io_en = _T_802 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_73_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_73_io_en = _T_805 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_74_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_74_io_en = _T_808 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_75_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_75_io_en = _T_811 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_76_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_76_io_en = _T_814 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_77_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_77_io_en = _T_817 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_78_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_78_io_en = _T_820 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_79_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_79_io_en = _T_823 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_80_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_80_io_en = _T_826 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_81_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_81_io_en = _T_829 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_82_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_82_io_en = _T_832 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_83_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_83_io_en = _T_835 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_84_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_84_io_en = _T_838 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_85_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_85_io_en = _T_841 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_86_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_86_io_en = _T_844 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_87_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_87_io_en = _T_847 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_88_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_88_io_en = _T_850 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_89_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_89_io_en = _T_853 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_90_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_90_io_en = _T_856 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_91_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_91_io_en = _T_859 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_92_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_92_io_en = _T_862 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_93_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_93_io_en = _T_865 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_94_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_94_io_en = _T_868 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_95_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_95_io_en = _T_871 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_96_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_96_io_en = _T_874 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_97_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_97_io_en = _T_877 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_98_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_98_io_en = _T_880 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_99_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_99_io_en = _T_883 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_100_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_100_io_en = _T_886 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_101_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_101_io_en = _T_889 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_102_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_102_io_en = _T_892 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_103_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_103_io_en = _T_895 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_104_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_104_io_en = _T_898 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_105_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_105_io_en = _T_901 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_106_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_106_io_en = _T_904 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_107_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_107_io_en = _T_907 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_108_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_108_io_en = _T_910 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_109_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_109_io_en = _T_913 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_110_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_110_io_en = _T_916 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_111_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_111_io_en = _T_919 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_112_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_112_io_en = _T_922 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_113_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_113_io_en = _T_925 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_114_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_114_io_en = _T_928 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_115_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_115_io_en = _T_931 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_116_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_116_io_en = _T_934 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_117_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_117_io_en = _T_937 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_118_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_118_io_en = _T_940 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_119_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_119_io_en = _T_943 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_120_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_120_io_en = _T_946 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_121_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_121_io_en = _T_949 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_122_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_122_io_en = _T_952 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_123_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_123_io_en = _T_955 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_124_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_124_io_en = _T_958 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_125_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_125_io_en = _T_961 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_126_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_126_io_en = _T_964 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_127_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_127_io_en = _T_967 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_128_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_128_io_en = _T_970 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_129_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_129_io_en = _T_973 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_130_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_130_io_en = _T_976 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_131_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_131_io_en = _T_979 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_132_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_132_io_en = _T_982 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_133_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_133_io_en = _T_985 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_134_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_134_io_en = _T_988 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_135_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_135_io_en = _T_991 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_136_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_136_io_en = _T_994 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_137_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_137_io_en = _T_997 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_138_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_138_io_en = _T_1000 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_139_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_139_io_en = _T_1003 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_140_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_140_io_en = _T_1006 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_141_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_141_io_en = _T_1009 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_142_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_142_io_en = _T_1012 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_143_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_143_io_en = _T_1015 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_144_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_144_io_en = _T_1018 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_145_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_145_io_en = _T_1021 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_146_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_146_io_en = _T_1024 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_147_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_147_io_en = _T_1027 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_148_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_148_io_en = _T_1030 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_149_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_149_io_en = _T_1033 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_150_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_150_io_en = _T_1036 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_151_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_151_io_en = _T_1039 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_152_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_152_io_en = _T_1042 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_153_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_153_io_en = _T_1045 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_154_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_154_io_en = _T_1048 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_155_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_155_io_en = _T_1051 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_156_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_156_io_en = _T_1054 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_157_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_157_io_en = _T_1057 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_158_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_158_io_en = _T_1060 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_159_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_159_io_en = _T_1063 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_160_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_160_io_en = _T_1066 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_161_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_161_io_en = _T_1069 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_162_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_162_io_en = _T_1072 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_163_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_163_io_en = _T_1075 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_164_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_164_io_en = _T_1078 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_165_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_165_io_en = _T_1081 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_166_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_166_io_en = _T_1084 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_167_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_167_io_en = _T_1087 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_168_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_168_io_en = _T_1090 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_169_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_169_io_en = _T_1093 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_170_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_170_io_en = _T_1096 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_171_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_171_io_en = _T_1099 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_172_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_172_io_en = _T_1102 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_173_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_173_io_en = _T_1105 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_174_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_174_io_en = _T_1108 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_175_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_175_io_en = _T_1111 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_176_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_176_io_en = _T_1114 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_177_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_177_io_en = _T_1117 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_178_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_178_io_en = _T_1120 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_179_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_179_io_en = _T_1123 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_180_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_180_io_en = _T_1126 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_181_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_181_io_en = _T_1129 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_182_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_182_io_en = _T_1132 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_183_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_183_io_en = _T_1135 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_184_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_184_io_en = _T_1138 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_185_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_185_io_en = _T_1141 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_186_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_186_io_en = _T_1144 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_187_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_187_io_en = _T_1147 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_188_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_188_io_en = _T_1150 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_189_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_189_io_en = _T_1153 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_190_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_190_io_en = _T_1156 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_191_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_191_io_en = _T_1159 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_192_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_192_io_en = _T_1162 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_193_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_193_io_en = _T_1165 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_194_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_194_io_en = _T_1168 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_195_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_195_io_en = _T_1171 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_196_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_196_io_en = _T_1174 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_197_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_197_io_en = _T_1177 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_198_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_198_io_en = _T_1180 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_199_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_199_io_en = _T_1183 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_200_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_200_io_en = _T_1186 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_201_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_201_io_en = _T_1189 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_202_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_202_io_en = _T_1192 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_203_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_203_io_en = _T_1195 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_204_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_204_io_en = _T_1198 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_205_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_205_io_en = _T_1201 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_206_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_206_io_en = _T_1204 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_207_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_207_io_en = _T_1207 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_208_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_208_io_en = _T_1210 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_209_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_209_io_en = _T_1213 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_210_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_210_io_en = _T_1216 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_211_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_211_io_en = _T_1219 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_212_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_212_io_en = _T_1222 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_213_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_213_io_en = _T_1225 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_214_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_214_io_en = _T_1228 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_215_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_215_io_en = _T_1231 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_216_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_216_io_en = _T_1234 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_217_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_217_io_en = _T_1237 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_218_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_218_io_en = _T_1240 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_219_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_219_io_en = _T_1243 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_220_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_220_io_en = _T_1246 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_221_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_221_io_en = _T_1249 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_222_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_222_io_en = _T_1252 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_223_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_223_io_en = _T_1255 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_224_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_224_io_en = _T_1258 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_225_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_225_io_en = _T_1261 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_226_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_226_io_en = _T_1264 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_227_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_227_io_en = _T_1267 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_228_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_228_io_en = _T_1270 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_229_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_229_io_en = _T_1273 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_230_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_230_io_en = _T_1276 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_231_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_231_io_en = _T_1279 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_232_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_232_io_en = _T_1282 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_233_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_233_io_en = _T_1285 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_234_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_234_io_en = _T_1288 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_235_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_235_io_en = _T_1291 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_236_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_236_io_en = _T_1294 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_237_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_237_io_en = _T_1297 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_238_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_238_io_en = _T_1300 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_239_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_239_io_en = _T_1303 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_240_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_240_io_en = _T_1306 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_241_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_241_io_en = _T_1309 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_242_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_242_io_en = _T_1312 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_243_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_243_io_en = _T_1315 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_244_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_244_io_en = _T_1318 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_245_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_245_io_en = _T_1321 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_246_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_246_io_en = _T_1324 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_247_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_247_io_en = _T_1327 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_248_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_248_io_en = _T_1330 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_249_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_249_io_en = _T_1333 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_250_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_250_io_en = _T_1336 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_251_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_251_io_en = _T_1339 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_252_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_252_io_en = _T_1342 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_253_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_253_io_en = _T_1345 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_254_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_254_io_en = _T_1348 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_255_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_255_io_en = _T_1351 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_256_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_256_io_en = _T_1354 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_257_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_257_io_en = _T_1357 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_258_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_258_io_en = _T_1360 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_259_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_259_io_en = _T_1363 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_260_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_260_io_en = _T_1366 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_261_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_261_io_en = _T_1369 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_262_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_262_io_en = _T_1372 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_263_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_263_io_en = _T_1375 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_264_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_264_io_en = _T_1378 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_265_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_265_io_en = _T_613 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_266_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_266_io_en = _T_616 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_267_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_267_io_en = _T_619 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_268_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_268_io_en = _T_622 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_269_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_269_io_en = _T_625 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_270_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_270_io_en = _T_628 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_271_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_271_io_en = _T_631 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_272_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_272_io_en = _T_634 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_273_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_273_io_en = _T_637 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_274_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_274_io_en = _T_640 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_275_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_275_io_en = _T_643 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_276_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_276_io_en = _T_646 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_277_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_277_io_en = _T_649 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_278_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_278_io_en = _T_652 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_279_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_279_io_en = _T_655 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_280_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_280_io_en = _T_658 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_281_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_281_io_en = _T_661 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_282_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_282_io_en = _T_664 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_283_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_283_io_en = _T_667 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_284_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_284_io_en = _T_670 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_285_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_285_io_en = _T_673 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_286_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_286_io_en = _T_676 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_287_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_287_io_en = _T_679 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_288_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_288_io_en = _T_682 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_289_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_289_io_en = _T_685 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_290_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_290_io_en = _T_688 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_291_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_291_io_en = _T_691 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_292_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_292_io_en = _T_694 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_293_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_293_io_en = _T_697 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_294_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_294_io_en = _T_700 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_295_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_295_io_en = _T_703 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_296_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_296_io_en = _T_706 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_297_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_297_io_en = _T_709 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_298_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_298_io_en = _T_712 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_299_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_299_io_en = _T_715 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_300_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_300_io_en = _T_718 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_301_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_301_io_en = _T_721 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_302_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_302_io_en = _T_724 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_303_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_303_io_en = _T_727 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_304_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_304_io_en = _T_730 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_305_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_305_io_en = _T_733 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_306_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_306_io_en = _T_736 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_307_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_307_io_en = _T_739 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_308_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_308_io_en = _T_742 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_309_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_309_io_en = _T_745 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_310_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_310_io_en = _T_748 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_311_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_311_io_en = _T_751 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_312_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_312_io_en = _T_754 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_313_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_313_io_en = _T_757 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_314_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_314_io_en = _T_760 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_315_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_315_io_en = _T_763 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_316_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_316_io_en = _T_766 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_317_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_317_io_en = _T_769 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_318_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_318_io_en = _T_772 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_319_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_319_io_en = _T_775 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_320_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_320_io_en = _T_778 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_321_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_321_io_en = _T_781 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_322_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_322_io_en = _T_784 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_323_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_323_io_en = _T_787 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_324_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_324_io_en = _T_790 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_325_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_325_io_en = _T_793 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_326_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_326_io_en = _T_796 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_327_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_327_io_en = _T_799 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_328_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_328_io_en = _T_802 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_329_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_329_io_en = _T_805 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_330_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_330_io_en = _T_808 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_331_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_331_io_en = _T_811 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_332_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_332_io_en = _T_814 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_333_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_333_io_en = _T_817 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_334_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_334_io_en = _T_820 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_335_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_335_io_en = _T_823 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_336_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_336_io_en = _T_826 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_337_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_337_io_en = _T_829 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_338_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_338_io_en = _T_832 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_339_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_339_io_en = _T_835 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_340_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_340_io_en = _T_838 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_341_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_341_io_en = _T_841 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_342_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_342_io_en = _T_844 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_343_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_343_io_en = _T_847 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_344_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_344_io_en = _T_850 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_345_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_345_io_en = _T_853 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_346_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_346_io_en = _T_856 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_347_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_347_io_en = _T_859 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_348_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_348_io_en = _T_862 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_349_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_349_io_en = _T_865 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_350_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_350_io_en = _T_868 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_351_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_351_io_en = _T_871 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_352_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_352_io_en = _T_874 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_353_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_353_io_en = _T_877 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_354_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_354_io_en = _T_880 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_355_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_355_io_en = _T_883 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_356_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_356_io_en = _T_886 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_357_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_357_io_en = _T_889 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_358_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_358_io_en = _T_892 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_359_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_359_io_en = _T_895 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_360_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_360_io_en = _T_898 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_361_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_361_io_en = _T_901 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_362_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_362_io_en = _T_904 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_363_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_363_io_en = _T_907 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_364_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_364_io_en = _T_910 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_365_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_365_io_en = _T_913 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_366_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_366_io_en = _T_916 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_367_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_367_io_en = _T_919 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_368_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_368_io_en = _T_922 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_369_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_369_io_en = _T_925 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_370_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_370_io_en = _T_928 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_371_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_371_io_en = _T_931 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_372_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_372_io_en = _T_934 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_373_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_373_io_en = _T_937 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_374_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_374_io_en = _T_940 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_375_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_375_io_en = _T_943 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_376_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_376_io_en = _T_946 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_377_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_377_io_en = _T_949 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_378_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_378_io_en = _T_952 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_379_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_379_io_en = _T_955 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_380_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_380_io_en = _T_958 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_381_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_381_io_en = _T_961 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_382_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_382_io_en = _T_964 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_383_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_383_io_en = _T_967 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_384_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_384_io_en = _T_970 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_385_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_385_io_en = _T_973 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_386_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_386_io_en = _T_976 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_387_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_387_io_en = _T_979 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_388_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_388_io_en = _T_982 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_389_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_389_io_en = _T_985 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_390_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_390_io_en = _T_988 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_391_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_391_io_en = _T_991 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_392_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_392_io_en = _T_994 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_393_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_393_io_en = _T_997 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_394_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_394_io_en = _T_1000 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_395_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_395_io_en = _T_1003 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_396_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_396_io_en = _T_1006 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_397_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_397_io_en = _T_1009 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_398_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_398_io_en = _T_1012 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_399_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_399_io_en = _T_1015 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_400_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_400_io_en = _T_1018 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_401_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_401_io_en = _T_1021 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_402_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_402_io_en = _T_1024 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_403_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_403_io_en = _T_1027 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_404_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_404_io_en = _T_1030 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_405_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_405_io_en = _T_1033 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_406_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_406_io_en = _T_1036 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_407_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_407_io_en = _T_1039 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_408_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_408_io_en = _T_1042 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_409_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_409_io_en = _T_1045 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_410_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_410_io_en = _T_1048 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_411_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_411_io_en = _T_1051 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_412_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_412_io_en = _T_1054 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_413_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_413_io_en = _T_1057 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_414_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_414_io_en = _T_1060 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_415_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_415_io_en = _T_1063 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_416_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_416_io_en = _T_1066 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_417_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_417_io_en = _T_1069 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_418_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_418_io_en = _T_1072 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_419_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_419_io_en = _T_1075 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_420_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_420_io_en = _T_1078 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_421_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_421_io_en = _T_1081 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_422_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_422_io_en = _T_1084 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_423_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_423_io_en = _T_1087 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_424_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_424_io_en = _T_1090 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_425_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_425_io_en = _T_1093 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_426_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_426_io_en = _T_1096 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_427_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_427_io_en = _T_1099 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_428_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_428_io_en = _T_1102 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_429_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_429_io_en = _T_1105 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_430_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_430_io_en = _T_1108 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_431_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_431_io_en = _T_1111 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_432_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_432_io_en = _T_1114 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_433_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_433_io_en = _T_1117 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_434_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_434_io_en = _T_1120 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_435_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_435_io_en = _T_1123 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_436_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_436_io_en = _T_1126 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_437_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_437_io_en = _T_1129 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_438_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_438_io_en = _T_1132 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_439_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_439_io_en = _T_1135 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_440_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_440_io_en = _T_1138 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_441_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_441_io_en = _T_1141 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_442_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_442_io_en = _T_1144 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_443_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_443_io_en = _T_1147 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_444_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_444_io_en = _T_1150 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_445_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_445_io_en = _T_1153 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_446_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_446_io_en = _T_1156 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_447_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_447_io_en = _T_1159 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_448_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_448_io_en = _T_1162 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_449_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_449_io_en = _T_1165 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_450_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_450_io_en = _T_1168 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_451_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_451_io_en = _T_1171 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_452_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_452_io_en = _T_1174 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_453_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_453_io_en = _T_1177 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_454_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_454_io_en = _T_1180 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_455_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_455_io_en = _T_1183 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_456_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_456_io_en = _T_1186 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_457_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_457_io_en = _T_1189 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_458_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_458_io_en = _T_1192 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_459_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_459_io_en = _T_1195 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_460_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_460_io_en = _T_1198 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_461_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_461_io_en = _T_1201 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_462_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_462_io_en = _T_1204 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_463_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_463_io_en = _T_1207 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_464_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_464_io_en = _T_1210 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_465_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_465_io_en = _T_1213 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_466_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_466_io_en = _T_1216 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_467_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_467_io_en = _T_1219 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_468_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_468_io_en = _T_1222 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_469_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_469_io_en = _T_1225 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_470_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_470_io_en = _T_1228 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_471_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_471_io_en = _T_1231 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_472_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_472_io_en = _T_1234 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_473_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_473_io_en = _T_1237 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_474_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_474_io_en = _T_1240 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_475_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_475_io_en = _T_1243 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_476_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_476_io_en = _T_1246 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_477_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_477_io_en = _T_1249 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_478_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_478_io_en = _T_1252 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_479_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_479_io_en = _T_1255 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_480_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_480_io_en = _T_1258 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_481_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_481_io_en = _T_1261 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_482_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_482_io_en = _T_1264 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_483_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_483_io_en = _T_1267 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_484_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_484_io_en = _T_1270 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_485_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_485_io_en = _T_1273 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_486_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_486_io_en = _T_1276 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_487_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_487_io_en = _T_1279 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_488_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_488_io_en = _T_1282 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_489_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_489_io_en = _T_1285 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_490_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_490_io_en = _T_1288 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_491_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_491_io_en = _T_1291 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_492_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_492_io_en = _T_1294 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_493_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_493_io_en = _T_1297 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_494_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_494_io_en = _T_1300 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_495_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_495_io_en = _T_1303 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_496_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_496_io_en = _T_1306 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_497_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_497_io_en = _T_1309 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_498_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_498_io_en = _T_1312 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_499_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_499_io_en = _T_1315 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_500_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_500_io_en = _T_1318 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_501_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_501_io_en = _T_1321 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_502_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_502_io_en = _T_1324 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_503_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_503_io_en = _T_1327 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_504_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_504_io_en = _T_1330 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_505_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_505_io_en = _T_1333 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_506_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_506_io_en = _T_1336 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_507_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_507_io_en = _T_1339 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_508_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_508_io_en = _T_1342 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_509_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_509_io_en = _T_1345 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_510_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_510_io_en = _T_1348 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_511_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_511_io_en = _T_1351 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_512_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_512_io_en = _T_1354 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_513_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_513_io_en = _T_1357 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_514_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_514_io_en = _T_1360 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_515_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_515_io_en = _T_1363 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_516_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_516_io_en = _T_1366 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_517_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_517_io_en = _T_1369 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_518_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_518_io_en = _T_1372 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_519_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_519_io_en = _T_1375 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_520_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_520_io_en = _T_1378 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_521_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_521_io_en = _T_6249 | _T_6254; // @[lib.scala 345:16]
  assign rvclkhdr_522_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_522_io_en = _T_6260 | _T_6265; // @[lib.scala 345:16]
  assign rvclkhdr_523_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_523_io_en = _T_6271 | _T_6276; // @[lib.scala 345:16]
  assign rvclkhdr_524_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_524_io_en = _T_6282 | _T_6287; // @[lib.scala 345:16]
  assign rvclkhdr_525_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_525_io_en = _T_6293 | _T_6298; // @[lib.scala 345:16]
  assign rvclkhdr_526_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_526_io_en = _T_6304 | _T_6309; // @[lib.scala 345:16]
  assign rvclkhdr_527_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_527_io_en = _T_6315 | _T_6320; // @[lib.scala 345:16]
  assign rvclkhdr_528_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_528_io_en = _T_6326 | _T_6331; // @[lib.scala 345:16]
  assign rvclkhdr_529_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_529_io_en = _T_6337 | _T_6342; // @[lib.scala 345:16]
  assign rvclkhdr_530_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_530_io_en = _T_6348 | _T_6353; // @[lib.scala 345:16]
  assign rvclkhdr_531_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_531_io_en = _T_6359 | _T_6364; // @[lib.scala 345:16]
  assign rvclkhdr_532_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_532_io_en = _T_6370 | _T_6375; // @[lib.scala 345:16]
  assign rvclkhdr_533_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_533_io_en = _T_6381 | _T_6386; // @[lib.scala 345:16]
  assign rvclkhdr_534_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_534_io_en = _T_6392 | _T_6397; // @[lib.scala 345:16]
  assign rvclkhdr_535_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_535_io_en = _T_6403 | _T_6408; // @[lib.scala 345:16]
  assign rvclkhdr_536_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_536_io_en = _T_6414 | _T_6419; // @[lib.scala 345:16]
  assign rvclkhdr_537_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_537_io_en = _T_6425 | _T_6430; // @[lib.scala 345:16]
  assign rvclkhdr_538_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_538_io_en = _T_6436 | _T_6441; // @[lib.scala 345:16]
  assign rvclkhdr_539_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_539_io_en = _T_6447 | _T_6452; // @[lib.scala 345:16]
  assign rvclkhdr_540_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_540_io_en = _T_6458 | _T_6463; // @[lib.scala 345:16]
  assign rvclkhdr_541_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_541_io_en = _T_6469 | _T_6474; // @[lib.scala 345:16]
  assign rvclkhdr_542_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_542_io_en = _T_6480 | _T_6485; // @[lib.scala 345:16]
  assign rvclkhdr_543_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_543_io_en = _T_6491 | _T_6496; // @[lib.scala 345:16]
  assign rvclkhdr_544_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_544_io_en = _T_6502 | _T_6507; // @[lib.scala 345:16]
  assign rvclkhdr_545_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_545_io_en = _T_6513 | _T_6518; // @[lib.scala 345:16]
  assign rvclkhdr_546_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_546_io_en = _T_6524 | _T_6529; // @[lib.scala 345:16]
  assign rvclkhdr_547_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_547_io_en = _T_6535 | _T_6540; // @[lib.scala 345:16]
  assign rvclkhdr_548_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_548_io_en = _T_6546 | _T_6551; // @[lib.scala 345:16]
  assign rvclkhdr_549_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_549_io_en = _T_6557 | _T_6562; // @[lib.scala 345:16]
  assign rvclkhdr_550_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_550_io_en = _T_6568 | _T_6573; // @[lib.scala 345:16]
  assign rvclkhdr_551_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_551_io_en = _T_6579 | _T_6584; // @[lib.scala 345:16]
  assign rvclkhdr_552_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_552_io_en = _T_6590 | _T_6595; // @[lib.scala 345:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_0 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_1 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_2 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_3 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_4 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_5 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_6 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_7 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_8 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_9 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_10 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_11 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_12 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_13 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_14 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_15 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_16 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_17 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_18 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_19 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_20 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_21 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_22 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_23 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_24 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_25 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_26 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_27 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_28 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_29 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_30 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_31 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_32 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_33 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_34 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_35 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_36 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_37 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_38 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_39 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_40 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_41 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_42 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_43 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_44 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_45 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_46 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_47 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_48 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_49 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_50 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_51 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_52 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_53 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_54 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_55 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_56 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_57 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_58 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_59 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_60 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_61 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_62 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_63 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_64 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_65 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_66 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_67 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_68 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_69 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_70 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_71 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_72 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_73 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_74 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_75 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_76 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_77 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_78 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_79 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_80 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_81 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_82 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_83 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_84 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_85 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_86 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_87 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_88 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_89 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_90 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_91 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_92 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_93 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_94 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_95 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_96 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_97 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_98 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_99 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_100 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_101 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_102 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_103 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_104 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_105 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_106 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_107 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_108 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_109 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_110 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_111 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_112 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_113 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_114 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_115 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_116 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_117 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_118 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_119 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_120 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_121 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_122 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_123 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_124 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_125 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_126 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_127 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_128 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_129 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_130 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_131 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_132 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_133 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_134 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_135 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_136 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_137 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_138 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_139 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_140 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_141 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_142 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_143 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_144 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_145 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_146 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_147 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_148 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_149 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_150 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_151 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_152 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_153 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_154 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_155 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_156 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_157 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_158 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_159 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_160 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_161 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_162 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_163 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_164 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_165 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_166 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_167 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_168 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_169 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_170 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_171 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_172 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_173 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_174 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_175 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_176 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_177 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_178 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_179 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_180 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_181 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_182 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_183 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_184 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_185 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_186 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_187 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_188 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_189 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_190 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_191 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_192 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_193 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_194 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_195 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_196 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_197 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_198 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_199 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_200 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_201 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_202 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_203 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_204 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_205 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_206 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_207 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_208 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_209 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_210 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_211 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_212 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_213 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_214 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_215 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_216 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_217 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_218 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_219 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_220 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_221 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_222 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_223 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_224 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_225 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_226 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_227 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_228 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_229 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_230 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_231 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_232 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_233 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_234 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_235 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_236 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_237 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_238 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_239 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_240 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_241 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_242 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_243 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_244 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_245 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_246 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_247 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_248 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_249 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_250 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_251 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_252 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_253 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_254 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_255 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_0 = _RAND_257[21:0];
  _RAND_258 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_1 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_2 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_3 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_4 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_5 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_6 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_7 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_8 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_9 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_10 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_11 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_12 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_13 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_14 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_15 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_16 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_17 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_18 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_19 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_20 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_21 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_22 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_23 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_24 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_25 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_26 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_27 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_28 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_29 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_30 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_31 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_32 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_33 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_34 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_35 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_36 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_37 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_38 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_39 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_40 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_41 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_42 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_43 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_44 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_45 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_46 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_47 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_48 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_49 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_50 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_51 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_52 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_53 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_54 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_55 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_56 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_57 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_58 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_59 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_60 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_61 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_62 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_63 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_64 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_65 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_66 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_67 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_68 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_69 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_70 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_71 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_72 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_73 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_74 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_75 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_76 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_77 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_78 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_79 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_80 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_81 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_82 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_83 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_84 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_85 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_86 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_87 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_88 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_89 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_90 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_91 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_92 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_93 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_94 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_95 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_96 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_97 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_98 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_99 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_100 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_101 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_102 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_103 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_104 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_105 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_106 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_107 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_108 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_109 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_110 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_111 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_112 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_113 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_114 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_115 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_116 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_117 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_118 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_119 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_120 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_121 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_122 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_123 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_124 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_125 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_126 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_127 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_128 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_129 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_130 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_131 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_132 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_133 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_134 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_135 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_136 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_137 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_138 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_139 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_140 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_141 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_142 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_143 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_144 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_145 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_146 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_147 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_148 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_149 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_150 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_151 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_152 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_153 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_154 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_155 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_156 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_157 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_158 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_159 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_160 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_161 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_162 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_163 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_164 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_165 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_166 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_167 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_168 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_169 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_170 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_171 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_172 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_173 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_174 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_175 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_176 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_177 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_178 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_179 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_180 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_181 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_182 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_183 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_184 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_185 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_186 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_187 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_188 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_189 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_190 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_191 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_192 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_193 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_194 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_195 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_196 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_197 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_198 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_199 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_200 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_201 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_202 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_203 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_204 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_205 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_206 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_207 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_208 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_209 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_210 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_211 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_212 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_213 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_214 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_215 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_216 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_217 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_218 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_219 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_220 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_221 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_222 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_223 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_224 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_225 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_226 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_227 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_228 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_229 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_230 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_231 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_232 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_233 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_234 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_235 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_236 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_237 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_238 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_239 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_240 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_241 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_242 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_243 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_244 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_245 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_246 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_247 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_248 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_249 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_250 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_251 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_252 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_253 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_254 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_255 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  fghr = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1026[0:0];
  _RAND_1027 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1027[255:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1029[29:0];
  _RAND_1030 = {1{`RANDOM}};
  rets_out_0 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_1 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_2 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_3 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_4 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_5 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_6 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_7 = _RAND_1037[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    leak_one_f_d1 = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_255 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_255 = 22'h0;
  end
  if (reset) begin
    fghr = 8'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_255 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_255 = 2'h0;
  end
  if (reset) begin
    exu_mp_way_f = 1'h0;
  end
  if (reset) begin
    btb_lru_b0_f = 256'h0;
  end
  if (reset) begin
    exu_flush_final_d1 = 1'h0;
  end
  if (reset) begin
    ifc_fetch_adder_prior = 30'h0;
  end
  if (reset) begin
    rets_out_0 = 32'h0;
  end
  if (reset) begin
    rets_out_1 = 32'h0;
  end
  if (reset) begin
    rets_out_2 = 32'h0;
  end
  if (reset) begin
    rets_out_3 = 32'h0;
  end
  if (reset) begin
    rets_out_4 = 32'h0;
  end
  if (reset) begin
    rets_out_5 = 32'h0;
  end
  if (reset) begin
    rets_out_6 = 32'h0;
  end
  if (reset) begin
    rets_out_7 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else if (_T_337) begin
      leak_one_f_d1 <= leak_one_f;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_0 <= 22'h0;
    end else if (_T_614) begin
      btb_bank0_rd_data_way0_out_0 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_1 <= 22'h0;
    end else if (_T_617) begin
      btb_bank0_rd_data_way0_out_1 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_2 <= 22'h0;
    end else if (_T_620) begin
      btb_bank0_rd_data_way0_out_2 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_3 <= 22'h0;
    end else if (_T_623) begin
      btb_bank0_rd_data_way0_out_3 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_4 <= 22'h0;
    end else if (_T_626) begin
      btb_bank0_rd_data_way0_out_4 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_5 <= 22'h0;
    end else if (_T_629) begin
      btb_bank0_rd_data_way0_out_5 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_6 <= 22'h0;
    end else if (_T_632) begin
      btb_bank0_rd_data_way0_out_6 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_7 <= 22'h0;
    end else if (_T_635) begin
      btb_bank0_rd_data_way0_out_7 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_8 <= 22'h0;
    end else if (_T_638) begin
      btb_bank0_rd_data_way0_out_8 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_9 <= 22'h0;
    end else if (_T_641) begin
      btb_bank0_rd_data_way0_out_9 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_10 <= 22'h0;
    end else if (_T_644) begin
      btb_bank0_rd_data_way0_out_10 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_11 <= 22'h0;
    end else if (_T_647) begin
      btb_bank0_rd_data_way0_out_11 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_12 <= 22'h0;
    end else if (_T_650) begin
      btb_bank0_rd_data_way0_out_12 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_13 <= 22'h0;
    end else if (_T_653) begin
      btb_bank0_rd_data_way0_out_13 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_14 <= 22'h0;
    end else if (_T_656) begin
      btb_bank0_rd_data_way0_out_14 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_15 <= 22'h0;
    end else if (_T_659) begin
      btb_bank0_rd_data_way0_out_15 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_16 <= 22'h0;
    end else if (_T_662) begin
      btb_bank0_rd_data_way0_out_16 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_17 <= 22'h0;
    end else if (_T_665) begin
      btb_bank0_rd_data_way0_out_17 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_18 <= 22'h0;
    end else if (_T_668) begin
      btb_bank0_rd_data_way0_out_18 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_19 <= 22'h0;
    end else if (_T_671) begin
      btb_bank0_rd_data_way0_out_19 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_20 <= 22'h0;
    end else if (_T_674) begin
      btb_bank0_rd_data_way0_out_20 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_21 <= 22'h0;
    end else if (_T_677) begin
      btb_bank0_rd_data_way0_out_21 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_22 <= 22'h0;
    end else if (_T_680) begin
      btb_bank0_rd_data_way0_out_22 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_23 <= 22'h0;
    end else if (_T_683) begin
      btb_bank0_rd_data_way0_out_23 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_24 <= 22'h0;
    end else if (_T_686) begin
      btb_bank0_rd_data_way0_out_24 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_25 <= 22'h0;
    end else if (_T_689) begin
      btb_bank0_rd_data_way0_out_25 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_26 <= 22'h0;
    end else if (_T_692) begin
      btb_bank0_rd_data_way0_out_26 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_27 <= 22'h0;
    end else if (_T_695) begin
      btb_bank0_rd_data_way0_out_27 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_28 <= 22'h0;
    end else if (_T_698) begin
      btb_bank0_rd_data_way0_out_28 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_29 <= 22'h0;
    end else if (_T_701) begin
      btb_bank0_rd_data_way0_out_29 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_30 <= 22'h0;
    end else if (_T_704) begin
      btb_bank0_rd_data_way0_out_30 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_31 <= 22'h0;
    end else if (_T_707) begin
      btb_bank0_rd_data_way0_out_31 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_32 <= 22'h0;
    end else if (_T_710) begin
      btb_bank0_rd_data_way0_out_32 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_33 <= 22'h0;
    end else if (_T_713) begin
      btb_bank0_rd_data_way0_out_33 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_34 <= 22'h0;
    end else if (_T_716) begin
      btb_bank0_rd_data_way0_out_34 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_35 <= 22'h0;
    end else if (_T_719) begin
      btb_bank0_rd_data_way0_out_35 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_36 <= 22'h0;
    end else if (_T_722) begin
      btb_bank0_rd_data_way0_out_36 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_37 <= 22'h0;
    end else if (_T_725) begin
      btb_bank0_rd_data_way0_out_37 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_38 <= 22'h0;
    end else if (_T_728) begin
      btb_bank0_rd_data_way0_out_38 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_39 <= 22'h0;
    end else if (_T_731) begin
      btb_bank0_rd_data_way0_out_39 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_40 <= 22'h0;
    end else if (_T_734) begin
      btb_bank0_rd_data_way0_out_40 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_41 <= 22'h0;
    end else if (_T_737) begin
      btb_bank0_rd_data_way0_out_41 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_42 <= 22'h0;
    end else if (_T_740) begin
      btb_bank0_rd_data_way0_out_42 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_43 <= 22'h0;
    end else if (_T_743) begin
      btb_bank0_rd_data_way0_out_43 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_44 <= 22'h0;
    end else if (_T_746) begin
      btb_bank0_rd_data_way0_out_44 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_45 <= 22'h0;
    end else if (_T_749) begin
      btb_bank0_rd_data_way0_out_45 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_46 <= 22'h0;
    end else if (_T_752) begin
      btb_bank0_rd_data_way0_out_46 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_47 <= 22'h0;
    end else if (_T_755) begin
      btb_bank0_rd_data_way0_out_47 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_48 <= 22'h0;
    end else if (_T_758) begin
      btb_bank0_rd_data_way0_out_48 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_49 <= 22'h0;
    end else if (_T_761) begin
      btb_bank0_rd_data_way0_out_49 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_50 <= 22'h0;
    end else if (_T_764) begin
      btb_bank0_rd_data_way0_out_50 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_51 <= 22'h0;
    end else if (_T_767) begin
      btb_bank0_rd_data_way0_out_51 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_52 <= 22'h0;
    end else if (_T_770) begin
      btb_bank0_rd_data_way0_out_52 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_53 <= 22'h0;
    end else if (_T_773) begin
      btb_bank0_rd_data_way0_out_53 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_54 <= 22'h0;
    end else if (_T_776) begin
      btb_bank0_rd_data_way0_out_54 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_55 <= 22'h0;
    end else if (_T_779) begin
      btb_bank0_rd_data_way0_out_55 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_56 <= 22'h0;
    end else if (_T_782) begin
      btb_bank0_rd_data_way0_out_56 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_57 <= 22'h0;
    end else if (_T_785) begin
      btb_bank0_rd_data_way0_out_57 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_58 <= 22'h0;
    end else if (_T_788) begin
      btb_bank0_rd_data_way0_out_58 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_59 <= 22'h0;
    end else if (_T_791) begin
      btb_bank0_rd_data_way0_out_59 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_60 <= 22'h0;
    end else if (_T_794) begin
      btb_bank0_rd_data_way0_out_60 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_61 <= 22'h0;
    end else if (_T_797) begin
      btb_bank0_rd_data_way0_out_61 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_62 <= 22'h0;
    end else if (_T_800) begin
      btb_bank0_rd_data_way0_out_62 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_63 <= 22'h0;
    end else if (_T_803) begin
      btb_bank0_rd_data_way0_out_63 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_64 <= 22'h0;
    end else if (_T_806) begin
      btb_bank0_rd_data_way0_out_64 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_65 <= 22'h0;
    end else if (_T_809) begin
      btb_bank0_rd_data_way0_out_65 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_66 <= 22'h0;
    end else if (_T_812) begin
      btb_bank0_rd_data_way0_out_66 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_67 <= 22'h0;
    end else if (_T_815) begin
      btb_bank0_rd_data_way0_out_67 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_68 <= 22'h0;
    end else if (_T_818) begin
      btb_bank0_rd_data_way0_out_68 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_69 <= 22'h0;
    end else if (_T_821) begin
      btb_bank0_rd_data_way0_out_69 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_70 <= 22'h0;
    end else if (_T_824) begin
      btb_bank0_rd_data_way0_out_70 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_71 <= 22'h0;
    end else if (_T_827) begin
      btb_bank0_rd_data_way0_out_71 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_72 <= 22'h0;
    end else if (_T_830) begin
      btb_bank0_rd_data_way0_out_72 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_73 <= 22'h0;
    end else if (_T_833) begin
      btb_bank0_rd_data_way0_out_73 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_74 <= 22'h0;
    end else if (_T_836) begin
      btb_bank0_rd_data_way0_out_74 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_75 <= 22'h0;
    end else if (_T_839) begin
      btb_bank0_rd_data_way0_out_75 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_76 <= 22'h0;
    end else if (_T_842) begin
      btb_bank0_rd_data_way0_out_76 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_77 <= 22'h0;
    end else if (_T_845) begin
      btb_bank0_rd_data_way0_out_77 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_78 <= 22'h0;
    end else if (_T_848) begin
      btb_bank0_rd_data_way0_out_78 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_79 <= 22'h0;
    end else if (_T_851) begin
      btb_bank0_rd_data_way0_out_79 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_80 <= 22'h0;
    end else if (_T_854) begin
      btb_bank0_rd_data_way0_out_80 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_81 <= 22'h0;
    end else if (_T_857) begin
      btb_bank0_rd_data_way0_out_81 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_82 <= 22'h0;
    end else if (_T_860) begin
      btb_bank0_rd_data_way0_out_82 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_83 <= 22'h0;
    end else if (_T_863) begin
      btb_bank0_rd_data_way0_out_83 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_84 <= 22'h0;
    end else if (_T_866) begin
      btb_bank0_rd_data_way0_out_84 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_85 <= 22'h0;
    end else if (_T_869) begin
      btb_bank0_rd_data_way0_out_85 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_86 <= 22'h0;
    end else if (_T_872) begin
      btb_bank0_rd_data_way0_out_86 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_87 <= 22'h0;
    end else if (_T_875) begin
      btb_bank0_rd_data_way0_out_87 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_88 <= 22'h0;
    end else if (_T_878) begin
      btb_bank0_rd_data_way0_out_88 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_89 <= 22'h0;
    end else if (_T_881) begin
      btb_bank0_rd_data_way0_out_89 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_90 <= 22'h0;
    end else if (_T_884) begin
      btb_bank0_rd_data_way0_out_90 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_91 <= 22'h0;
    end else if (_T_887) begin
      btb_bank0_rd_data_way0_out_91 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_92 <= 22'h0;
    end else if (_T_890) begin
      btb_bank0_rd_data_way0_out_92 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_93 <= 22'h0;
    end else if (_T_893) begin
      btb_bank0_rd_data_way0_out_93 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_94 <= 22'h0;
    end else if (_T_896) begin
      btb_bank0_rd_data_way0_out_94 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_95 <= 22'h0;
    end else if (_T_899) begin
      btb_bank0_rd_data_way0_out_95 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_96 <= 22'h0;
    end else if (_T_902) begin
      btb_bank0_rd_data_way0_out_96 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_97 <= 22'h0;
    end else if (_T_905) begin
      btb_bank0_rd_data_way0_out_97 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_98 <= 22'h0;
    end else if (_T_908) begin
      btb_bank0_rd_data_way0_out_98 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_99 <= 22'h0;
    end else if (_T_911) begin
      btb_bank0_rd_data_way0_out_99 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_100 <= 22'h0;
    end else if (_T_914) begin
      btb_bank0_rd_data_way0_out_100 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_101 <= 22'h0;
    end else if (_T_917) begin
      btb_bank0_rd_data_way0_out_101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_102 <= 22'h0;
    end else if (_T_920) begin
      btb_bank0_rd_data_way0_out_102 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_103 <= 22'h0;
    end else if (_T_923) begin
      btb_bank0_rd_data_way0_out_103 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_104 <= 22'h0;
    end else if (_T_926) begin
      btb_bank0_rd_data_way0_out_104 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_105 <= 22'h0;
    end else if (_T_929) begin
      btb_bank0_rd_data_way0_out_105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_106 <= 22'h0;
    end else if (_T_932) begin
      btb_bank0_rd_data_way0_out_106 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_107 <= 22'h0;
    end else if (_T_935) begin
      btb_bank0_rd_data_way0_out_107 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_108 <= 22'h0;
    end else if (_T_938) begin
      btb_bank0_rd_data_way0_out_108 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_109 <= 22'h0;
    end else if (_T_941) begin
      btb_bank0_rd_data_way0_out_109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_110 <= 22'h0;
    end else if (_T_944) begin
      btb_bank0_rd_data_way0_out_110 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_111 <= 22'h0;
    end else if (_T_947) begin
      btb_bank0_rd_data_way0_out_111 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_112 <= 22'h0;
    end else if (_T_950) begin
      btb_bank0_rd_data_way0_out_112 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_113 <= 22'h0;
    end else if (_T_953) begin
      btb_bank0_rd_data_way0_out_113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_114 <= 22'h0;
    end else if (_T_956) begin
      btb_bank0_rd_data_way0_out_114 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_115 <= 22'h0;
    end else if (_T_959) begin
      btb_bank0_rd_data_way0_out_115 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_116 <= 22'h0;
    end else if (_T_962) begin
      btb_bank0_rd_data_way0_out_116 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_117 <= 22'h0;
    end else if (_T_965) begin
      btb_bank0_rd_data_way0_out_117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_118 <= 22'h0;
    end else if (_T_968) begin
      btb_bank0_rd_data_way0_out_118 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_119 <= 22'h0;
    end else if (_T_971) begin
      btb_bank0_rd_data_way0_out_119 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_120 <= 22'h0;
    end else if (_T_974) begin
      btb_bank0_rd_data_way0_out_120 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_121 <= 22'h0;
    end else if (_T_977) begin
      btb_bank0_rd_data_way0_out_121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_122 <= 22'h0;
    end else if (_T_980) begin
      btb_bank0_rd_data_way0_out_122 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_123 <= 22'h0;
    end else if (_T_983) begin
      btb_bank0_rd_data_way0_out_123 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_124 <= 22'h0;
    end else if (_T_986) begin
      btb_bank0_rd_data_way0_out_124 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_125 <= 22'h0;
    end else if (_T_989) begin
      btb_bank0_rd_data_way0_out_125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_126 <= 22'h0;
    end else if (_T_992) begin
      btb_bank0_rd_data_way0_out_126 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_127 <= 22'h0;
    end else if (_T_995) begin
      btb_bank0_rd_data_way0_out_127 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_128 <= 22'h0;
    end else if (_T_998) begin
      btb_bank0_rd_data_way0_out_128 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_129 <= 22'h0;
    end else if (_T_1001) begin
      btb_bank0_rd_data_way0_out_129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_130 <= 22'h0;
    end else if (_T_1004) begin
      btb_bank0_rd_data_way0_out_130 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_131 <= 22'h0;
    end else if (_T_1007) begin
      btb_bank0_rd_data_way0_out_131 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_132 <= 22'h0;
    end else if (_T_1010) begin
      btb_bank0_rd_data_way0_out_132 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_133 <= 22'h0;
    end else if (_T_1013) begin
      btb_bank0_rd_data_way0_out_133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_134 <= 22'h0;
    end else if (_T_1016) begin
      btb_bank0_rd_data_way0_out_134 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_135 <= 22'h0;
    end else if (_T_1019) begin
      btb_bank0_rd_data_way0_out_135 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_136 <= 22'h0;
    end else if (_T_1022) begin
      btb_bank0_rd_data_way0_out_136 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_137 <= 22'h0;
    end else if (_T_1025) begin
      btb_bank0_rd_data_way0_out_137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_138 <= 22'h0;
    end else if (_T_1028) begin
      btb_bank0_rd_data_way0_out_138 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_139 <= 22'h0;
    end else if (_T_1031) begin
      btb_bank0_rd_data_way0_out_139 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_140 <= 22'h0;
    end else if (_T_1034) begin
      btb_bank0_rd_data_way0_out_140 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_141 <= 22'h0;
    end else if (_T_1037) begin
      btb_bank0_rd_data_way0_out_141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_142 <= 22'h0;
    end else if (_T_1040) begin
      btb_bank0_rd_data_way0_out_142 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_143 <= 22'h0;
    end else if (_T_1043) begin
      btb_bank0_rd_data_way0_out_143 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_144 <= 22'h0;
    end else if (_T_1046) begin
      btb_bank0_rd_data_way0_out_144 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_145 <= 22'h0;
    end else if (_T_1049) begin
      btb_bank0_rd_data_way0_out_145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_146 <= 22'h0;
    end else if (_T_1052) begin
      btb_bank0_rd_data_way0_out_146 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_147 <= 22'h0;
    end else if (_T_1055) begin
      btb_bank0_rd_data_way0_out_147 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_148 <= 22'h0;
    end else if (_T_1058) begin
      btb_bank0_rd_data_way0_out_148 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_149 <= 22'h0;
    end else if (_T_1061) begin
      btb_bank0_rd_data_way0_out_149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_150 <= 22'h0;
    end else if (_T_1064) begin
      btb_bank0_rd_data_way0_out_150 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_151 <= 22'h0;
    end else if (_T_1067) begin
      btb_bank0_rd_data_way0_out_151 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_152 <= 22'h0;
    end else if (_T_1070) begin
      btb_bank0_rd_data_way0_out_152 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_153 <= 22'h0;
    end else if (_T_1073) begin
      btb_bank0_rd_data_way0_out_153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_154 <= 22'h0;
    end else if (_T_1076) begin
      btb_bank0_rd_data_way0_out_154 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_155 <= 22'h0;
    end else if (_T_1079) begin
      btb_bank0_rd_data_way0_out_155 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_156 <= 22'h0;
    end else if (_T_1082) begin
      btb_bank0_rd_data_way0_out_156 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_157 <= 22'h0;
    end else if (_T_1085) begin
      btb_bank0_rd_data_way0_out_157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_158 <= 22'h0;
    end else if (_T_1088) begin
      btb_bank0_rd_data_way0_out_158 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_159 <= 22'h0;
    end else if (_T_1091) begin
      btb_bank0_rd_data_way0_out_159 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_160 <= 22'h0;
    end else if (_T_1094) begin
      btb_bank0_rd_data_way0_out_160 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_161 <= 22'h0;
    end else if (_T_1097) begin
      btb_bank0_rd_data_way0_out_161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_162 <= 22'h0;
    end else if (_T_1100) begin
      btb_bank0_rd_data_way0_out_162 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_163 <= 22'h0;
    end else if (_T_1103) begin
      btb_bank0_rd_data_way0_out_163 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_164 <= 22'h0;
    end else if (_T_1106) begin
      btb_bank0_rd_data_way0_out_164 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_165 <= 22'h0;
    end else if (_T_1109) begin
      btb_bank0_rd_data_way0_out_165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_166 <= 22'h0;
    end else if (_T_1112) begin
      btb_bank0_rd_data_way0_out_166 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_167 <= 22'h0;
    end else if (_T_1115) begin
      btb_bank0_rd_data_way0_out_167 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_168 <= 22'h0;
    end else if (_T_1118) begin
      btb_bank0_rd_data_way0_out_168 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_169 <= 22'h0;
    end else if (_T_1121) begin
      btb_bank0_rd_data_way0_out_169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_170 <= 22'h0;
    end else if (_T_1124) begin
      btb_bank0_rd_data_way0_out_170 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_171 <= 22'h0;
    end else if (_T_1127) begin
      btb_bank0_rd_data_way0_out_171 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_172 <= 22'h0;
    end else if (_T_1130) begin
      btb_bank0_rd_data_way0_out_172 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_173 <= 22'h0;
    end else if (_T_1133) begin
      btb_bank0_rd_data_way0_out_173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_174 <= 22'h0;
    end else if (_T_1136) begin
      btb_bank0_rd_data_way0_out_174 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_175 <= 22'h0;
    end else if (_T_1139) begin
      btb_bank0_rd_data_way0_out_175 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_176 <= 22'h0;
    end else if (_T_1142) begin
      btb_bank0_rd_data_way0_out_176 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_177 <= 22'h0;
    end else if (_T_1145) begin
      btb_bank0_rd_data_way0_out_177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_178 <= 22'h0;
    end else if (_T_1148) begin
      btb_bank0_rd_data_way0_out_178 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_179 <= 22'h0;
    end else if (_T_1151) begin
      btb_bank0_rd_data_way0_out_179 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_180 <= 22'h0;
    end else if (_T_1154) begin
      btb_bank0_rd_data_way0_out_180 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_181 <= 22'h0;
    end else if (_T_1157) begin
      btb_bank0_rd_data_way0_out_181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_182 <= 22'h0;
    end else if (_T_1160) begin
      btb_bank0_rd_data_way0_out_182 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_183 <= 22'h0;
    end else if (_T_1163) begin
      btb_bank0_rd_data_way0_out_183 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_184 <= 22'h0;
    end else if (_T_1166) begin
      btb_bank0_rd_data_way0_out_184 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_185 <= 22'h0;
    end else if (_T_1169) begin
      btb_bank0_rd_data_way0_out_185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_186 <= 22'h0;
    end else if (_T_1172) begin
      btb_bank0_rd_data_way0_out_186 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_187 <= 22'h0;
    end else if (_T_1175) begin
      btb_bank0_rd_data_way0_out_187 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_188 <= 22'h0;
    end else if (_T_1178) begin
      btb_bank0_rd_data_way0_out_188 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_189 <= 22'h0;
    end else if (_T_1181) begin
      btb_bank0_rd_data_way0_out_189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_190 <= 22'h0;
    end else if (_T_1184) begin
      btb_bank0_rd_data_way0_out_190 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_191 <= 22'h0;
    end else if (_T_1187) begin
      btb_bank0_rd_data_way0_out_191 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_192 <= 22'h0;
    end else if (_T_1190) begin
      btb_bank0_rd_data_way0_out_192 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_193 <= 22'h0;
    end else if (_T_1193) begin
      btb_bank0_rd_data_way0_out_193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_194 <= 22'h0;
    end else if (_T_1196) begin
      btb_bank0_rd_data_way0_out_194 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_195 <= 22'h0;
    end else if (_T_1199) begin
      btb_bank0_rd_data_way0_out_195 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_196 <= 22'h0;
    end else if (_T_1202) begin
      btb_bank0_rd_data_way0_out_196 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_197 <= 22'h0;
    end else if (_T_1205) begin
      btb_bank0_rd_data_way0_out_197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_198 <= 22'h0;
    end else if (_T_1208) begin
      btb_bank0_rd_data_way0_out_198 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_199 <= 22'h0;
    end else if (_T_1211) begin
      btb_bank0_rd_data_way0_out_199 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_200 <= 22'h0;
    end else if (_T_1214) begin
      btb_bank0_rd_data_way0_out_200 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_201 <= 22'h0;
    end else if (_T_1217) begin
      btb_bank0_rd_data_way0_out_201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_202 <= 22'h0;
    end else if (_T_1220) begin
      btb_bank0_rd_data_way0_out_202 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_203 <= 22'h0;
    end else if (_T_1223) begin
      btb_bank0_rd_data_way0_out_203 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_204 <= 22'h0;
    end else if (_T_1226) begin
      btb_bank0_rd_data_way0_out_204 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_205 <= 22'h0;
    end else if (_T_1229) begin
      btb_bank0_rd_data_way0_out_205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_206 <= 22'h0;
    end else if (_T_1232) begin
      btb_bank0_rd_data_way0_out_206 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_207 <= 22'h0;
    end else if (_T_1235) begin
      btb_bank0_rd_data_way0_out_207 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_208 <= 22'h0;
    end else if (_T_1238) begin
      btb_bank0_rd_data_way0_out_208 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_209 <= 22'h0;
    end else if (_T_1241) begin
      btb_bank0_rd_data_way0_out_209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_210 <= 22'h0;
    end else if (_T_1244) begin
      btb_bank0_rd_data_way0_out_210 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_211 <= 22'h0;
    end else if (_T_1247) begin
      btb_bank0_rd_data_way0_out_211 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_212 <= 22'h0;
    end else if (_T_1250) begin
      btb_bank0_rd_data_way0_out_212 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_213 <= 22'h0;
    end else if (_T_1253) begin
      btb_bank0_rd_data_way0_out_213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_214 <= 22'h0;
    end else if (_T_1256) begin
      btb_bank0_rd_data_way0_out_214 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_215 <= 22'h0;
    end else if (_T_1259) begin
      btb_bank0_rd_data_way0_out_215 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_216 <= 22'h0;
    end else if (_T_1262) begin
      btb_bank0_rd_data_way0_out_216 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_217 <= 22'h0;
    end else if (_T_1265) begin
      btb_bank0_rd_data_way0_out_217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_218 <= 22'h0;
    end else if (_T_1268) begin
      btb_bank0_rd_data_way0_out_218 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_219 <= 22'h0;
    end else if (_T_1271) begin
      btb_bank0_rd_data_way0_out_219 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_220 <= 22'h0;
    end else if (_T_1274) begin
      btb_bank0_rd_data_way0_out_220 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_221 <= 22'h0;
    end else if (_T_1277) begin
      btb_bank0_rd_data_way0_out_221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_222 <= 22'h0;
    end else if (_T_1280) begin
      btb_bank0_rd_data_way0_out_222 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_223 <= 22'h0;
    end else if (_T_1283) begin
      btb_bank0_rd_data_way0_out_223 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_224 <= 22'h0;
    end else if (_T_1286) begin
      btb_bank0_rd_data_way0_out_224 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_225 <= 22'h0;
    end else if (_T_1289) begin
      btb_bank0_rd_data_way0_out_225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_226 <= 22'h0;
    end else if (_T_1292) begin
      btb_bank0_rd_data_way0_out_226 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_227 <= 22'h0;
    end else if (_T_1295) begin
      btb_bank0_rd_data_way0_out_227 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_228 <= 22'h0;
    end else if (_T_1298) begin
      btb_bank0_rd_data_way0_out_228 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_229 <= 22'h0;
    end else if (_T_1301) begin
      btb_bank0_rd_data_way0_out_229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_230 <= 22'h0;
    end else if (_T_1304) begin
      btb_bank0_rd_data_way0_out_230 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_231 <= 22'h0;
    end else if (_T_1307) begin
      btb_bank0_rd_data_way0_out_231 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_232 <= 22'h0;
    end else if (_T_1310) begin
      btb_bank0_rd_data_way0_out_232 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_233 <= 22'h0;
    end else if (_T_1313) begin
      btb_bank0_rd_data_way0_out_233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_234 <= 22'h0;
    end else if (_T_1316) begin
      btb_bank0_rd_data_way0_out_234 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_235 <= 22'h0;
    end else if (_T_1319) begin
      btb_bank0_rd_data_way0_out_235 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_236 <= 22'h0;
    end else if (_T_1322) begin
      btb_bank0_rd_data_way0_out_236 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_237 <= 22'h0;
    end else if (_T_1325) begin
      btb_bank0_rd_data_way0_out_237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_238 <= 22'h0;
    end else if (_T_1328) begin
      btb_bank0_rd_data_way0_out_238 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_239 <= 22'h0;
    end else if (_T_1331) begin
      btb_bank0_rd_data_way0_out_239 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_240 <= 22'h0;
    end else if (_T_1334) begin
      btb_bank0_rd_data_way0_out_240 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_241 <= 22'h0;
    end else if (_T_1337) begin
      btb_bank0_rd_data_way0_out_241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_242 <= 22'h0;
    end else if (_T_1340) begin
      btb_bank0_rd_data_way0_out_242 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_243 <= 22'h0;
    end else if (_T_1343) begin
      btb_bank0_rd_data_way0_out_243 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_244 <= 22'h0;
    end else if (_T_1346) begin
      btb_bank0_rd_data_way0_out_244 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_245 <= 22'h0;
    end else if (_T_1349) begin
      btb_bank0_rd_data_way0_out_245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_246 <= 22'h0;
    end else if (_T_1352) begin
      btb_bank0_rd_data_way0_out_246 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_247 <= 22'h0;
    end else if (_T_1355) begin
      btb_bank0_rd_data_way0_out_247 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_248 <= 22'h0;
    end else if (_T_1358) begin
      btb_bank0_rd_data_way0_out_248 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_249 <= 22'h0;
    end else if (_T_1361) begin
      btb_bank0_rd_data_way0_out_249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_250 <= 22'h0;
    end else if (_T_1364) begin
      btb_bank0_rd_data_way0_out_250 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_251 <= 22'h0;
    end else if (_T_1367) begin
      btb_bank0_rd_data_way0_out_251 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_252 <= 22'h0;
    end else if (_T_1370) begin
      btb_bank0_rd_data_way0_out_252 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_253 <= 22'h0;
    end else if (_T_1373) begin
      btb_bank0_rd_data_way0_out_253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_254 <= 22'h0;
    end else if (_T_1376) begin
      btb_bank0_rd_data_way0_out_254 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_255 <= 22'h0;
    end else if (_T_1379) begin
      btb_bank0_rd_data_way0_out_255 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_0 <= 22'h0;
    end else if (_T_1382) begin
      btb_bank0_rd_data_way1_out_0 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_1 <= 22'h0;
    end else if (_T_1385) begin
      btb_bank0_rd_data_way1_out_1 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_2 <= 22'h0;
    end else if (_T_1388) begin
      btb_bank0_rd_data_way1_out_2 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_3 <= 22'h0;
    end else if (_T_1391) begin
      btb_bank0_rd_data_way1_out_3 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_4 <= 22'h0;
    end else if (_T_1394) begin
      btb_bank0_rd_data_way1_out_4 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_5 <= 22'h0;
    end else if (_T_1397) begin
      btb_bank0_rd_data_way1_out_5 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_6 <= 22'h0;
    end else if (_T_1400) begin
      btb_bank0_rd_data_way1_out_6 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_7 <= 22'h0;
    end else if (_T_1403) begin
      btb_bank0_rd_data_way1_out_7 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_8 <= 22'h0;
    end else if (_T_1406) begin
      btb_bank0_rd_data_way1_out_8 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_9 <= 22'h0;
    end else if (_T_1409) begin
      btb_bank0_rd_data_way1_out_9 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_10 <= 22'h0;
    end else if (_T_1412) begin
      btb_bank0_rd_data_way1_out_10 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_11 <= 22'h0;
    end else if (_T_1415) begin
      btb_bank0_rd_data_way1_out_11 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_12 <= 22'h0;
    end else if (_T_1418) begin
      btb_bank0_rd_data_way1_out_12 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_13 <= 22'h0;
    end else if (_T_1421) begin
      btb_bank0_rd_data_way1_out_13 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_14 <= 22'h0;
    end else if (_T_1424) begin
      btb_bank0_rd_data_way1_out_14 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_15 <= 22'h0;
    end else if (_T_1427) begin
      btb_bank0_rd_data_way1_out_15 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_16 <= 22'h0;
    end else if (_T_1430) begin
      btb_bank0_rd_data_way1_out_16 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_17 <= 22'h0;
    end else if (_T_1433) begin
      btb_bank0_rd_data_way1_out_17 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_18 <= 22'h0;
    end else if (_T_1436) begin
      btb_bank0_rd_data_way1_out_18 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_19 <= 22'h0;
    end else if (_T_1439) begin
      btb_bank0_rd_data_way1_out_19 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_20 <= 22'h0;
    end else if (_T_1442) begin
      btb_bank0_rd_data_way1_out_20 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_21 <= 22'h0;
    end else if (_T_1445) begin
      btb_bank0_rd_data_way1_out_21 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_22 <= 22'h0;
    end else if (_T_1448) begin
      btb_bank0_rd_data_way1_out_22 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_23 <= 22'h0;
    end else if (_T_1451) begin
      btb_bank0_rd_data_way1_out_23 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_24 <= 22'h0;
    end else if (_T_1454) begin
      btb_bank0_rd_data_way1_out_24 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_25 <= 22'h0;
    end else if (_T_1457) begin
      btb_bank0_rd_data_way1_out_25 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_26 <= 22'h0;
    end else if (_T_1460) begin
      btb_bank0_rd_data_way1_out_26 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_27 <= 22'h0;
    end else if (_T_1463) begin
      btb_bank0_rd_data_way1_out_27 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_28 <= 22'h0;
    end else if (_T_1466) begin
      btb_bank0_rd_data_way1_out_28 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_29 <= 22'h0;
    end else if (_T_1469) begin
      btb_bank0_rd_data_way1_out_29 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_30 <= 22'h0;
    end else if (_T_1472) begin
      btb_bank0_rd_data_way1_out_30 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_31 <= 22'h0;
    end else if (_T_1475) begin
      btb_bank0_rd_data_way1_out_31 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_32 <= 22'h0;
    end else if (_T_1478) begin
      btb_bank0_rd_data_way1_out_32 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_33 <= 22'h0;
    end else if (_T_1481) begin
      btb_bank0_rd_data_way1_out_33 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_34 <= 22'h0;
    end else if (_T_1484) begin
      btb_bank0_rd_data_way1_out_34 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_35 <= 22'h0;
    end else if (_T_1487) begin
      btb_bank0_rd_data_way1_out_35 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_36 <= 22'h0;
    end else if (_T_1490) begin
      btb_bank0_rd_data_way1_out_36 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_37 <= 22'h0;
    end else if (_T_1493) begin
      btb_bank0_rd_data_way1_out_37 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_38 <= 22'h0;
    end else if (_T_1496) begin
      btb_bank0_rd_data_way1_out_38 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_39 <= 22'h0;
    end else if (_T_1499) begin
      btb_bank0_rd_data_way1_out_39 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_40 <= 22'h0;
    end else if (_T_1502) begin
      btb_bank0_rd_data_way1_out_40 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_41 <= 22'h0;
    end else if (_T_1505) begin
      btb_bank0_rd_data_way1_out_41 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_42 <= 22'h0;
    end else if (_T_1508) begin
      btb_bank0_rd_data_way1_out_42 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_43 <= 22'h0;
    end else if (_T_1511) begin
      btb_bank0_rd_data_way1_out_43 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_44 <= 22'h0;
    end else if (_T_1514) begin
      btb_bank0_rd_data_way1_out_44 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_45 <= 22'h0;
    end else if (_T_1517) begin
      btb_bank0_rd_data_way1_out_45 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_46 <= 22'h0;
    end else if (_T_1520) begin
      btb_bank0_rd_data_way1_out_46 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_47 <= 22'h0;
    end else if (_T_1523) begin
      btb_bank0_rd_data_way1_out_47 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_48 <= 22'h0;
    end else if (_T_1526) begin
      btb_bank0_rd_data_way1_out_48 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_49 <= 22'h0;
    end else if (_T_1529) begin
      btb_bank0_rd_data_way1_out_49 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_50 <= 22'h0;
    end else if (_T_1532) begin
      btb_bank0_rd_data_way1_out_50 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_51 <= 22'h0;
    end else if (_T_1535) begin
      btb_bank0_rd_data_way1_out_51 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_52 <= 22'h0;
    end else if (_T_1538) begin
      btb_bank0_rd_data_way1_out_52 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_53 <= 22'h0;
    end else if (_T_1541) begin
      btb_bank0_rd_data_way1_out_53 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_54 <= 22'h0;
    end else if (_T_1544) begin
      btb_bank0_rd_data_way1_out_54 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_55 <= 22'h0;
    end else if (_T_1547) begin
      btb_bank0_rd_data_way1_out_55 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_56 <= 22'h0;
    end else if (_T_1550) begin
      btb_bank0_rd_data_way1_out_56 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_57 <= 22'h0;
    end else if (_T_1553) begin
      btb_bank0_rd_data_way1_out_57 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_58 <= 22'h0;
    end else if (_T_1556) begin
      btb_bank0_rd_data_way1_out_58 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_59 <= 22'h0;
    end else if (_T_1559) begin
      btb_bank0_rd_data_way1_out_59 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_60 <= 22'h0;
    end else if (_T_1562) begin
      btb_bank0_rd_data_way1_out_60 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_61 <= 22'h0;
    end else if (_T_1565) begin
      btb_bank0_rd_data_way1_out_61 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_62 <= 22'h0;
    end else if (_T_1568) begin
      btb_bank0_rd_data_way1_out_62 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_63 <= 22'h0;
    end else if (_T_1571) begin
      btb_bank0_rd_data_way1_out_63 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_64 <= 22'h0;
    end else if (_T_1574) begin
      btb_bank0_rd_data_way1_out_64 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_65 <= 22'h0;
    end else if (_T_1577) begin
      btb_bank0_rd_data_way1_out_65 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_66 <= 22'h0;
    end else if (_T_1580) begin
      btb_bank0_rd_data_way1_out_66 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_67 <= 22'h0;
    end else if (_T_1583) begin
      btb_bank0_rd_data_way1_out_67 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_68 <= 22'h0;
    end else if (_T_1586) begin
      btb_bank0_rd_data_way1_out_68 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_69 <= 22'h0;
    end else if (_T_1589) begin
      btb_bank0_rd_data_way1_out_69 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_70 <= 22'h0;
    end else if (_T_1592) begin
      btb_bank0_rd_data_way1_out_70 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_71 <= 22'h0;
    end else if (_T_1595) begin
      btb_bank0_rd_data_way1_out_71 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_72 <= 22'h0;
    end else if (_T_1598) begin
      btb_bank0_rd_data_way1_out_72 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_73 <= 22'h0;
    end else if (_T_1601) begin
      btb_bank0_rd_data_way1_out_73 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_74 <= 22'h0;
    end else if (_T_1604) begin
      btb_bank0_rd_data_way1_out_74 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_75 <= 22'h0;
    end else if (_T_1607) begin
      btb_bank0_rd_data_way1_out_75 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_76 <= 22'h0;
    end else if (_T_1610) begin
      btb_bank0_rd_data_way1_out_76 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_77 <= 22'h0;
    end else if (_T_1613) begin
      btb_bank0_rd_data_way1_out_77 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_78 <= 22'h0;
    end else if (_T_1616) begin
      btb_bank0_rd_data_way1_out_78 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_79 <= 22'h0;
    end else if (_T_1619) begin
      btb_bank0_rd_data_way1_out_79 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_80 <= 22'h0;
    end else if (_T_1622) begin
      btb_bank0_rd_data_way1_out_80 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_81 <= 22'h0;
    end else if (_T_1625) begin
      btb_bank0_rd_data_way1_out_81 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_82 <= 22'h0;
    end else if (_T_1628) begin
      btb_bank0_rd_data_way1_out_82 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_83 <= 22'h0;
    end else if (_T_1631) begin
      btb_bank0_rd_data_way1_out_83 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_84 <= 22'h0;
    end else if (_T_1634) begin
      btb_bank0_rd_data_way1_out_84 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_85 <= 22'h0;
    end else if (_T_1637) begin
      btb_bank0_rd_data_way1_out_85 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_86 <= 22'h0;
    end else if (_T_1640) begin
      btb_bank0_rd_data_way1_out_86 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_87 <= 22'h0;
    end else if (_T_1643) begin
      btb_bank0_rd_data_way1_out_87 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_88 <= 22'h0;
    end else if (_T_1646) begin
      btb_bank0_rd_data_way1_out_88 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_89 <= 22'h0;
    end else if (_T_1649) begin
      btb_bank0_rd_data_way1_out_89 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_90 <= 22'h0;
    end else if (_T_1652) begin
      btb_bank0_rd_data_way1_out_90 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_91 <= 22'h0;
    end else if (_T_1655) begin
      btb_bank0_rd_data_way1_out_91 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_92 <= 22'h0;
    end else if (_T_1658) begin
      btb_bank0_rd_data_way1_out_92 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_93 <= 22'h0;
    end else if (_T_1661) begin
      btb_bank0_rd_data_way1_out_93 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_94 <= 22'h0;
    end else if (_T_1664) begin
      btb_bank0_rd_data_way1_out_94 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_95 <= 22'h0;
    end else if (_T_1667) begin
      btb_bank0_rd_data_way1_out_95 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_96 <= 22'h0;
    end else if (_T_1670) begin
      btb_bank0_rd_data_way1_out_96 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_97 <= 22'h0;
    end else if (_T_1673) begin
      btb_bank0_rd_data_way1_out_97 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_98 <= 22'h0;
    end else if (_T_1676) begin
      btb_bank0_rd_data_way1_out_98 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_99 <= 22'h0;
    end else if (_T_1679) begin
      btb_bank0_rd_data_way1_out_99 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_100 <= 22'h0;
    end else if (_T_1682) begin
      btb_bank0_rd_data_way1_out_100 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_101 <= 22'h0;
    end else if (_T_1685) begin
      btb_bank0_rd_data_way1_out_101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_102 <= 22'h0;
    end else if (_T_1688) begin
      btb_bank0_rd_data_way1_out_102 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_103 <= 22'h0;
    end else if (_T_1691) begin
      btb_bank0_rd_data_way1_out_103 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_104 <= 22'h0;
    end else if (_T_1694) begin
      btb_bank0_rd_data_way1_out_104 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_105 <= 22'h0;
    end else if (_T_1697) begin
      btb_bank0_rd_data_way1_out_105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_106 <= 22'h0;
    end else if (_T_1700) begin
      btb_bank0_rd_data_way1_out_106 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_107 <= 22'h0;
    end else if (_T_1703) begin
      btb_bank0_rd_data_way1_out_107 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_108 <= 22'h0;
    end else if (_T_1706) begin
      btb_bank0_rd_data_way1_out_108 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_109 <= 22'h0;
    end else if (_T_1709) begin
      btb_bank0_rd_data_way1_out_109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_110 <= 22'h0;
    end else if (_T_1712) begin
      btb_bank0_rd_data_way1_out_110 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_111 <= 22'h0;
    end else if (_T_1715) begin
      btb_bank0_rd_data_way1_out_111 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_112 <= 22'h0;
    end else if (_T_1718) begin
      btb_bank0_rd_data_way1_out_112 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_113 <= 22'h0;
    end else if (_T_1721) begin
      btb_bank0_rd_data_way1_out_113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_114 <= 22'h0;
    end else if (_T_1724) begin
      btb_bank0_rd_data_way1_out_114 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_115 <= 22'h0;
    end else if (_T_1727) begin
      btb_bank0_rd_data_way1_out_115 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_116 <= 22'h0;
    end else if (_T_1730) begin
      btb_bank0_rd_data_way1_out_116 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_117 <= 22'h0;
    end else if (_T_1733) begin
      btb_bank0_rd_data_way1_out_117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_118 <= 22'h0;
    end else if (_T_1736) begin
      btb_bank0_rd_data_way1_out_118 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_119 <= 22'h0;
    end else if (_T_1739) begin
      btb_bank0_rd_data_way1_out_119 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_120 <= 22'h0;
    end else if (_T_1742) begin
      btb_bank0_rd_data_way1_out_120 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_121 <= 22'h0;
    end else if (_T_1745) begin
      btb_bank0_rd_data_way1_out_121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_122 <= 22'h0;
    end else if (_T_1748) begin
      btb_bank0_rd_data_way1_out_122 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_123 <= 22'h0;
    end else if (_T_1751) begin
      btb_bank0_rd_data_way1_out_123 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_124 <= 22'h0;
    end else if (_T_1754) begin
      btb_bank0_rd_data_way1_out_124 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_125 <= 22'h0;
    end else if (_T_1757) begin
      btb_bank0_rd_data_way1_out_125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_126 <= 22'h0;
    end else if (_T_1760) begin
      btb_bank0_rd_data_way1_out_126 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_127 <= 22'h0;
    end else if (_T_1763) begin
      btb_bank0_rd_data_way1_out_127 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_128 <= 22'h0;
    end else if (_T_1766) begin
      btb_bank0_rd_data_way1_out_128 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_129 <= 22'h0;
    end else if (_T_1769) begin
      btb_bank0_rd_data_way1_out_129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_130 <= 22'h0;
    end else if (_T_1772) begin
      btb_bank0_rd_data_way1_out_130 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_131 <= 22'h0;
    end else if (_T_1775) begin
      btb_bank0_rd_data_way1_out_131 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_132 <= 22'h0;
    end else if (_T_1778) begin
      btb_bank0_rd_data_way1_out_132 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_133 <= 22'h0;
    end else if (_T_1781) begin
      btb_bank0_rd_data_way1_out_133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_134 <= 22'h0;
    end else if (_T_1784) begin
      btb_bank0_rd_data_way1_out_134 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_135 <= 22'h0;
    end else if (_T_1787) begin
      btb_bank0_rd_data_way1_out_135 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_136 <= 22'h0;
    end else if (_T_1790) begin
      btb_bank0_rd_data_way1_out_136 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_137 <= 22'h0;
    end else if (_T_1793) begin
      btb_bank0_rd_data_way1_out_137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_138 <= 22'h0;
    end else if (_T_1796) begin
      btb_bank0_rd_data_way1_out_138 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_139 <= 22'h0;
    end else if (_T_1799) begin
      btb_bank0_rd_data_way1_out_139 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_140 <= 22'h0;
    end else if (_T_1802) begin
      btb_bank0_rd_data_way1_out_140 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_141 <= 22'h0;
    end else if (_T_1805) begin
      btb_bank0_rd_data_way1_out_141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_142 <= 22'h0;
    end else if (_T_1808) begin
      btb_bank0_rd_data_way1_out_142 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_143 <= 22'h0;
    end else if (_T_1811) begin
      btb_bank0_rd_data_way1_out_143 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_144 <= 22'h0;
    end else if (_T_1814) begin
      btb_bank0_rd_data_way1_out_144 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_145 <= 22'h0;
    end else if (_T_1817) begin
      btb_bank0_rd_data_way1_out_145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_146 <= 22'h0;
    end else if (_T_1820) begin
      btb_bank0_rd_data_way1_out_146 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_147 <= 22'h0;
    end else if (_T_1823) begin
      btb_bank0_rd_data_way1_out_147 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_148 <= 22'h0;
    end else if (_T_1826) begin
      btb_bank0_rd_data_way1_out_148 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_149 <= 22'h0;
    end else if (_T_1829) begin
      btb_bank0_rd_data_way1_out_149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_150 <= 22'h0;
    end else if (_T_1832) begin
      btb_bank0_rd_data_way1_out_150 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_151 <= 22'h0;
    end else if (_T_1835) begin
      btb_bank0_rd_data_way1_out_151 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_152 <= 22'h0;
    end else if (_T_1838) begin
      btb_bank0_rd_data_way1_out_152 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_153 <= 22'h0;
    end else if (_T_1841) begin
      btb_bank0_rd_data_way1_out_153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_154 <= 22'h0;
    end else if (_T_1844) begin
      btb_bank0_rd_data_way1_out_154 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_155 <= 22'h0;
    end else if (_T_1847) begin
      btb_bank0_rd_data_way1_out_155 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_156 <= 22'h0;
    end else if (_T_1850) begin
      btb_bank0_rd_data_way1_out_156 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_157 <= 22'h0;
    end else if (_T_1853) begin
      btb_bank0_rd_data_way1_out_157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_158 <= 22'h0;
    end else if (_T_1856) begin
      btb_bank0_rd_data_way1_out_158 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_159 <= 22'h0;
    end else if (_T_1859) begin
      btb_bank0_rd_data_way1_out_159 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_160 <= 22'h0;
    end else if (_T_1862) begin
      btb_bank0_rd_data_way1_out_160 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_161 <= 22'h0;
    end else if (_T_1865) begin
      btb_bank0_rd_data_way1_out_161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_162 <= 22'h0;
    end else if (_T_1868) begin
      btb_bank0_rd_data_way1_out_162 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_163 <= 22'h0;
    end else if (_T_1871) begin
      btb_bank0_rd_data_way1_out_163 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_164 <= 22'h0;
    end else if (_T_1874) begin
      btb_bank0_rd_data_way1_out_164 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_165 <= 22'h0;
    end else if (_T_1877) begin
      btb_bank0_rd_data_way1_out_165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_166 <= 22'h0;
    end else if (_T_1880) begin
      btb_bank0_rd_data_way1_out_166 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_167 <= 22'h0;
    end else if (_T_1883) begin
      btb_bank0_rd_data_way1_out_167 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_168 <= 22'h0;
    end else if (_T_1886) begin
      btb_bank0_rd_data_way1_out_168 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_169 <= 22'h0;
    end else if (_T_1889) begin
      btb_bank0_rd_data_way1_out_169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_170 <= 22'h0;
    end else if (_T_1892) begin
      btb_bank0_rd_data_way1_out_170 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_171 <= 22'h0;
    end else if (_T_1895) begin
      btb_bank0_rd_data_way1_out_171 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_172 <= 22'h0;
    end else if (_T_1898) begin
      btb_bank0_rd_data_way1_out_172 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_173 <= 22'h0;
    end else if (_T_1901) begin
      btb_bank0_rd_data_way1_out_173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_174 <= 22'h0;
    end else if (_T_1904) begin
      btb_bank0_rd_data_way1_out_174 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_175 <= 22'h0;
    end else if (_T_1907) begin
      btb_bank0_rd_data_way1_out_175 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_176 <= 22'h0;
    end else if (_T_1910) begin
      btb_bank0_rd_data_way1_out_176 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_177 <= 22'h0;
    end else if (_T_1913) begin
      btb_bank0_rd_data_way1_out_177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_178 <= 22'h0;
    end else if (_T_1916) begin
      btb_bank0_rd_data_way1_out_178 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_179 <= 22'h0;
    end else if (_T_1919) begin
      btb_bank0_rd_data_way1_out_179 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_180 <= 22'h0;
    end else if (_T_1922) begin
      btb_bank0_rd_data_way1_out_180 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_181 <= 22'h0;
    end else if (_T_1925) begin
      btb_bank0_rd_data_way1_out_181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_182 <= 22'h0;
    end else if (_T_1928) begin
      btb_bank0_rd_data_way1_out_182 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_183 <= 22'h0;
    end else if (_T_1931) begin
      btb_bank0_rd_data_way1_out_183 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_184 <= 22'h0;
    end else if (_T_1934) begin
      btb_bank0_rd_data_way1_out_184 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_185 <= 22'h0;
    end else if (_T_1937) begin
      btb_bank0_rd_data_way1_out_185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_186 <= 22'h0;
    end else if (_T_1940) begin
      btb_bank0_rd_data_way1_out_186 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_187 <= 22'h0;
    end else if (_T_1943) begin
      btb_bank0_rd_data_way1_out_187 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_188 <= 22'h0;
    end else if (_T_1946) begin
      btb_bank0_rd_data_way1_out_188 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_189 <= 22'h0;
    end else if (_T_1949) begin
      btb_bank0_rd_data_way1_out_189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_190 <= 22'h0;
    end else if (_T_1952) begin
      btb_bank0_rd_data_way1_out_190 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_191 <= 22'h0;
    end else if (_T_1955) begin
      btb_bank0_rd_data_way1_out_191 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_192 <= 22'h0;
    end else if (_T_1958) begin
      btb_bank0_rd_data_way1_out_192 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_193 <= 22'h0;
    end else if (_T_1961) begin
      btb_bank0_rd_data_way1_out_193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_194 <= 22'h0;
    end else if (_T_1964) begin
      btb_bank0_rd_data_way1_out_194 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_195 <= 22'h0;
    end else if (_T_1967) begin
      btb_bank0_rd_data_way1_out_195 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_196 <= 22'h0;
    end else if (_T_1970) begin
      btb_bank0_rd_data_way1_out_196 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_197 <= 22'h0;
    end else if (_T_1973) begin
      btb_bank0_rd_data_way1_out_197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_198 <= 22'h0;
    end else if (_T_1976) begin
      btb_bank0_rd_data_way1_out_198 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_199 <= 22'h0;
    end else if (_T_1979) begin
      btb_bank0_rd_data_way1_out_199 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_200 <= 22'h0;
    end else if (_T_1982) begin
      btb_bank0_rd_data_way1_out_200 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_201 <= 22'h0;
    end else if (_T_1985) begin
      btb_bank0_rd_data_way1_out_201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_202 <= 22'h0;
    end else if (_T_1988) begin
      btb_bank0_rd_data_way1_out_202 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_203 <= 22'h0;
    end else if (_T_1991) begin
      btb_bank0_rd_data_way1_out_203 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_204 <= 22'h0;
    end else if (_T_1994) begin
      btb_bank0_rd_data_way1_out_204 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_205 <= 22'h0;
    end else if (_T_1997) begin
      btb_bank0_rd_data_way1_out_205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_206 <= 22'h0;
    end else if (_T_2000) begin
      btb_bank0_rd_data_way1_out_206 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_207 <= 22'h0;
    end else if (_T_2003) begin
      btb_bank0_rd_data_way1_out_207 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_208 <= 22'h0;
    end else if (_T_2006) begin
      btb_bank0_rd_data_way1_out_208 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_209 <= 22'h0;
    end else if (_T_2009) begin
      btb_bank0_rd_data_way1_out_209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_210 <= 22'h0;
    end else if (_T_2012) begin
      btb_bank0_rd_data_way1_out_210 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_211 <= 22'h0;
    end else if (_T_2015) begin
      btb_bank0_rd_data_way1_out_211 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_212 <= 22'h0;
    end else if (_T_2018) begin
      btb_bank0_rd_data_way1_out_212 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_213 <= 22'h0;
    end else if (_T_2021) begin
      btb_bank0_rd_data_way1_out_213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_214 <= 22'h0;
    end else if (_T_2024) begin
      btb_bank0_rd_data_way1_out_214 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_215 <= 22'h0;
    end else if (_T_2027) begin
      btb_bank0_rd_data_way1_out_215 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_216 <= 22'h0;
    end else if (_T_2030) begin
      btb_bank0_rd_data_way1_out_216 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_217 <= 22'h0;
    end else if (_T_2033) begin
      btb_bank0_rd_data_way1_out_217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_218 <= 22'h0;
    end else if (_T_2036) begin
      btb_bank0_rd_data_way1_out_218 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_219 <= 22'h0;
    end else if (_T_2039) begin
      btb_bank0_rd_data_way1_out_219 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_220 <= 22'h0;
    end else if (_T_2042) begin
      btb_bank0_rd_data_way1_out_220 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_221 <= 22'h0;
    end else if (_T_2045) begin
      btb_bank0_rd_data_way1_out_221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_222 <= 22'h0;
    end else if (_T_2048) begin
      btb_bank0_rd_data_way1_out_222 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_223 <= 22'h0;
    end else if (_T_2051) begin
      btb_bank0_rd_data_way1_out_223 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_224 <= 22'h0;
    end else if (_T_2054) begin
      btb_bank0_rd_data_way1_out_224 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_225 <= 22'h0;
    end else if (_T_2057) begin
      btb_bank0_rd_data_way1_out_225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_226 <= 22'h0;
    end else if (_T_2060) begin
      btb_bank0_rd_data_way1_out_226 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_227 <= 22'h0;
    end else if (_T_2063) begin
      btb_bank0_rd_data_way1_out_227 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_228 <= 22'h0;
    end else if (_T_2066) begin
      btb_bank0_rd_data_way1_out_228 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_229 <= 22'h0;
    end else if (_T_2069) begin
      btb_bank0_rd_data_way1_out_229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_230 <= 22'h0;
    end else if (_T_2072) begin
      btb_bank0_rd_data_way1_out_230 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_231 <= 22'h0;
    end else if (_T_2075) begin
      btb_bank0_rd_data_way1_out_231 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_232 <= 22'h0;
    end else if (_T_2078) begin
      btb_bank0_rd_data_way1_out_232 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_233 <= 22'h0;
    end else if (_T_2081) begin
      btb_bank0_rd_data_way1_out_233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_234 <= 22'h0;
    end else if (_T_2084) begin
      btb_bank0_rd_data_way1_out_234 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_235 <= 22'h0;
    end else if (_T_2087) begin
      btb_bank0_rd_data_way1_out_235 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_236 <= 22'h0;
    end else if (_T_2090) begin
      btb_bank0_rd_data_way1_out_236 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_237 <= 22'h0;
    end else if (_T_2093) begin
      btb_bank0_rd_data_way1_out_237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_238 <= 22'h0;
    end else if (_T_2096) begin
      btb_bank0_rd_data_way1_out_238 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_239 <= 22'h0;
    end else if (_T_2099) begin
      btb_bank0_rd_data_way1_out_239 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_240 <= 22'h0;
    end else if (_T_2102) begin
      btb_bank0_rd_data_way1_out_240 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_241 <= 22'h0;
    end else if (_T_2105) begin
      btb_bank0_rd_data_way1_out_241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_242 <= 22'h0;
    end else if (_T_2108) begin
      btb_bank0_rd_data_way1_out_242 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_243 <= 22'h0;
    end else if (_T_2111) begin
      btb_bank0_rd_data_way1_out_243 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_244 <= 22'h0;
    end else if (_T_2114) begin
      btb_bank0_rd_data_way1_out_244 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_245 <= 22'h0;
    end else if (_T_2117) begin
      btb_bank0_rd_data_way1_out_245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_246 <= 22'h0;
    end else if (_T_2120) begin
      btb_bank0_rd_data_way1_out_246 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_247 <= 22'h0;
    end else if (_T_2123) begin
      btb_bank0_rd_data_way1_out_247 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_248 <= 22'h0;
    end else if (_T_2126) begin
      btb_bank0_rd_data_way1_out_248 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_249 <= 22'h0;
    end else if (_T_2129) begin
      btb_bank0_rd_data_way1_out_249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_250 <= 22'h0;
    end else if (_T_2132) begin
      btb_bank0_rd_data_way1_out_250 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_251 <= 22'h0;
    end else if (_T_2135) begin
      btb_bank0_rd_data_way1_out_251 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_252 <= 22'h0;
    end else if (_T_2138) begin
      btb_bank0_rd_data_way1_out_252 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_253 <= 22'h0;
    end else if (_T_2141) begin
      btb_bank0_rd_data_way1_out_253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_254 <= 22'h0;
    end else if (_T_2144) begin
      btb_bank0_rd_data_way1_out_254 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_255 <= 22'h0;
    end else if (_T_2147) begin
      btb_bank0_rd_data_way1_out_255 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      fghr <= 8'h0;
    end else if (_T_349) begin
      fghr <= fghr_ns;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_8908) begin
        bht_bank_rd_data_out_1_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_8917) begin
        bht_bank_rd_data_out_1_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_8926) begin
        bht_bank_rd_data_out_1_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_8935) begin
        bht_bank_rd_data_out_1_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_8944) begin
        bht_bank_rd_data_out_1_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_8953) begin
        bht_bank_rd_data_out_1_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_8962) begin
        bht_bank_rd_data_out_1_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_8971) begin
        bht_bank_rd_data_out_1_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_8980) begin
        bht_bank_rd_data_out_1_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_8989) begin
        bht_bank_rd_data_out_1_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_8998) begin
        bht_bank_rd_data_out_1_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_9007) begin
        bht_bank_rd_data_out_1_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_9016) begin
        bht_bank_rd_data_out_1_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_9025) begin
        bht_bank_rd_data_out_1_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_9034) begin
        bht_bank_rd_data_out_1_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_9043) begin
        bht_bank_rd_data_out_1_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_9052) begin
        bht_bank_rd_data_out_1_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_9061) begin
        bht_bank_rd_data_out_1_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_9070) begin
        bht_bank_rd_data_out_1_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_9079) begin
        bht_bank_rd_data_out_1_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_9088) begin
        bht_bank_rd_data_out_1_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_9097) begin
        bht_bank_rd_data_out_1_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_9106) begin
        bht_bank_rd_data_out_1_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_9115) begin
        bht_bank_rd_data_out_1_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_9124) begin
        bht_bank_rd_data_out_1_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_9133) begin
        bht_bank_rd_data_out_1_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_9142) begin
        bht_bank_rd_data_out_1_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_9151) begin
        bht_bank_rd_data_out_1_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_9160) begin
        bht_bank_rd_data_out_1_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_9169) begin
        bht_bank_rd_data_out_1_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_9178) begin
        bht_bank_rd_data_out_1_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_9187) begin
        bht_bank_rd_data_out_1_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_9196) begin
        bht_bank_rd_data_out_1_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_9205) begin
        bht_bank_rd_data_out_1_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_9214) begin
        bht_bank_rd_data_out_1_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_9223) begin
        bht_bank_rd_data_out_1_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_9232) begin
        bht_bank_rd_data_out_1_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_9241) begin
        bht_bank_rd_data_out_1_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_9250) begin
        bht_bank_rd_data_out_1_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_9259) begin
        bht_bank_rd_data_out_1_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_9268) begin
        bht_bank_rd_data_out_1_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_9277) begin
        bht_bank_rd_data_out_1_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_9286) begin
        bht_bank_rd_data_out_1_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_9295) begin
        bht_bank_rd_data_out_1_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_9304) begin
        bht_bank_rd_data_out_1_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_9313) begin
        bht_bank_rd_data_out_1_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_9322) begin
        bht_bank_rd_data_out_1_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_9331) begin
        bht_bank_rd_data_out_1_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_9340) begin
        bht_bank_rd_data_out_1_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_9349) begin
        bht_bank_rd_data_out_1_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_9358) begin
        bht_bank_rd_data_out_1_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_9367) begin
        bht_bank_rd_data_out_1_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_9376) begin
        bht_bank_rd_data_out_1_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_9385) begin
        bht_bank_rd_data_out_1_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9394) begin
        bht_bank_rd_data_out_1_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9403) begin
        bht_bank_rd_data_out_1_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9412) begin
        bht_bank_rd_data_out_1_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9421) begin
        bht_bank_rd_data_out_1_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9430) begin
        bht_bank_rd_data_out_1_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9439) begin
        bht_bank_rd_data_out_1_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9448) begin
        bht_bank_rd_data_out_1_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9457) begin
        bht_bank_rd_data_out_1_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_9466) begin
        bht_bank_rd_data_out_1_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_9475) begin
        bht_bank_rd_data_out_1_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_9484) begin
        bht_bank_rd_data_out_1_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_9493) begin
        bht_bank_rd_data_out_1_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_9502) begin
        bht_bank_rd_data_out_1_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_9511) begin
        bht_bank_rd_data_out_1_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_9520) begin
        bht_bank_rd_data_out_1_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_9529) begin
        bht_bank_rd_data_out_1_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_9538) begin
        bht_bank_rd_data_out_1_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_9547) begin
        bht_bank_rd_data_out_1_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_9556) begin
        bht_bank_rd_data_out_1_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_9565) begin
        bht_bank_rd_data_out_1_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_9574) begin
        bht_bank_rd_data_out_1_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_9583) begin
        bht_bank_rd_data_out_1_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_9592) begin
        bht_bank_rd_data_out_1_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_9601) begin
        bht_bank_rd_data_out_1_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_9610) begin
        bht_bank_rd_data_out_1_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_9619) begin
        bht_bank_rd_data_out_1_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_9628) begin
        bht_bank_rd_data_out_1_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_9637) begin
        bht_bank_rd_data_out_1_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_9646) begin
        bht_bank_rd_data_out_1_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_9655) begin
        bht_bank_rd_data_out_1_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_9664) begin
        bht_bank_rd_data_out_1_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_9673) begin
        bht_bank_rd_data_out_1_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_9682) begin
        bht_bank_rd_data_out_1_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_9691) begin
        bht_bank_rd_data_out_1_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_9700) begin
        bht_bank_rd_data_out_1_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_9709) begin
        bht_bank_rd_data_out_1_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_9718) begin
        bht_bank_rd_data_out_1_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_9727) begin
        bht_bank_rd_data_out_1_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_9736) begin
        bht_bank_rd_data_out_1_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_9745) begin
        bht_bank_rd_data_out_1_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_9754) begin
        bht_bank_rd_data_out_1_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_9763) begin
        bht_bank_rd_data_out_1_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_9772) begin
        bht_bank_rd_data_out_1_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_9781) begin
        bht_bank_rd_data_out_1_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_9790) begin
        bht_bank_rd_data_out_1_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_9799) begin
        bht_bank_rd_data_out_1_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_9808) begin
        bht_bank_rd_data_out_1_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_9817) begin
        bht_bank_rd_data_out_1_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_9826) begin
        bht_bank_rd_data_out_1_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_9835) begin
        bht_bank_rd_data_out_1_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_9844) begin
        bht_bank_rd_data_out_1_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_9853) begin
        bht_bank_rd_data_out_1_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_9862) begin
        bht_bank_rd_data_out_1_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_9871) begin
        bht_bank_rd_data_out_1_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_9880) begin
        bht_bank_rd_data_out_1_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_9889) begin
        bht_bank_rd_data_out_1_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_9898) begin
        bht_bank_rd_data_out_1_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_9907) begin
        bht_bank_rd_data_out_1_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_9916) begin
        bht_bank_rd_data_out_1_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_9925) begin
        bht_bank_rd_data_out_1_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_9934) begin
        bht_bank_rd_data_out_1_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_9943) begin
        bht_bank_rd_data_out_1_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_9952) begin
        bht_bank_rd_data_out_1_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_9961) begin
        bht_bank_rd_data_out_1_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_9970) begin
        bht_bank_rd_data_out_1_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_9979) begin
        bht_bank_rd_data_out_1_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_9988) begin
        bht_bank_rd_data_out_1_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_9997) begin
        bht_bank_rd_data_out_1_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_10006) begin
        bht_bank_rd_data_out_1_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_10015) begin
        bht_bank_rd_data_out_1_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_10024) begin
        bht_bank_rd_data_out_1_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_10033) begin
        bht_bank_rd_data_out_1_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_10042) begin
        bht_bank_rd_data_out_1_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_10051) begin
        bht_bank_rd_data_out_1_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_10060) begin
        bht_bank_rd_data_out_1_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_10069) begin
        bht_bank_rd_data_out_1_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_10078) begin
        bht_bank_rd_data_out_1_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_10087) begin
        bht_bank_rd_data_out_1_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_10096) begin
        bht_bank_rd_data_out_1_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_10105) begin
        bht_bank_rd_data_out_1_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_10114) begin
        bht_bank_rd_data_out_1_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_10123) begin
        bht_bank_rd_data_out_1_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_10132) begin
        bht_bank_rd_data_out_1_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_10141) begin
        bht_bank_rd_data_out_1_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_10150) begin
        bht_bank_rd_data_out_1_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_10159) begin
        bht_bank_rd_data_out_1_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_10168) begin
        bht_bank_rd_data_out_1_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_10177) begin
        bht_bank_rd_data_out_1_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_10186) begin
        bht_bank_rd_data_out_1_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_10195) begin
        bht_bank_rd_data_out_1_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_10204) begin
        bht_bank_rd_data_out_1_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_10213) begin
        bht_bank_rd_data_out_1_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_10222) begin
        bht_bank_rd_data_out_1_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_10231) begin
        bht_bank_rd_data_out_1_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_10240) begin
        bht_bank_rd_data_out_1_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_10249) begin
        bht_bank_rd_data_out_1_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_10258) begin
        bht_bank_rd_data_out_1_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_10267) begin
        bht_bank_rd_data_out_1_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_10276) begin
        bht_bank_rd_data_out_1_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_10285) begin
        bht_bank_rd_data_out_1_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_10294) begin
        bht_bank_rd_data_out_1_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_10303) begin
        bht_bank_rd_data_out_1_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_10312) begin
        bht_bank_rd_data_out_1_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_10321) begin
        bht_bank_rd_data_out_1_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_10330) begin
        bht_bank_rd_data_out_1_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_10339) begin
        bht_bank_rd_data_out_1_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_10348) begin
        bht_bank_rd_data_out_1_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_10357) begin
        bht_bank_rd_data_out_1_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_10366) begin
        bht_bank_rd_data_out_1_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_10375) begin
        bht_bank_rd_data_out_1_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_10384) begin
        bht_bank_rd_data_out_1_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_10393) begin
        bht_bank_rd_data_out_1_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10402) begin
        bht_bank_rd_data_out_1_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10411) begin
        bht_bank_rd_data_out_1_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10420) begin
        bht_bank_rd_data_out_1_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10429) begin
        bht_bank_rd_data_out_1_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10438) begin
        bht_bank_rd_data_out_1_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10447) begin
        bht_bank_rd_data_out_1_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10456) begin
        bht_bank_rd_data_out_1_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_10465) begin
        bht_bank_rd_data_out_1_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_10474) begin
        bht_bank_rd_data_out_1_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_10483) begin
        bht_bank_rd_data_out_1_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_10492) begin
        bht_bank_rd_data_out_1_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_10501) begin
        bht_bank_rd_data_out_1_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_10510) begin
        bht_bank_rd_data_out_1_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_10519) begin
        bht_bank_rd_data_out_1_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_10528) begin
        bht_bank_rd_data_out_1_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_10537) begin
        bht_bank_rd_data_out_1_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_10546) begin
        bht_bank_rd_data_out_1_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_10555) begin
        bht_bank_rd_data_out_1_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_10564) begin
        bht_bank_rd_data_out_1_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_10573) begin
        bht_bank_rd_data_out_1_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_10582) begin
        bht_bank_rd_data_out_1_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_10591) begin
        bht_bank_rd_data_out_1_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_10600) begin
        bht_bank_rd_data_out_1_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_10609) begin
        bht_bank_rd_data_out_1_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_10618) begin
        bht_bank_rd_data_out_1_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_10627) begin
        bht_bank_rd_data_out_1_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_10636) begin
        bht_bank_rd_data_out_1_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_10645) begin
        bht_bank_rd_data_out_1_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_10654) begin
        bht_bank_rd_data_out_1_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_10663) begin
        bht_bank_rd_data_out_1_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_10672) begin
        bht_bank_rd_data_out_1_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_10681) begin
        bht_bank_rd_data_out_1_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_10690) begin
        bht_bank_rd_data_out_1_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_10699) begin
        bht_bank_rd_data_out_1_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_10708) begin
        bht_bank_rd_data_out_1_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_10717) begin
        bht_bank_rd_data_out_1_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_10726) begin
        bht_bank_rd_data_out_1_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_10735) begin
        bht_bank_rd_data_out_1_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_10744) begin
        bht_bank_rd_data_out_1_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_10753) begin
        bht_bank_rd_data_out_1_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_10762) begin
        bht_bank_rd_data_out_1_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_10771) begin
        bht_bank_rd_data_out_1_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_10780) begin
        bht_bank_rd_data_out_1_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_10789) begin
        bht_bank_rd_data_out_1_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_10798) begin
        bht_bank_rd_data_out_1_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_10807) begin
        bht_bank_rd_data_out_1_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_10816) begin
        bht_bank_rd_data_out_1_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_10825) begin
        bht_bank_rd_data_out_1_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_10834) begin
        bht_bank_rd_data_out_1_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_10843) begin
        bht_bank_rd_data_out_1_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_10852) begin
        bht_bank_rd_data_out_1_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_10861) begin
        bht_bank_rd_data_out_1_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_10870) begin
        bht_bank_rd_data_out_1_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_10879) begin
        bht_bank_rd_data_out_1_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_10888) begin
        bht_bank_rd_data_out_1_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_10897) begin
        bht_bank_rd_data_out_1_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_10906) begin
        bht_bank_rd_data_out_1_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_10915) begin
        bht_bank_rd_data_out_1_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_10924) begin
        bht_bank_rd_data_out_1_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_10933) begin
        bht_bank_rd_data_out_1_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_10942) begin
        bht_bank_rd_data_out_1_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_10951) begin
        bht_bank_rd_data_out_1_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_10960) begin
        bht_bank_rd_data_out_1_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_10969) begin
        bht_bank_rd_data_out_1_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_10978) begin
        bht_bank_rd_data_out_1_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_10987) begin
        bht_bank_rd_data_out_1_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_10996) begin
        bht_bank_rd_data_out_1_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_11005) begin
        bht_bank_rd_data_out_1_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_11014) begin
        bht_bank_rd_data_out_1_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_11023) begin
        bht_bank_rd_data_out_1_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_11032) begin
        bht_bank_rd_data_out_1_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_11041) begin
        bht_bank_rd_data_out_1_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_11050) begin
        bht_bank_rd_data_out_1_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_11059) begin
        bht_bank_rd_data_out_1_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_11068) begin
        bht_bank_rd_data_out_1_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_11077) begin
        bht_bank_rd_data_out_1_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_11086) begin
        bht_bank_rd_data_out_1_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_11095) begin
        bht_bank_rd_data_out_1_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_11104) begin
        bht_bank_rd_data_out_1_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_11113) begin
        bht_bank_rd_data_out_1_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_11122) begin
        bht_bank_rd_data_out_1_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_11131) begin
        bht_bank_rd_data_out_1_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_11140) begin
        bht_bank_rd_data_out_1_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_11149) begin
        bht_bank_rd_data_out_1_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_11158) begin
        bht_bank_rd_data_out_1_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_11167) begin
        bht_bank_rd_data_out_1_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_11176) begin
        bht_bank_rd_data_out_1_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_11185) begin
        bht_bank_rd_data_out_1_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_11194) begin
        bht_bank_rd_data_out_1_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_11203) begin
        bht_bank_rd_data_out_1_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_6604) begin
        bht_bank_rd_data_out_0_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_6613) begin
        bht_bank_rd_data_out_0_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_6622) begin
        bht_bank_rd_data_out_0_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_6631) begin
        bht_bank_rd_data_out_0_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_6640) begin
        bht_bank_rd_data_out_0_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_6649) begin
        bht_bank_rd_data_out_0_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_6658) begin
        bht_bank_rd_data_out_0_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_6667) begin
        bht_bank_rd_data_out_0_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_6676) begin
        bht_bank_rd_data_out_0_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_6685) begin
        bht_bank_rd_data_out_0_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_6694) begin
        bht_bank_rd_data_out_0_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_6703) begin
        bht_bank_rd_data_out_0_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_6712) begin
        bht_bank_rd_data_out_0_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_6721) begin
        bht_bank_rd_data_out_0_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_6730) begin
        bht_bank_rd_data_out_0_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_6739) begin
        bht_bank_rd_data_out_0_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_6748) begin
        bht_bank_rd_data_out_0_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_6757) begin
        bht_bank_rd_data_out_0_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_6766) begin
        bht_bank_rd_data_out_0_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_6775) begin
        bht_bank_rd_data_out_0_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_6784) begin
        bht_bank_rd_data_out_0_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_6793) begin
        bht_bank_rd_data_out_0_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_6802) begin
        bht_bank_rd_data_out_0_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_6811) begin
        bht_bank_rd_data_out_0_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_6820) begin
        bht_bank_rd_data_out_0_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_6829) begin
        bht_bank_rd_data_out_0_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_6838) begin
        bht_bank_rd_data_out_0_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_6847) begin
        bht_bank_rd_data_out_0_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_6856) begin
        bht_bank_rd_data_out_0_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_6865) begin
        bht_bank_rd_data_out_0_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_6874) begin
        bht_bank_rd_data_out_0_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_6883) begin
        bht_bank_rd_data_out_0_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_6892) begin
        bht_bank_rd_data_out_0_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_6901) begin
        bht_bank_rd_data_out_0_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_6910) begin
        bht_bank_rd_data_out_0_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_6919) begin
        bht_bank_rd_data_out_0_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_6928) begin
        bht_bank_rd_data_out_0_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_6937) begin
        bht_bank_rd_data_out_0_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_6946) begin
        bht_bank_rd_data_out_0_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_6955) begin
        bht_bank_rd_data_out_0_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_6964) begin
        bht_bank_rd_data_out_0_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_6973) begin
        bht_bank_rd_data_out_0_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_6982) begin
        bht_bank_rd_data_out_0_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_6991) begin
        bht_bank_rd_data_out_0_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_7000) begin
        bht_bank_rd_data_out_0_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_7009) begin
        bht_bank_rd_data_out_0_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_7018) begin
        bht_bank_rd_data_out_0_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_7027) begin
        bht_bank_rd_data_out_0_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_7036) begin
        bht_bank_rd_data_out_0_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_7045) begin
        bht_bank_rd_data_out_0_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_7054) begin
        bht_bank_rd_data_out_0_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_7063) begin
        bht_bank_rd_data_out_0_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_7072) begin
        bht_bank_rd_data_out_0_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_7081) begin
        bht_bank_rd_data_out_0_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_7090) begin
        bht_bank_rd_data_out_0_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_7099) begin
        bht_bank_rd_data_out_0_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_7108) begin
        bht_bank_rd_data_out_0_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_7117) begin
        bht_bank_rd_data_out_0_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_7126) begin
        bht_bank_rd_data_out_0_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_7135) begin
        bht_bank_rd_data_out_0_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_7144) begin
        bht_bank_rd_data_out_0_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_7153) begin
        bht_bank_rd_data_out_0_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_7162) begin
        bht_bank_rd_data_out_0_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_7171) begin
        bht_bank_rd_data_out_0_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_7180) begin
        bht_bank_rd_data_out_0_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_7189) begin
        bht_bank_rd_data_out_0_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_7198) begin
        bht_bank_rd_data_out_0_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_7207) begin
        bht_bank_rd_data_out_0_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_7216) begin
        bht_bank_rd_data_out_0_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_7225) begin
        bht_bank_rd_data_out_0_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_7234) begin
        bht_bank_rd_data_out_0_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_7243) begin
        bht_bank_rd_data_out_0_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_7252) begin
        bht_bank_rd_data_out_0_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_7261) begin
        bht_bank_rd_data_out_0_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_7270) begin
        bht_bank_rd_data_out_0_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_7279) begin
        bht_bank_rd_data_out_0_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_7288) begin
        bht_bank_rd_data_out_0_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_7297) begin
        bht_bank_rd_data_out_0_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_7306) begin
        bht_bank_rd_data_out_0_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_7315) begin
        bht_bank_rd_data_out_0_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_7324) begin
        bht_bank_rd_data_out_0_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_7333) begin
        bht_bank_rd_data_out_0_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_7342) begin
        bht_bank_rd_data_out_0_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_7351) begin
        bht_bank_rd_data_out_0_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_7360) begin
        bht_bank_rd_data_out_0_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_7369) begin
        bht_bank_rd_data_out_0_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_7378) begin
        bht_bank_rd_data_out_0_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_7387) begin
        bht_bank_rd_data_out_0_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7396) begin
        bht_bank_rd_data_out_0_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7405) begin
        bht_bank_rd_data_out_0_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7414) begin
        bht_bank_rd_data_out_0_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7423) begin
        bht_bank_rd_data_out_0_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7432) begin
        bht_bank_rd_data_out_0_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7441) begin
        bht_bank_rd_data_out_0_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7450) begin
        bht_bank_rd_data_out_0_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_7459) begin
        bht_bank_rd_data_out_0_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_7468) begin
        bht_bank_rd_data_out_0_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_7477) begin
        bht_bank_rd_data_out_0_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_7486) begin
        bht_bank_rd_data_out_0_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_7495) begin
        bht_bank_rd_data_out_0_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_7504) begin
        bht_bank_rd_data_out_0_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_7513) begin
        bht_bank_rd_data_out_0_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_7522) begin
        bht_bank_rd_data_out_0_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_7531) begin
        bht_bank_rd_data_out_0_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_7540) begin
        bht_bank_rd_data_out_0_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_7549) begin
        bht_bank_rd_data_out_0_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_7558) begin
        bht_bank_rd_data_out_0_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_7567) begin
        bht_bank_rd_data_out_0_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_7576) begin
        bht_bank_rd_data_out_0_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_7585) begin
        bht_bank_rd_data_out_0_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_7594) begin
        bht_bank_rd_data_out_0_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_7603) begin
        bht_bank_rd_data_out_0_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_7612) begin
        bht_bank_rd_data_out_0_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_7621) begin
        bht_bank_rd_data_out_0_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_7630) begin
        bht_bank_rd_data_out_0_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_7639) begin
        bht_bank_rd_data_out_0_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_7648) begin
        bht_bank_rd_data_out_0_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_7657) begin
        bht_bank_rd_data_out_0_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_7666) begin
        bht_bank_rd_data_out_0_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_7675) begin
        bht_bank_rd_data_out_0_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_7684) begin
        bht_bank_rd_data_out_0_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_7693) begin
        bht_bank_rd_data_out_0_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_7702) begin
        bht_bank_rd_data_out_0_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_7711) begin
        bht_bank_rd_data_out_0_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_7720) begin
        bht_bank_rd_data_out_0_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_7729) begin
        bht_bank_rd_data_out_0_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_7738) begin
        bht_bank_rd_data_out_0_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_7747) begin
        bht_bank_rd_data_out_0_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_7756) begin
        bht_bank_rd_data_out_0_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_7765) begin
        bht_bank_rd_data_out_0_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_7774) begin
        bht_bank_rd_data_out_0_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_7783) begin
        bht_bank_rd_data_out_0_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_7792) begin
        bht_bank_rd_data_out_0_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_7801) begin
        bht_bank_rd_data_out_0_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_7810) begin
        bht_bank_rd_data_out_0_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_7819) begin
        bht_bank_rd_data_out_0_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_7828) begin
        bht_bank_rd_data_out_0_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_7837) begin
        bht_bank_rd_data_out_0_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_7846) begin
        bht_bank_rd_data_out_0_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_7855) begin
        bht_bank_rd_data_out_0_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_7864) begin
        bht_bank_rd_data_out_0_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_7873) begin
        bht_bank_rd_data_out_0_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_7882) begin
        bht_bank_rd_data_out_0_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_7891) begin
        bht_bank_rd_data_out_0_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_7900) begin
        bht_bank_rd_data_out_0_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_7909) begin
        bht_bank_rd_data_out_0_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_7918) begin
        bht_bank_rd_data_out_0_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_7927) begin
        bht_bank_rd_data_out_0_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_7936) begin
        bht_bank_rd_data_out_0_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_7945) begin
        bht_bank_rd_data_out_0_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_7954) begin
        bht_bank_rd_data_out_0_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_7963) begin
        bht_bank_rd_data_out_0_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_7972) begin
        bht_bank_rd_data_out_0_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_7981) begin
        bht_bank_rd_data_out_0_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_7990) begin
        bht_bank_rd_data_out_0_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_7999) begin
        bht_bank_rd_data_out_0_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_8008) begin
        bht_bank_rd_data_out_0_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_8017) begin
        bht_bank_rd_data_out_0_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_8026) begin
        bht_bank_rd_data_out_0_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_8035) begin
        bht_bank_rd_data_out_0_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_8044) begin
        bht_bank_rd_data_out_0_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_8053) begin
        bht_bank_rd_data_out_0_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_8062) begin
        bht_bank_rd_data_out_0_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_8071) begin
        bht_bank_rd_data_out_0_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_8080) begin
        bht_bank_rd_data_out_0_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_8089) begin
        bht_bank_rd_data_out_0_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_8098) begin
        bht_bank_rd_data_out_0_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_8107) begin
        bht_bank_rd_data_out_0_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_8116) begin
        bht_bank_rd_data_out_0_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_8125) begin
        bht_bank_rd_data_out_0_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_8134) begin
        bht_bank_rd_data_out_0_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_8143) begin
        bht_bank_rd_data_out_0_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_8152) begin
        bht_bank_rd_data_out_0_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_8161) begin
        bht_bank_rd_data_out_0_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_8170) begin
        bht_bank_rd_data_out_0_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_8179) begin
        bht_bank_rd_data_out_0_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_8188) begin
        bht_bank_rd_data_out_0_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_8197) begin
        bht_bank_rd_data_out_0_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_8206) begin
        bht_bank_rd_data_out_0_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_8215) begin
        bht_bank_rd_data_out_0_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_8224) begin
        bht_bank_rd_data_out_0_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_8233) begin
        bht_bank_rd_data_out_0_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_8242) begin
        bht_bank_rd_data_out_0_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_8251) begin
        bht_bank_rd_data_out_0_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_8260) begin
        bht_bank_rd_data_out_0_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_8269) begin
        bht_bank_rd_data_out_0_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_8278) begin
        bht_bank_rd_data_out_0_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_8287) begin
        bht_bank_rd_data_out_0_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_8296) begin
        bht_bank_rd_data_out_0_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_8305) begin
        bht_bank_rd_data_out_0_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_8314) begin
        bht_bank_rd_data_out_0_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_8323) begin
        bht_bank_rd_data_out_0_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_8332) begin
        bht_bank_rd_data_out_0_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_8341) begin
        bht_bank_rd_data_out_0_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_8350) begin
        bht_bank_rd_data_out_0_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_8359) begin
        bht_bank_rd_data_out_0_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_8368) begin
        bht_bank_rd_data_out_0_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_8377) begin
        bht_bank_rd_data_out_0_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_8386) begin
        bht_bank_rd_data_out_0_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8395) begin
        bht_bank_rd_data_out_0_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8404) begin
        bht_bank_rd_data_out_0_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8413) begin
        bht_bank_rd_data_out_0_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8422) begin
        bht_bank_rd_data_out_0_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8431) begin
        bht_bank_rd_data_out_0_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8440) begin
        bht_bank_rd_data_out_0_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8449) begin
        bht_bank_rd_data_out_0_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8458) begin
        bht_bank_rd_data_out_0_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_8467) begin
        bht_bank_rd_data_out_0_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_8476) begin
        bht_bank_rd_data_out_0_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_8485) begin
        bht_bank_rd_data_out_0_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_8494) begin
        bht_bank_rd_data_out_0_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_8503) begin
        bht_bank_rd_data_out_0_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_8512) begin
        bht_bank_rd_data_out_0_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_8521) begin
        bht_bank_rd_data_out_0_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_8530) begin
        bht_bank_rd_data_out_0_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_8539) begin
        bht_bank_rd_data_out_0_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_8548) begin
        bht_bank_rd_data_out_0_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_8557) begin
        bht_bank_rd_data_out_0_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_8566) begin
        bht_bank_rd_data_out_0_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_8575) begin
        bht_bank_rd_data_out_0_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_8584) begin
        bht_bank_rd_data_out_0_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_8593) begin
        bht_bank_rd_data_out_0_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_8602) begin
        bht_bank_rd_data_out_0_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_8611) begin
        bht_bank_rd_data_out_0_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_8620) begin
        bht_bank_rd_data_out_0_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_8629) begin
        bht_bank_rd_data_out_0_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_8638) begin
        bht_bank_rd_data_out_0_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_8647) begin
        bht_bank_rd_data_out_0_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_8656) begin
        bht_bank_rd_data_out_0_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_8665) begin
        bht_bank_rd_data_out_0_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_8674) begin
        bht_bank_rd_data_out_0_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_8683) begin
        bht_bank_rd_data_out_0_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_8692) begin
        bht_bank_rd_data_out_0_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_8701) begin
        bht_bank_rd_data_out_0_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_8710) begin
        bht_bank_rd_data_out_0_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_8719) begin
        bht_bank_rd_data_out_0_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_8728) begin
        bht_bank_rd_data_out_0_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_8737) begin
        bht_bank_rd_data_out_0_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_8746) begin
        bht_bank_rd_data_out_0_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_8755) begin
        bht_bank_rd_data_out_0_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_8764) begin
        bht_bank_rd_data_out_0_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_8773) begin
        bht_bank_rd_data_out_0_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_8782) begin
        bht_bank_rd_data_out_0_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_8791) begin
        bht_bank_rd_data_out_0_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_8800) begin
        bht_bank_rd_data_out_0_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_8809) begin
        bht_bank_rd_data_out_0_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_8818) begin
        bht_bank_rd_data_out_0_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_8827) begin
        bht_bank_rd_data_out_0_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_8836) begin
        bht_bank_rd_data_out_0_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_8845) begin
        bht_bank_rd_data_out_0_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_8854) begin
        bht_bank_rd_data_out_0_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_8863) begin
        bht_bank_rd_data_out_0_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_8872) begin
        bht_bank_rd_data_out_0_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_8881) begin
        bht_bank_rd_data_out_0_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_8890) begin
        bht_bank_rd_data_out_0_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_8899) begin
        bht_bank_rd_data_out_0_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else if (_T_341) begin
      exu_mp_way_f <= io_exu_bp_exu_mp_pkt_bits_way;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else if (_T_208) begin
      btb_lru_b0_f <= btb_lru_b0_ns;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else if (_T_345) begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_fetch_adder_prior <= 30'h0;
    end else if (_T_385) begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f[30:1];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else if (rsenable_0) begin
      rets_out_0 <= rets_in_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_1 <= rets_in_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_2 <= rets_in_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_3 <= rets_in_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_4 <= rets_in_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_5 <= rets_in_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_6 <= rets_in_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else if (rs_push) begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
