module el2_ifu_compress_ctl(
  input         clock,
  input         reset,
  input  [15:0] io_in,
  output [31:0] io_out
);
  wire  _T_4 = ~io_in[14]; // @[el2_ifu_compress_ctl.scala 18:34]
  wire  _T_5 = io_in[15] & _T_4; // @[el2_ifu_compress_ctl.scala 18:32]
  wire  _T_7 = ~io_in[13]; // @[el2_ifu_compress_ctl.scala 18:47]
  wire  _T_8 = _T_5 & _T_7; // @[el2_ifu_compress_ctl.scala 18:45]
  wire  _T_10 = _T_8 & io_in[10]; // @[el2_ifu_compress_ctl.scala 18:58]
  wire  _T_12 = ~io_in[6]; // @[el2_ifu_compress_ctl.scala 18:70]
  wire  _T_13 = _T_10 & _T_12; // @[el2_ifu_compress_ctl.scala 18:68]
  wire  _T_15 = ~io_in[5]; // @[el2_ifu_compress_ctl.scala 18:82]
  wire  _T_16 = _T_13 & _T_15; // @[el2_ifu_compress_ctl.scala 18:80]
  wire  _T_18 = _T_16 & io_in[0]; // @[el2_ifu_compress_ctl.scala 18:92]
  wire  _T_22 = io_in[14] & _T_4; // @[el2_ifu_compress_ctl.scala 19:27]
  wire  _T_25 = _T_22 & _T_7; // @[el2_ifu_compress_ctl.scala 19:40]
  wire  _T_27 = ~io_in[11]; // @[el2_ifu_compress_ctl.scala 19:55]
  wire  _T_28 = _T_25 & _T_27; // @[el2_ifu_compress_ctl.scala 19:53]
  wire  _T_30 = _T_28 & io_in[10]; // @[el2_ifu_compress_ctl.scala 19:66]
  wire  _T_32 = _T_30 & io_in[0]; // @[el2_ifu_compress_ctl.scala 19:76]
  wire  _T_33 = _T_18 | _T_32; // @[el2_ifu_compress_ctl.scala 19:15]
  wire  _T_38 = _T_4 & io_in[12]; // @[el2_ifu_compress_ctl.scala 20:25]
  wire  _T_41 = _T_38 & _T_27; // @[el2_ifu_compress_ctl.scala 20:35]
  wire  _T_43 = ~io_in[10]; // @[el2_ifu_compress_ctl.scala 20:50]
  wire  _T_44 = _T_41 & _T_43; // @[el2_ifu_compress_ctl.scala 20:48]
  wire  _T_46 = ~io_in[9]; // @[el2_ifu_compress_ctl.scala 20:63]
  wire  _T_47 = _T_44 & _T_46; // @[el2_ifu_compress_ctl.scala 20:61]
  wire  _T_49 = ~io_in[8]; // @[el2_ifu_compress_ctl.scala 20:75]
  wire  _T_50 = _T_47 & _T_49; // @[el2_ifu_compress_ctl.scala 20:73]
  wire  _T_52 = ~io_in[7]; // @[el2_ifu_compress_ctl.scala 20:87]
  wire  _T_53 = _T_50 & _T_52; // @[el2_ifu_compress_ctl.scala 20:85]
  wire  _T_56 = _T_53 & _T_12; // @[el2_ifu_compress_ctl.scala 20:97]
  wire  _T_59 = _T_56 & _T_15; // @[el2_ifu_compress_ctl.scala 20:109]
  wire  _T_61 = ~io_in[4]; // @[el2_ifu_compress_ctl.scala 21:16]
  wire  _T_62 = _T_59 & _T_61; // @[el2_ifu_compress_ctl.scala 20:121]
  wire  _T_64 = ~io_in[3]; // @[el2_ifu_compress_ctl.scala 21:28]
  wire  _T_65 = _T_62 & _T_64; // @[el2_ifu_compress_ctl.scala 21:26]
  wire  _T_67 = ~io_in[2]; // @[el2_ifu_compress_ctl.scala 21:40]
  wire  _T_68 = _T_65 & _T_67; // @[el2_ifu_compress_ctl.scala 21:38]
  wire  _T_70 = _T_68 & io_in[1]; // @[el2_ifu_compress_ctl.scala 21:50]
  wire  _T_81 = _T_8 & _T_27; // @[el2_ifu_compress_ctl.scala 22:50]
  wire  _T_83 = _T_81 & io_in[0]; // @[el2_ifu_compress_ctl.scala 22:63]
  wire  _T_93 = _T_8 & _T_43; // @[el2_ifu_compress_ctl.scala 23:51]
  wire  _T_95 = _T_93 & io_in[0]; // @[el2_ifu_compress_ctl.scala 23:64]
  wire  _T_96 = _T_83 | _T_95; // @[el2_ifu_compress_ctl.scala 23:15]
  wire  _T_105 = _T_8 & io_in[6]; // @[el2_ifu_compress_ctl.scala 24:51]
  wire  _T_107 = _T_105 & io_in[0]; // @[el2_ifu_compress_ctl.scala 24:60]
  wire  _T_108 = _T_96 | _T_107; // @[el2_ifu_compress_ctl.scala 24:15]
  wire  _T_117 = _T_8 & io_in[5]; // @[el2_ifu_compress_ctl.scala 25:51]
  wire  _T_119 = _T_117 & io_in[0]; // @[el2_ifu_compress_ctl.scala 25:60]
  wire  _T_120 = _T_108 | _T_119; // @[el2_ifu_compress_ctl.scala 25:15]
  wire  _T_131 = _T_105 & io_in[5]; // @[el2_ifu_compress_ctl.scala 26:59]
  wire  _T_133 = _T_131 & io_in[0]; // @[el2_ifu_compress_ctl.scala 26:68]
  wire  _T_146 = _T_133 | _T_83; // @[el2_ifu_compress_ctl.scala 27:15]
  wire  _T_159 = _T_146 | _T_95; // @[el2_ifu_compress_ctl.scala 28:15]
  wire  _T_161 = ~io_in[15]; // @[el2_ifu_compress_ctl.scala 29:17]
  wire  _T_164 = _T_161 & _T_4; // @[el2_ifu_compress_ctl.scala 29:28]
  wire  _T_166 = _T_164 & io_in[1]; // @[el2_ifu_compress_ctl.scala 29:41]
  wire  _T_167 = _T_159 | _T_166; // @[el2_ifu_compress_ctl.scala 29:15]
  wire  _T_170 = io_in[15] & io_in[14]; // @[el2_ifu_compress_ctl.scala 29:62]
  wire  _T_172 = _T_170 & io_in[13]; // @[el2_ifu_compress_ctl.scala 29:72]
  wire  _T_173 = _T_167 | _T_172; // @[el2_ifu_compress_ctl.scala 29:51]
  wire  _T_234 = _T_5 & _T_12; // @[el2_ifu_compress_ctl.scala 34:37]
  wire  _T_237 = _T_234 & _T_15; // @[el2_ifu_compress_ctl.scala 34:49]
  wire  _T_240 = _T_237 & _T_61; // @[el2_ifu_compress_ctl.scala 34:61]
  wire  _T_243 = _T_240 & _T_64; // @[el2_ifu_compress_ctl.scala 34:73]
  wire  _T_246 = _T_243 & _T_67; // @[el2_ifu_compress_ctl.scala 34:85]
  wire  _T_248 = ~io_in[0]; // @[el2_ifu_compress_ctl.scala 34:99]
  wire  _T_249 = _T_246 & _T_248; // @[el2_ifu_compress_ctl.scala 34:97]
  wire  _T_253 = _T_4 & io_in[13]; // @[el2_ifu_compress_ctl.scala 35:28]
  wire  _T_254 = _T_249 | _T_253; // @[el2_ifu_compress_ctl.scala 35:15]
  wire  _T_259 = _T_170 & io_in[0]; // @[el2_ifu_compress_ctl.scala 35:60]
  wire  _T_260 = _T_254 | _T_259; // @[el2_ifu_compress_ctl.scala 35:39]
  wire  _T_264 = io_in[15] & _T_248; // @[el2_ifu_compress_ctl.scala 35:80]
  wire  _T_267 = io_in[15] & io_in[11]; // @[el2_ifu_compress_ctl.scala 36:25]
  wire  _T_269 = _T_267 & io_in[10]; // @[el2_ifu_compress_ctl.scala 36:35]
  wire  _T_270 = _T_264 | _T_269; // @[el2_ifu_compress_ctl.scala 36:15]
  wire  _T_274 = io_in[13] & _T_49; // @[el2_ifu_compress_ctl.scala 36:57]
  wire  _T_275 = _T_270 | _T_274; // @[el2_ifu_compress_ctl.scala 36:46]
  wire  _T_280 = _T_275 | _T_274; // @[el2_ifu_compress_ctl.scala 37:15]
  wire  _T_283 = io_in[13] & io_in[7]; // @[el2_ifu_compress_ctl.scala 37:47]
  wire  _T_284 = _T_280 | _T_283; // @[el2_ifu_compress_ctl.scala 37:37]
  wire  _T_287 = io_in[13] & io_in[9]; // @[el2_ifu_compress_ctl.scala 37:66]
  wire  _T_288 = _T_284 | _T_287; // @[el2_ifu_compress_ctl.scala 37:56]
  wire  _T_291 = io_in[13] & io_in[10]; // @[el2_ifu_compress_ctl.scala 37:85]
  wire  _T_292 = _T_288 | _T_291; // @[el2_ifu_compress_ctl.scala 37:75]
  wire  _T_295 = io_in[13] & io_in[11]; // @[el2_ifu_compress_ctl.scala 38:25]
  wire  _T_296 = _T_292 | _T_295; // @[el2_ifu_compress_ctl.scala 38:15]
  wire  _T_300 = io_in[13] & _T_4; // @[el2_ifu_compress_ctl.scala 38:45]
  wire  _T_301 = _T_296 | _T_300; // @[el2_ifu_compress_ctl.scala 38:35]
  wire  _T_304 = io_in[14] & io_in[15]; // @[el2_ifu_compress_ctl.scala 38:68]
  wire  _T_305 = _T_301 | _T_304; // @[el2_ifu_compress_ctl.scala 38:58]
  wire  _T_310 = _T_4 & _T_27; // @[el2_ifu_compress_ctl.scala 39:25]
  wire  _T_313 = _T_310 & _T_43; // @[el2_ifu_compress_ctl.scala 39:38]
  wire  _T_316 = _T_313 & _T_46; // @[el2_ifu_compress_ctl.scala 39:51]
  wire  _T_319 = _T_316 & _T_49; // @[el2_ifu_compress_ctl.scala 39:63]
  wire  _T_322 = _T_319 & _T_52; // @[el2_ifu_compress_ctl.scala 39:75]
  wire  _T_325 = _T_322 & _T_248; // @[el2_ifu_compress_ctl.scala 39:87]
  wire  _T_333 = _T_164 & _T_248; // @[el2_ifu_compress_ctl.scala 40:41]
  wire  _T_334 = _T_325 | _T_333; // @[el2_ifu_compress_ctl.scala 40:15]
  wire  _T_338 = _T_4 & io_in[6]; // @[el2_ifu_compress_ctl.scala 40:66]
  wire  _T_341 = _T_338 & _T_248; // @[el2_ifu_compress_ctl.scala 40:75]
  wire  _T_342 = _T_334 | _T_341; // @[el2_ifu_compress_ctl.scala 40:53]
  wire  _T_346 = _T_161 & io_in[14]; // @[el2_ifu_compress_ctl.scala 41:28]
  wire  _T_348 = _T_346 & io_in[0]; // @[el2_ifu_compress_ctl.scala 41:38]
  wire  _T_349 = _T_342 | _T_348; // @[el2_ifu_compress_ctl.scala 41:15]
  wire  _T_353 = _T_4 & io_in[5]; // @[el2_ifu_compress_ctl.scala 41:60]
  wire  _T_356 = _T_353 & _T_248; // @[el2_ifu_compress_ctl.scala 41:69]
  wire  _T_357 = _T_349 | _T_356; // @[el2_ifu_compress_ctl.scala 41:47]
  wire  _T_361 = _T_4 & io_in[4]; // @[el2_ifu_compress_ctl.scala 42:28]
  wire  _T_364 = _T_361 & _T_248; // @[el2_ifu_compress_ctl.scala 42:37]
  wire  _T_365 = _T_357 | _T_364; // @[el2_ifu_compress_ctl.scala 42:15]
  wire  _T_370 = _T_4 & _T_7; // @[el2_ifu_compress_ctl.scala 42:64]
  wire  _T_372 = _T_370 & io_in[0]; // @[el2_ifu_compress_ctl.scala 42:77]
  wire  _T_373 = _T_365 | _T_372; // @[el2_ifu_compress_ctl.scala 42:50]
  wire  _T_377 = _T_4 & io_in[3]; // @[el2_ifu_compress_ctl.scala 43:28]
  wire  _T_380 = _T_377 & _T_248; // @[el2_ifu_compress_ctl.scala 43:37]
  wire  _T_381 = _T_373 | _T_380; // @[el2_ifu_compress_ctl.scala 43:15]
  wire  _T_385 = _T_4 & io_in[2]; // @[el2_ifu_compress_ctl.scala 43:64]
  wire  _T_388 = _T_385 & _T_248; // @[el2_ifu_compress_ctl.scala 43:73]
  wire  _T_389 = _T_381 | _T_388; // @[el2_ifu_compress_ctl.scala 43:50]
  wire  _T_399 = _T_38 & io_in[11]; // @[el2_ifu_compress_ctl.scala 45:35]
  wire  _T_402 = _T_399 & _T_12; // @[el2_ifu_compress_ctl.scala 45:45]
  wire  _T_405 = _T_402 & _T_15; // @[el2_ifu_compress_ctl.scala 45:57]
  wire  _T_408 = _T_405 & _T_61; // @[el2_ifu_compress_ctl.scala 45:69]
  wire  _T_411 = _T_408 & _T_64; // @[el2_ifu_compress_ctl.scala 45:81]
  wire  _T_414 = _T_411 & _T_67; // @[el2_ifu_compress_ctl.scala 45:93]
  wire  _T_416 = _T_414 & io_in[1]; // @[el2_ifu_compress_ctl.scala 45:105]
  wire  _T_422 = _T_38 & io_in[10]; // @[el2_ifu_compress_ctl.scala 46:38]
  wire  _T_425 = _T_422 & _T_12; // @[el2_ifu_compress_ctl.scala 46:48]
  wire  _T_428 = _T_425 & _T_15; // @[el2_ifu_compress_ctl.scala 46:60]
  wire  _T_431 = _T_428 & _T_61; // @[el2_ifu_compress_ctl.scala 46:72]
  wire  _T_434 = _T_431 & _T_64; // @[el2_ifu_compress_ctl.scala 46:84]
  wire  _T_437 = _T_434 & _T_67; // @[el2_ifu_compress_ctl.scala 46:96]
  wire  _T_439 = _T_437 & io_in[1]; // @[el2_ifu_compress_ctl.scala 46:108]
  wire  _T_440 = _T_416 | _T_439; // @[el2_ifu_compress_ctl.scala 46:15]
  wire  _T_446 = _T_38 & io_in[9]; // @[el2_ifu_compress_ctl.scala 47:38]
  wire  _T_449 = _T_446 & _T_12; // @[el2_ifu_compress_ctl.scala 47:47]
  wire  _T_452 = _T_449 & _T_15; // @[el2_ifu_compress_ctl.scala 47:59]
  wire  _T_455 = _T_452 & _T_61; // @[el2_ifu_compress_ctl.scala 47:71]
  wire  _T_458 = _T_455 & _T_64; // @[el2_ifu_compress_ctl.scala 47:83]
  wire  _T_461 = _T_458 & _T_67; // @[el2_ifu_compress_ctl.scala 47:95]
  wire  _T_463 = _T_461 & io_in[1]; // @[el2_ifu_compress_ctl.scala 47:107]
  wire  _T_464 = _T_440 | _T_463; // @[el2_ifu_compress_ctl.scala 47:15]
  wire  _T_470 = _T_38 & io_in[8]; // @[el2_ifu_compress_ctl.scala 48:38]
  wire  _T_473 = _T_470 & _T_12; // @[el2_ifu_compress_ctl.scala 48:47]
  wire  _T_476 = _T_473 & _T_15; // @[el2_ifu_compress_ctl.scala 48:59]
  wire  _T_479 = _T_476 & _T_61; // @[el2_ifu_compress_ctl.scala 48:71]
  wire  _T_482 = _T_479 & _T_64; // @[el2_ifu_compress_ctl.scala 48:83]
  wire  _T_485 = _T_482 & _T_67; // @[el2_ifu_compress_ctl.scala 48:95]
  wire  _T_487 = _T_485 & io_in[1]; // @[el2_ifu_compress_ctl.scala 48:107]
  wire  _T_488 = _T_464 | _T_487; // @[el2_ifu_compress_ctl.scala 48:15]
  wire  _T_494 = _T_38 & io_in[7]; // @[el2_ifu_compress_ctl.scala 49:38]
  wire  _T_497 = _T_494 & _T_12; // @[el2_ifu_compress_ctl.scala 49:47]
  wire  _T_500 = _T_497 & _T_15; // @[el2_ifu_compress_ctl.scala 49:59]
  wire  _T_503 = _T_500 & _T_61; // @[el2_ifu_compress_ctl.scala 49:71]
  wire  _T_506 = _T_503 & _T_64; // @[el2_ifu_compress_ctl.scala 49:83]
  wire  _T_509 = _T_506 & _T_67; // @[el2_ifu_compress_ctl.scala 49:95]
  wire  _T_511 = _T_509 & io_in[1]; // @[el2_ifu_compress_ctl.scala 49:107]
  wire  _T_512 = _T_488 | _T_511; // @[el2_ifu_compress_ctl.scala 49:15]
  wire  _T_518 = ~io_in[12]; // @[el2_ifu_compress_ctl.scala 50:40]
  wire  _T_519 = _T_5 & _T_518; // @[el2_ifu_compress_ctl.scala 50:38]
  wire  _T_522 = _T_519 & _T_12; // @[el2_ifu_compress_ctl.scala 50:51]
  wire  _T_525 = _T_522 & _T_15; // @[el2_ifu_compress_ctl.scala 50:63]
  wire  _T_528 = _T_525 & _T_61; // @[el2_ifu_compress_ctl.scala 50:75]
  wire  _T_531 = _T_528 & _T_64; // @[el2_ifu_compress_ctl.scala 50:87]
  wire  _T_534 = _T_531 & _T_67; // @[el2_ifu_compress_ctl.scala 50:99]
  wire  _T_537 = _T_534 & _T_248; // @[el2_ifu_compress_ctl.scala 50:111]
  wire  _T_538 = _T_512 | _T_537; // @[el2_ifu_compress_ctl.scala 50:15]
  wire  _T_542 = _T_161 & io_in[13]; // @[el2_ifu_compress_ctl.scala 51:28]
  wire  _T_545 = _T_542 & _T_49; // @[el2_ifu_compress_ctl.scala 51:38]
  wire  _T_546 = _T_538 | _T_545; // @[el2_ifu_compress_ctl.scala 51:15]
  wire  _T_552 = _T_542 & io_in[7]; // @[el2_ifu_compress_ctl.scala 51:75]
  wire  _T_553 = _T_546 | _T_552; // @[el2_ifu_compress_ctl.scala 51:51]
  wire  _T_559 = _T_542 & io_in[9]; // @[el2_ifu_compress_ctl.scala 51:109]
  wire  _T_560 = _T_553 | _T_559; // @[el2_ifu_compress_ctl.scala 51:85]
  wire  _T_566 = _T_542 & io_in[10]; // @[el2_ifu_compress_ctl.scala 52:38]
  wire  _T_567 = _T_560 | _T_566; // @[el2_ifu_compress_ctl.scala 52:15]
  wire  _T_573 = _T_542 & io_in[11]; // @[el2_ifu_compress_ctl.scala 52:73]
  wire  _T_574 = _T_567 | _T_573; // @[el2_ifu_compress_ctl.scala 52:49]
  wire  _T_579 = _T_574 | _T_253; // @[el2_ifu_compress_ctl.scala 52:84]
  wire [11:0] _T_586 = {5'h0,_T_260,_T_305,_T_389,_T_253,_T_579,2'h3}; // @[Cat.scala 29:58]
  wire [19:0] _T_593 = {1'h0,_T_33,9'h0,_T_70,5'h0,_T_120,_T_173,_T_173}; // @[Cat.scala 29:58]
  assign io_out = {_T_593,_T_586}; // @[el2_ifu_compress_ctl.scala 111:10]
endmodule
