module inv_sbox(
  input        clock,
  input        reset,
  input  [7:0] io_byte_in,
  output [7:0] io_byte_out
);
  wire  _T = io_byte_in == 8'h0; // @[cipher.scala 63:56]
  wire  _T_1 = io_byte_in == 8'h1; // @[cipher.scala 63:56]
  wire  _T_2 = io_byte_in == 8'h2; // @[cipher.scala 63:56]
  wire  _T_3 = io_byte_in == 8'h3; // @[cipher.scala 63:56]
  wire  _T_4 = io_byte_in == 8'h4; // @[cipher.scala 63:56]
  wire  _T_5 = io_byte_in == 8'h5; // @[cipher.scala 63:56]
  wire  _T_6 = io_byte_in == 8'h6; // @[cipher.scala 63:56]
  wire  _T_7 = io_byte_in == 8'h7; // @[cipher.scala 63:56]
  wire  _T_8 = io_byte_in == 8'h8; // @[cipher.scala 63:56]
  wire  _T_9 = io_byte_in == 8'h9; // @[cipher.scala 63:56]
  wire  _T_10 = io_byte_in == 8'ha; // @[cipher.scala 63:56]
  wire  _T_11 = io_byte_in == 8'hb; // @[cipher.scala 63:56]
  wire  _T_12 = io_byte_in == 8'hc; // @[cipher.scala 63:56]
  wire  _T_13 = io_byte_in == 8'hd; // @[cipher.scala 63:56]
  wire  _T_14 = io_byte_in == 8'he; // @[cipher.scala 63:56]
  wire  _T_15 = io_byte_in == 8'hf; // @[cipher.scala 63:56]
  wire  _T_16 = io_byte_in == 8'h10; // @[cipher.scala 63:56]
  wire  _T_17 = io_byte_in == 8'h11; // @[cipher.scala 63:56]
  wire  _T_18 = io_byte_in == 8'h12; // @[cipher.scala 63:56]
  wire  _T_19 = io_byte_in == 8'h13; // @[cipher.scala 63:56]
  wire  _T_20 = io_byte_in == 8'h14; // @[cipher.scala 63:56]
  wire  _T_21 = io_byte_in == 8'h15; // @[cipher.scala 63:56]
  wire  _T_22 = io_byte_in == 8'h16; // @[cipher.scala 63:56]
  wire  _T_23 = io_byte_in == 8'h17; // @[cipher.scala 63:56]
  wire  _T_24 = io_byte_in == 8'h18; // @[cipher.scala 63:56]
  wire  _T_25 = io_byte_in == 8'h19; // @[cipher.scala 63:56]
  wire  _T_26 = io_byte_in == 8'h1a; // @[cipher.scala 63:56]
  wire  _T_27 = io_byte_in == 8'h1b; // @[cipher.scala 63:56]
  wire  _T_28 = io_byte_in == 8'h1c; // @[cipher.scala 63:56]
  wire  _T_29 = io_byte_in == 8'h1d; // @[cipher.scala 63:56]
  wire  _T_30 = io_byte_in == 8'h1e; // @[cipher.scala 63:56]
  wire  _T_31 = io_byte_in == 8'h1f; // @[cipher.scala 63:56]
  wire  _T_32 = io_byte_in == 8'h20; // @[cipher.scala 63:56]
  wire  _T_33 = io_byte_in == 8'h21; // @[cipher.scala 63:56]
  wire  _T_34 = io_byte_in == 8'h22; // @[cipher.scala 63:56]
  wire  _T_35 = io_byte_in == 8'h23; // @[cipher.scala 63:56]
  wire  _T_36 = io_byte_in == 8'h24; // @[cipher.scala 63:56]
  wire  _T_37 = io_byte_in == 8'h25; // @[cipher.scala 63:56]
  wire  _T_38 = io_byte_in == 8'h26; // @[cipher.scala 63:56]
  wire  _T_39 = io_byte_in == 8'h27; // @[cipher.scala 63:56]
  wire  _T_40 = io_byte_in == 8'h28; // @[cipher.scala 63:56]
  wire  _T_41 = io_byte_in == 8'h29; // @[cipher.scala 63:56]
  wire  _T_42 = io_byte_in == 8'h2a; // @[cipher.scala 63:56]
  wire  _T_43 = io_byte_in == 8'h2b; // @[cipher.scala 63:56]
  wire  _T_44 = io_byte_in == 8'h2c; // @[cipher.scala 63:56]
  wire  _T_45 = io_byte_in == 8'h2d; // @[cipher.scala 63:56]
  wire  _T_46 = io_byte_in == 8'h2e; // @[cipher.scala 63:56]
  wire  _T_47 = io_byte_in == 8'h2f; // @[cipher.scala 63:56]
  wire  _T_48 = io_byte_in == 8'h30; // @[cipher.scala 63:56]
  wire  _T_49 = io_byte_in == 8'h31; // @[cipher.scala 63:56]
  wire  _T_50 = io_byte_in == 8'h32; // @[cipher.scala 63:56]
  wire  _T_51 = io_byte_in == 8'h33; // @[cipher.scala 63:56]
  wire  _T_52 = io_byte_in == 8'h34; // @[cipher.scala 63:56]
  wire  _T_53 = io_byte_in == 8'h35; // @[cipher.scala 63:56]
  wire  _T_54 = io_byte_in == 8'h36; // @[cipher.scala 63:56]
  wire  _T_55 = io_byte_in == 8'h37; // @[cipher.scala 63:56]
  wire  _T_56 = io_byte_in == 8'h38; // @[cipher.scala 63:56]
  wire  _T_57 = io_byte_in == 8'h39; // @[cipher.scala 63:56]
  wire  _T_58 = io_byte_in == 8'h3a; // @[cipher.scala 63:56]
  wire  _T_59 = io_byte_in == 8'h3b; // @[cipher.scala 63:56]
  wire  _T_60 = io_byte_in == 8'h3c; // @[cipher.scala 63:56]
  wire  _T_61 = io_byte_in == 8'h3d; // @[cipher.scala 63:56]
  wire  _T_62 = io_byte_in == 8'h3e; // @[cipher.scala 63:56]
  wire  _T_63 = io_byte_in == 8'h3f; // @[cipher.scala 63:56]
  wire  _T_64 = io_byte_in == 8'h40; // @[cipher.scala 63:56]
  wire  _T_65 = io_byte_in == 8'h41; // @[cipher.scala 63:56]
  wire  _T_66 = io_byte_in == 8'h42; // @[cipher.scala 63:56]
  wire  _T_67 = io_byte_in == 8'h43; // @[cipher.scala 63:56]
  wire  _T_68 = io_byte_in == 8'h44; // @[cipher.scala 63:56]
  wire  _T_69 = io_byte_in == 8'h45; // @[cipher.scala 63:56]
  wire  _T_70 = io_byte_in == 8'h46; // @[cipher.scala 63:56]
  wire  _T_71 = io_byte_in == 8'h47; // @[cipher.scala 63:56]
  wire  _T_72 = io_byte_in == 8'h48; // @[cipher.scala 63:56]
  wire  _T_73 = io_byte_in == 8'h49; // @[cipher.scala 63:56]
  wire  _T_74 = io_byte_in == 8'h4a; // @[cipher.scala 63:56]
  wire  _T_75 = io_byte_in == 8'h4b; // @[cipher.scala 63:56]
  wire  _T_76 = io_byte_in == 8'h4c; // @[cipher.scala 63:56]
  wire  _T_77 = io_byte_in == 8'h4d; // @[cipher.scala 63:56]
  wire  _T_78 = io_byte_in == 8'h4e; // @[cipher.scala 63:56]
  wire  _T_79 = io_byte_in == 8'h4f; // @[cipher.scala 63:56]
  wire  _T_80 = io_byte_in == 8'h50; // @[cipher.scala 63:56]
  wire  _T_81 = io_byte_in == 8'h51; // @[cipher.scala 63:56]
  wire  _T_82 = io_byte_in == 8'h52; // @[cipher.scala 63:56]
  wire  _T_83 = io_byte_in == 8'h53; // @[cipher.scala 63:56]
  wire  _T_84 = io_byte_in == 8'h54; // @[cipher.scala 63:56]
  wire  _T_85 = io_byte_in == 8'h55; // @[cipher.scala 63:56]
  wire  _T_86 = io_byte_in == 8'h56; // @[cipher.scala 63:56]
  wire  _T_87 = io_byte_in == 8'h57; // @[cipher.scala 63:56]
  wire  _T_88 = io_byte_in == 8'h58; // @[cipher.scala 63:56]
  wire  _T_89 = io_byte_in == 8'h59; // @[cipher.scala 63:56]
  wire  _T_90 = io_byte_in == 8'h5a; // @[cipher.scala 63:56]
  wire  _T_91 = io_byte_in == 8'h5b; // @[cipher.scala 63:56]
  wire  _T_92 = io_byte_in == 8'h5c; // @[cipher.scala 63:56]
  wire  _T_93 = io_byte_in == 8'h5d; // @[cipher.scala 63:56]
  wire  _T_94 = io_byte_in == 8'h5e; // @[cipher.scala 63:56]
  wire  _T_95 = io_byte_in == 8'h5f; // @[cipher.scala 63:56]
  wire  _T_96 = io_byte_in == 8'h60; // @[cipher.scala 63:56]
  wire  _T_97 = io_byte_in == 8'h61; // @[cipher.scala 63:56]
  wire  _T_98 = io_byte_in == 8'h62; // @[cipher.scala 63:56]
  wire  _T_100 = io_byte_in == 8'h64; // @[cipher.scala 63:56]
  wire  _T_101 = io_byte_in == 8'h65; // @[cipher.scala 63:56]
  wire  _T_102 = io_byte_in == 8'h66; // @[cipher.scala 63:56]
  wire  _T_103 = io_byte_in == 8'h67; // @[cipher.scala 63:56]
  wire  _T_104 = io_byte_in == 8'h68; // @[cipher.scala 63:56]
  wire  _T_105 = io_byte_in == 8'h69; // @[cipher.scala 63:56]
  wire  _T_106 = io_byte_in == 8'h6a; // @[cipher.scala 63:56]
  wire  _T_107 = io_byte_in == 8'h6b; // @[cipher.scala 63:56]
  wire  _T_108 = io_byte_in == 8'h6c; // @[cipher.scala 63:56]
  wire  _T_109 = io_byte_in == 8'h6d; // @[cipher.scala 63:56]
  wire  _T_110 = io_byte_in == 8'h6e; // @[cipher.scala 63:56]
  wire  _T_111 = io_byte_in == 8'h6f; // @[cipher.scala 63:56]
  wire  _T_112 = io_byte_in == 8'h70; // @[cipher.scala 63:56]
  wire  _T_113 = io_byte_in == 8'h71; // @[cipher.scala 63:56]
  wire  _T_114 = io_byte_in == 8'h72; // @[cipher.scala 63:56]
  wire  _T_115 = io_byte_in == 8'h73; // @[cipher.scala 63:56]
  wire  _T_116 = io_byte_in == 8'h74; // @[cipher.scala 63:56]
  wire  _T_117 = io_byte_in == 8'h75; // @[cipher.scala 63:56]
  wire  _T_118 = io_byte_in == 8'h76; // @[cipher.scala 63:56]
  wire  _T_119 = io_byte_in == 8'h77; // @[cipher.scala 63:56]
  wire  _T_120 = io_byte_in == 8'h78; // @[cipher.scala 63:56]
  wire  _T_121 = io_byte_in == 8'h79; // @[cipher.scala 63:56]
  wire  _T_122 = io_byte_in == 8'h7a; // @[cipher.scala 63:56]
  wire  _T_123 = io_byte_in == 8'h7b; // @[cipher.scala 63:56]
  wire  _T_124 = io_byte_in == 8'h7c; // @[cipher.scala 63:56]
  wire  _T_125 = io_byte_in == 8'h7d; // @[cipher.scala 63:56]
  wire  _T_126 = io_byte_in == 8'h7e; // @[cipher.scala 63:56]
  wire  _T_127 = io_byte_in == 8'h7f; // @[cipher.scala 63:56]
  wire  _T_128 = io_byte_in == 8'h80; // @[cipher.scala 63:56]
  wire  _T_129 = io_byte_in == 8'h81; // @[cipher.scala 63:56]
  wire  _T_130 = io_byte_in == 8'h82; // @[cipher.scala 63:56]
  wire  _T_131 = io_byte_in == 8'h83; // @[cipher.scala 63:56]
  wire  _T_132 = io_byte_in == 8'h84; // @[cipher.scala 63:56]
  wire  _T_133 = io_byte_in == 8'h85; // @[cipher.scala 63:56]
  wire  _T_134 = io_byte_in == 8'h86; // @[cipher.scala 63:56]
  wire  _T_135 = io_byte_in == 8'h87; // @[cipher.scala 63:56]
  wire  _T_136 = io_byte_in == 8'h88; // @[cipher.scala 63:56]
  wire  _T_137 = io_byte_in == 8'h89; // @[cipher.scala 63:56]
  wire  _T_138 = io_byte_in == 8'h8a; // @[cipher.scala 63:56]
  wire  _T_139 = io_byte_in == 8'h8b; // @[cipher.scala 63:56]
  wire  _T_140 = io_byte_in == 8'h8c; // @[cipher.scala 63:56]
  wire  _T_141 = io_byte_in == 8'h8d; // @[cipher.scala 63:56]
  wire  _T_142 = io_byte_in == 8'h8e; // @[cipher.scala 63:56]
  wire  _T_143 = io_byte_in == 8'h8f; // @[cipher.scala 63:56]
  wire  _T_144 = io_byte_in == 8'h90; // @[cipher.scala 63:56]
  wire  _T_145 = io_byte_in == 8'h91; // @[cipher.scala 63:56]
  wire  _T_146 = io_byte_in == 8'h92; // @[cipher.scala 63:56]
  wire  _T_147 = io_byte_in == 8'h93; // @[cipher.scala 63:56]
  wire  _T_148 = io_byte_in == 8'h94; // @[cipher.scala 63:56]
  wire  _T_149 = io_byte_in == 8'h95; // @[cipher.scala 63:56]
  wire  _T_150 = io_byte_in == 8'h96; // @[cipher.scala 63:56]
  wire  _T_151 = io_byte_in == 8'h97; // @[cipher.scala 63:56]
  wire  _T_152 = io_byte_in == 8'h98; // @[cipher.scala 63:56]
  wire  _T_153 = io_byte_in == 8'h99; // @[cipher.scala 63:56]
  wire  _T_154 = io_byte_in == 8'h9a; // @[cipher.scala 63:56]
  wire  _T_155 = io_byte_in == 8'h9b; // @[cipher.scala 63:56]
  wire  _T_156 = io_byte_in == 8'h9c; // @[cipher.scala 63:56]
  wire  _T_157 = io_byte_in == 8'h9d; // @[cipher.scala 63:56]
  wire  _T_158 = io_byte_in == 8'h9e; // @[cipher.scala 63:56]
  wire  _T_159 = io_byte_in == 8'h9f; // @[cipher.scala 63:56]
  wire  _T_160 = io_byte_in == 8'ha0; // @[cipher.scala 63:56]
  wire  _T_161 = io_byte_in == 8'ha1; // @[cipher.scala 63:56]
  wire  _T_162 = io_byte_in == 8'ha2; // @[cipher.scala 63:56]
  wire  _T_163 = io_byte_in == 8'ha3; // @[cipher.scala 63:56]
  wire  _T_164 = io_byte_in == 8'ha4; // @[cipher.scala 63:56]
  wire  _T_165 = io_byte_in == 8'ha5; // @[cipher.scala 63:56]
  wire  _T_166 = io_byte_in == 8'ha6; // @[cipher.scala 63:56]
  wire  _T_167 = io_byte_in == 8'ha7; // @[cipher.scala 63:56]
  wire  _T_168 = io_byte_in == 8'ha8; // @[cipher.scala 63:56]
  wire  _T_169 = io_byte_in == 8'ha9; // @[cipher.scala 63:56]
  wire  _T_170 = io_byte_in == 8'haa; // @[cipher.scala 63:56]
  wire  _T_171 = io_byte_in == 8'hab; // @[cipher.scala 63:56]
  wire  _T_172 = io_byte_in == 8'hac; // @[cipher.scala 63:56]
  wire  _T_173 = io_byte_in == 8'had; // @[cipher.scala 63:56]
  wire  _T_174 = io_byte_in == 8'hae; // @[cipher.scala 63:56]
  wire  _T_175 = io_byte_in == 8'haf; // @[cipher.scala 63:56]
  wire  _T_176 = io_byte_in == 8'hb0; // @[cipher.scala 63:56]
  wire  _T_177 = io_byte_in == 8'hb1; // @[cipher.scala 63:56]
  wire  _T_178 = io_byte_in == 8'hb2; // @[cipher.scala 63:56]
  wire  _T_179 = io_byte_in == 8'hb3; // @[cipher.scala 63:56]
  wire  _T_180 = io_byte_in == 8'hb4; // @[cipher.scala 63:56]
  wire  _T_181 = io_byte_in == 8'hb5; // @[cipher.scala 63:56]
  wire  _T_182 = io_byte_in == 8'hb6; // @[cipher.scala 63:56]
  wire  _T_183 = io_byte_in == 8'hb7; // @[cipher.scala 63:56]
  wire  _T_184 = io_byte_in == 8'hb8; // @[cipher.scala 63:56]
  wire  _T_185 = io_byte_in == 8'hb9; // @[cipher.scala 63:56]
  wire  _T_186 = io_byte_in == 8'hba; // @[cipher.scala 63:56]
  wire  _T_187 = io_byte_in == 8'hbb; // @[cipher.scala 63:56]
  wire  _T_188 = io_byte_in == 8'hbc; // @[cipher.scala 63:56]
  wire  _T_189 = io_byte_in == 8'hbd; // @[cipher.scala 63:56]
  wire  _T_190 = io_byte_in == 8'hbe; // @[cipher.scala 63:56]
  wire  _T_191 = io_byte_in == 8'hbf; // @[cipher.scala 63:56]
  wire  _T_192 = io_byte_in == 8'hc0; // @[cipher.scala 63:56]
  wire  _T_193 = io_byte_in == 8'hc1; // @[cipher.scala 63:56]
  wire  _T_194 = io_byte_in == 8'hc2; // @[cipher.scala 63:56]
  wire  _T_195 = io_byte_in == 8'hc3; // @[cipher.scala 63:56]
  wire  _T_196 = io_byte_in == 8'hc4; // @[cipher.scala 63:56]
  wire  _T_197 = io_byte_in == 8'hc5; // @[cipher.scala 63:56]
  wire  _T_198 = io_byte_in == 8'hc6; // @[cipher.scala 63:56]
  wire  _T_199 = io_byte_in == 8'hc7; // @[cipher.scala 63:56]
  wire  _T_200 = io_byte_in == 8'hc8; // @[cipher.scala 63:56]
  wire  _T_201 = io_byte_in == 8'hc9; // @[cipher.scala 63:56]
  wire  _T_202 = io_byte_in == 8'hca; // @[cipher.scala 63:56]
  wire  _T_203 = io_byte_in == 8'hcb; // @[cipher.scala 63:56]
  wire  _T_204 = io_byte_in == 8'hcc; // @[cipher.scala 63:56]
  wire  _T_205 = io_byte_in == 8'hcd; // @[cipher.scala 63:56]
  wire  _T_206 = io_byte_in == 8'hce; // @[cipher.scala 63:56]
  wire  _T_207 = io_byte_in == 8'hcf; // @[cipher.scala 63:56]
  wire  _T_208 = io_byte_in == 8'hd0; // @[cipher.scala 63:56]
  wire  _T_209 = io_byte_in == 8'hd1; // @[cipher.scala 63:56]
  wire  _T_210 = io_byte_in == 8'hd2; // @[cipher.scala 63:56]
  wire  _T_211 = io_byte_in == 8'hd3; // @[cipher.scala 63:56]
  wire  _T_212 = io_byte_in == 8'hd4; // @[cipher.scala 63:56]
  wire  _T_213 = io_byte_in == 8'hd5; // @[cipher.scala 63:56]
  wire  _T_214 = io_byte_in == 8'hd6; // @[cipher.scala 63:56]
  wire  _T_215 = io_byte_in == 8'hd7; // @[cipher.scala 63:56]
  wire  _T_216 = io_byte_in == 8'hd8; // @[cipher.scala 63:56]
  wire  _T_217 = io_byte_in == 8'hd9; // @[cipher.scala 63:56]
  wire  _T_218 = io_byte_in == 8'hda; // @[cipher.scala 63:56]
  wire  _T_219 = io_byte_in == 8'hdb; // @[cipher.scala 63:56]
  wire  _T_220 = io_byte_in == 8'hdc; // @[cipher.scala 63:56]
  wire  _T_221 = io_byte_in == 8'hdd; // @[cipher.scala 63:56]
  wire  _T_222 = io_byte_in == 8'hde; // @[cipher.scala 63:56]
  wire  _T_223 = io_byte_in == 8'hdf; // @[cipher.scala 63:56]
  wire  _T_224 = io_byte_in == 8'he0; // @[cipher.scala 63:56]
  wire  _T_225 = io_byte_in == 8'he1; // @[cipher.scala 63:56]
  wire  _T_226 = io_byte_in == 8'he2; // @[cipher.scala 63:56]
  wire  _T_227 = io_byte_in == 8'he3; // @[cipher.scala 63:56]
  wire  _T_228 = io_byte_in == 8'he4; // @[cipher.scala 63:56]
  wire  _T_229 = io_byte_in == 8'he5; // @[cipher.scala 63:56]
  wire  _T_230 = io_byte_in == 8'he6; // @[cipher.scala 63:56]
  wire  _T_231 = io_byte_in == 8'he7; // @[cipher.scala 63:56]
  wire  _T_232 = io_byte_in == 8'he8; // @[cipher.scala 63:56]
  wire  _T_233 = io_byte_in == 8'he9; // @[cipher.scala 63:56]
  wire  _T_234 = io_byte_in == 8'hea; // @[cipher.scala 63:56]
  wire  _T_235 = io_byte_in == 8'heb; // @[cipher.scala 63:56]
  wire  _T_236 = io_byte_in == 8'hec; // @[cipher.scala 63:56]
  wire  _T_237 = io_byte_in == 8'hed; // @[cipher.scala 63:56]
  wire  _T_238 = io_byte_in == 8'hee; // @[cipher.scala 63:56]
  wire  _T_239 = io_byte_in == 8'hef; // @[cipher.scala 63:56]
  wire  _T_240 = io_byte_in == 8'hf0; // @[cipher.scala 63:56]
  wire  _T_241 = io_byte_in == 8'hf1; // @[cipher.scala 63:56]
  wire  _T_242 = io_byte_in == 8'hf2; // @[cipher.scala 63:56]
  wire  _T_243 = io_byte_in == 8'hf3; // @[cipher.scala 63:56]
  wire  _T_244 = io_byte_in == 8'hf4; // @[cipher.scala 63:56]
  wire  _T_245 = io_byte_in == 8'hf5; // @[cipher.scala 63:56]
  wire  _T_246 = io_byte_in == 8'hf6; // @[cipher.scala 63:56]
  wire  _T_247 = io_byte_in == 8'hf7; // @[cipher.scala 63:56]
  wire  _T_248 = io_byte_in == 8'hf8; // @[cipher.scala 63:56]
  wire  _T_249 = io_byte_in == 8'hf9; // @[cipher.scala 63:56]
  wire  _T_250 = io_byte_in == 8'hfa; // @[cipher.scala 63:56]
  wire  _T_251 = io_byte_in == 8'hfb; // @[cipher.scala 63:56]
  wire  _T_252 = io_byte_in == 8'hfc; // @[cipher.scala 63:56]
  wire  _T_253 = io_byte_in == 8'hfd; // @[cipher.scala 63:56]
  wire  _T_254 = io_byte_in == 8'hfe; // @[cipher.scala 63:56]
  wire  _T_255 = io_byte_in == 8'hff; // @[cipher.scala 63:56]
  wire [6:0] _T_256 = _T ? 7'h52 : 7'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_257 = _T_1 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_258 = _T_2 ? 7'h6a : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_259 = _T_3 ? 8'hd5 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_260 = _T_4 ? 6'h30 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_261 = _T_5 ? 6'h36 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_262 = _T_6 ? 8'ha5 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_263 = _T_7 ? 6'h38 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_264 = _T_8 ? 8'hbf : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_265 = _T_9 ? 7'h40 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_266 = _T_10 ? 8'ha3 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_267 = _T_11 ? 8'h9e : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_268 = _T_12 ? 8'h81 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_269 = _T_13 ? 8'hf3 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_270 = _T_14 ? 8'hd7 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_271 = _T_15 ? 8'hfb : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_272 = _T_16 ? 7'h7c : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_273 = _T_17 ? 8'he3 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_274 = _T_18 ? 6'h39 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_275 = _T_19 ? 8'h82 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_276 = _T_20 ? 8'h9b : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_277 = _T_21 ? 6'h2f : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_278 = _T_22 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_279 = _T_23 ? 8'h87 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_280 = _T_24 ? 6'h34 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_281 = _T_25 ? 8'h8e : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_282 = _T_26 ? 7'h43 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_283 = _T_27 ? 7'h44 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_284 = _T_28 ? 8'hc4 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_285 = _T_29 ? 8'hde : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_286 = _T_30 ? 8'he9 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_287 = _T_31 ? 8'hcb : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_288 = _T_32 ? 7'h54 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_289 = _T_33 ? 7'h7b : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_290 = _T_34 ? 8'h94 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_291 = _T_35 ? 6'h32 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_292 = _T_36 ? 8'ha6 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_293 = _T_37 ? 8'hc2 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_294 = _T_38 ? 6'h23 : 6'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_295 = _T_39 ? 6'h3d : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_296 = _T_40 ? 8'hee : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_297 = _T_41 ? 7'h4c : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_298 = _T_42 ? 8'h95 : 8'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_299 = _T_43 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_300 = _T_44 ? 7'h42 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_301 = _T_45 ? 8'hfa : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_302 = _T_46 ? 8'hc3 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_303 = _T_47 ? 7'h4e : 7'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_304 = _T_48 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_305 = _T_49 ? 6'h2e : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_306 = _T_50 ? 8'ha1 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_307 = _T_51 ? 7'h66 : 7'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_308 = _T_52 ? 6'h28 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_309 = _T_53 ? 8'hd9 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_310 = _T_54 ? 6'h24 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_311 = _T_55 ? 8'hb2 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_312 = _T_56 ? 7'h76 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_313 = _T_57 ? 7'h5b : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_314 = _T_58 ? 8'ha2 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_315 = _T_59 ? 7'h49 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_316 = _T_60 ? 7'h6d : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_317 = _T_61 ? 8'h8b : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_318 = _T_62 ? 8'hd1 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_319 = _T_63 ? 6'h25 : 6'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_320 = _T_64 ? 7'h72 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_321 = _T_65 ? 8'hf8 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_322 = _T_66 ? 8'hf6 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_323 = _T_67 ? 7'h64 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_324 = _T_68 ? 8'h86 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_325 = _T_69 ? 7'h68 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_326 = _T_70 ? 8'h98 : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_327 = _T_71 ? 5'h16 : 5'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_328 = _T_72 ? 8'hd4 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_329 = _T_73 ? 8'ha4 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_330 = _T_74 ? 7'h5c : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_331 = _T_75 ? 8'hcc : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_332 = _T_76 ? 7'h5d : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_333 = _T_77 ? 7'h65 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_334 = _T_78 ? 8'hb6 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_335 = _T_79 ? 8'h92 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_336 = _T_80 ? 7'h6c : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_337 = _T_81 ? 7'h70 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_338 = _T_82 ? 7'h48 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_339 = _T_83 ? 7'h50 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_340 = _T_84 ? 8'hfd : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_341 = _T_85 ? 8'hed : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_342 = _T_86 ? 8'hb9 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_343 = _T_87 ? 8'hda : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_344 = _T_88 ? 7'h5e : 7'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_345 = _T_89 ? 5'h15 : 5'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_346 = _T_90 ? 7'h46 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_347 = _T_91 ? 7'h57 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_348 = _T_92 ? 8'ha7 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_349 = _T_93 ? 8'h8d : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_350 = _T_94 ? 8'h9d : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_351 = _T_95 ? 8'h84 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_352 = _T_96 ? 8'h90 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_353 = _T_97 ? 8'hd8 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_354 = _T_98 ? 8'hab : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_356 = _T_100 ? 8'h8c : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_357 = _T_101 ? 8'hbc : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_358 = _T_102 ? 8'hd3 : 8'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_359 = _T_103 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_360 = _T_104 ? 8'hf7 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_361 = _T_105 ? 8'he4 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_362 = _T_106 ? 7'h58 : 7'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_363 = _T_107 ? 3'h5 : 3'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_364 = _T_108 ? 8'hb8 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_365 = _T_109 ? 8'hb3 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_366 = _T_110 ? 7'h45 : 7'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_367 = _T_111 ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_368 = _T_112 ? 8'hd0 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_369 = _T_113 ? 6'h2c : 6'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_370 = _T_114 ? 5'h1e : 5'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_371 = _T_115 ? 8'h8f : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_372 = _T_116 ? 8'hca : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_373 = _T_117 ? 6'h3f : 6'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_374 = _T_118 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_375 = _T_119 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_376 = _T_120 ? 8'hc1 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_377 = _T_121 ? 8'haf : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_378 = _T_122 ? 8'hbd : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_379 = _T_123 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_381 = _T_125 ? 5'h13 : 5'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_382 = _T_126 ? 8'h8a : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_383 = _T_127 ? 7'h6b : 7'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_384 = _T_128 ? 6'h3a : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_385 = _T_129 ? 8'h91 : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_386 = _T_130 ? 5'h11 : 5'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_387 = _T_131 ? 7'h41 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_388 = _T_132 ? 7'h4f : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_389 = _T_133 ? 7'h67 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_390 = _T_134 ? 8'hdc : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_391 = _T_135 ? 8'hea : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_392 = _T_136 ? 8'h97 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_393 = _T_137 ? 8'hf2 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_394 = _T_138 ? 8'hcf : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_395 = _T_139 ? 8'hce : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_396 = _T_140 ? 8'hf0 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_397 = _T_141 ? 8'hb4 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_398 = _T_142 ? 8'he6 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_399 = _T_143 ? 7'h73 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_400 = _T_144 ? 8'h96 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_401 = _T_145 ? 8'hac : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_402 = _T_146 ? 7'h74 : 7'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_403 = _T_147 ? 6'h22 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_404 = _T_148 ? 8'he7 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_405 = _T_149 ? 8'had : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_406 = _T_150 ? 6'h35 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_407 = _T_151 ? 8'h85 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_408 = _T_152 ? 8'he2 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_409 = _T_153 ? 8'hf9 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_410 = _T_154 ? 6'h37 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_411 = _T_155 ? 8'he8 : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_412 = _T_156 ? 5'h1c : 5'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_413 = _T_157 ? 7'h75 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_414 = _T_158 ? 8'hdf : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_415 = _T_159 ? 7'h6e : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_416 = _T_160 ? 7'h47 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_417 = _T_161 ? 8'hf1 : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_418 = _T_162 ? 5'h1a : 5'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_419 = _T_163 ? 7'h71 : 7'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_420 = _T_164 ? 5'h1d : 5'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_421 = _T_165 ? 6'h29 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_422 = _T_166 ? 8'hc5 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_423 = _T_167 ? 8'h89 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_424 = _T_168 ? 7'h6f : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_425 = _T_169 ? 8'hb7 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_426 = _T_170 ? 7'h62 : 7'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_427 = _T_171 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_428 = _T_172 ? 8'haa : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_429 = _T_173 ? 5'h18 : 5'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_430 = _T_174 ? 8'hbe : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_431 = _T_175 ? 5'h1b : 5'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_432 = _T_176 ? 8'hfc : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_433 = _T_177 ? 7'h56 : 7'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_434 = _T_178 ? 6'h3e : 6'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_435 = _T_179 ? 7'h4b : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_436 = _T_180 ? 8'hc6 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_437 = _T_181 ? 8'hd2 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_438 = _T_182 ? 7'h79 : 7'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_439 = _T_183 ? 6'h20 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_440 = _T_184 ? 8'h9a : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_441 = _T_185 ? 8'hdb : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_442 = _T_186 ? 8'hc0 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_443 = _T_187 ? 8'hfe : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_444 = _T_188 ? 7'h78 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_445 = _T_189 ? 8'hcd : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_446 = _T_190 ? 7'h5a : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_447 = _T_191 ? 8'hf4 : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_448 = _T_192 ? 5'h1f : 5'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_449 = _T_193 ? 8'hdd : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_450 = _T_194 ? 8'ha8 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_451 = _T_195 ? 6'h33 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_452 = _T_196 ? 8'h88 : 8'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_453 = _T_197 ? 3'h7 : 3'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_454 = _T_198 ? 8'hc7 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_455 = _T_199 ? 6'h31 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_456 = _T_200 ? 8'hb1 : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_457 = _T_201 ? 5'h12 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_458 = _T_202 ? 5'h10 : 5'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_459 = _T_203 ? 7'h59 : 7'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_460 = _T_204 ? 6'h27 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_461 = _T_205 ? 8'h80 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_462 = _T_206 ? 8'hec : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_463 = _T_207 ? 7'h5f : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_464 = _T_208 ? 7'h60 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_465 = _T_209 ? 7'h51 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_466 = _T_210 ? 7'h7f : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_467 = _T_211 ? 8'ha9 : 8'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_468 = _T_212 ? 5'h19 : 5'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_469 = _T_213 ? 8'hb5 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_470 = _T_214 ? 7'h4a : 7'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_471 = _T_215 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_472 = _T_216 ? 6'h2d : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_473 = _T_217 ? 8'he5 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_474 = _T_218 ? 7'h7a : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_475 = _T_219 ? 8'h9f : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_476 = _T_220 ? 8'h93 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_477 = _T_221 ? 8'hc9 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_478 = _T_222 ? 8'h9c : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_479 = _T_223 ? 8'hef : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_480 = _T_224 ? 8'ha0 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_481 = _T_225 ? 8'he0 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_482 = _T_226 ? 6'h3b : 6'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_483 = _T_227 ? 7'h4d : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_484 = _T_228 ? 8'hae : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_485 = _T_229 ? 6'h2a : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_486 = _T_230 ? 8'hf5 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_487 = _T_231 ? 8'hb0 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_488 = _T_232 ? 8'hc8 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_489 = _T_233 ? 8'heb : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_490 = _T_234 ? 8'hbb : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_491 = _T_235 ? 6'h3c : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_492 = _T_236 ? 8'h83 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_493 = _T_237 ? 7'h53 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_494 = _T_238 ? 8'h99 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_495 = _T_239 ? 7'h61 : 7'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_496 = _T_240 ? 5'h17 : 5'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_497 = _T_241 ? 6'h2b : 6'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_498 = _T_242 ? 3'h4 : 3'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_499 = _T_243 ? 7'h7e : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_500 = _T_244 ? 8'hba : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_501 = _T_245 ? 7'h77 : 7'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_502 = _T_246 ? 8'hd6 : 8'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_503 = _T_247 ? 6'h26 : 6'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_504 = _T_248 ? 8'he1 : 8'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_505 = _T_249 ? 7'h69 : 7'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_506 = _T_250 ? 5'h14 : 5'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_507 = _T_251 ? 7'h63 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_508 = _T_252 ? 7'h55 : 7'h0; // @[Mux.scala 27:72]
  wire [5:0] _T_509 = _T_253 ? 6'h21 : 6'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_510 = _T_254 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_511 = _T_255 ? 7'h7d : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _GEN_0 = {{3'd0}, _T_257}; // @[Mux.scala 27:72]
  wire [6:0] _T_512 = _T_256 | _GEN_0; // @[Mux.scala 27:72]
  wire [6:0] _T_513 = _T_512 | _T_258; // @[Mux.scala 27:72]
  wire [7:0] _GEN_1 = {{1'd0}, _T_513}; // @[Mux.scala 27:72]
  wire [7:0] _T_514 = _GEN_1 | _T_259; // @[Mux.scala 27:72]
  wire [7:0] _GEN_2 = {{2'd0}, _T_260}; // @[Mux.scala 27:72]
  wire [7:0] _T_515 = _T_514 | _GEN_2; // @[Mux.scala 27:72]
  wire [7:0] _GEN_3 = {{2'd0}, _T_261}; // @[Mux.scala 27:72]
  wire [7:0] _T_516 = _T_515 | _GEN_3; // @[Mux.scala 27:72]
  wire [7:0] _T_517 = _T_516 | _T_262; // @[Mux.scala 27:72]
  wire [7:0] _GEN_4 = {{2'd0}, _T_263}; // @[Mux.scala 27:72]
  wire [7:0] _T_518 = _T_517 | _GEN_4; // @[Mux.scala 27:72]
  wire [7:0] _T_519 = _T_518 | _T_264; // @[Mux.scala 27:72]
  wire [7:0] _GEN_5 = {{1'd0}, _T_265}; // @[Mux.scala 27:72]
  wire [7:0] _T_520 = _T_519 | _GEN_5; // @[Mux.scala 27:72]
  wire [7:0] _T_521 = _T_520 | _T_266; // @[Mux.scala 27:72]
  wire [7:0] _T_522 = _T_521 | _T_267; // @[Mux.scala 27:72]
  wire [7:0] _T_523 = _T_522 | _T_268; // @[Mux.scala 27:72]
  wire [7:0] _T_524 = _T_523 | _T_269; // @[Mux.scala 27:72]
  wire [7:0] _T_525 = _T_524 | _T_270; // @[Mux.scala 27:72]
  wire [7:0] _T_526 = _T_525 | _T_271; // @[Mux.scala 27:72]
  wire [7:0] _GEN_6 = {{1'd0}, _T_272}; // @[Mux.scala 27:72]
  wire [7:0] _T_527 = _T_526 | _GEN_6; // @[Mux.scala 27:72]
  wire [7:0] _T_528 = _T_527 | _T_273; // @[Mux.scala 27:72]
  wire [7:0] _GEN_7 = {{2'd0}, _T_274}; // @[Mux.scala 27:72]
  wire [7:0] _T_529 = _T_528 | _GEN_7; // @[Mux.scala 27:72]
  wire [7:0] _T_530 = _T_529 | _T_275; // @[Mux.scala 27:72]
  wire [7:0] _T_531 = _T_530 | _T_276; // @[Mux.scala 27:72]
  wire [7:0] _GEN_8 = {{2'd0}, _T_277}; // @[Mux.scala 27:72]
  wire [7:0] _T_532 = _T_531 | _GEN_8; // @[Mux.scala 27:72]
  wire [7:0] _T_533 = _T_532 | _T_278; // @[Mux.scala 27:72]
  wire [7:0] _T_534 = _T_533 | _T_279; // @[Mux.scala 27:72]
  wire [7:0] _GEN_9 = {{2'd0}, _T_280}; // @[Mux.scala 27:72]
  wire [7:0] _T_535 = _T_534 | _GEN_9; // @[Mux.scala 27:72]
  wire [7:0] _T_536 = _T_535 | _T_281; // @[Mux.scala 27:72]
  wire [7:0] _GEN_10 = {{1'd0}, _T_282}; // @[Mux.scala 27:72]
  wire [7:0] _T_537 = _T_536 | _GEN_10; // @[Mux.scala 27:72]
  wire [7:0] _GEN_11 = {{1'd0}, _T_283}; // @[Mux.scala 27:72]
  wire [7:0] _T_538 = _T_537 | _GEN_11; // @[Mux.scala 27:72]
  wire [7:0] _T_539 = _T_538 | _T_284; // @[Mux.scala 27:72]
  wire [7:0] _T_540 = _T_539 | _T_285; // @[Mux.scala 27:72]
  wire [7:0] _T_541 = _T_540 | _T_286; // @[Mux.scala 27:72]
  wire [7:0] _T_542 = _T_541 | _T_287; // @[Mux.scala 27:72]
  wire [7:0] _GEN_12 = {{1'd0}, _T_288}; // @[Mux.scala 27:72]
  wire [7:0] _T_543 = _T_542 | _GEN_12; // @[Mux.scala 27:72]
  wire [7:0] _GEN_13 = {{1'd0}, _T_289}; // @[Mux.scala 27:72]
  wire [7:0] _T_544 = _T_543 | _GEN_13; // @[Mux.scala 27:72]
  wire [7:0] _T_545 = _T_544 | _T_290; // @[Mux.scala 27:72]
  wire [7:0] _GEN_14 = {{2'd0}, _T_291}; // @[Mux.scala 27:72]
  wire [7:0] _T_546 = _T_545 | _GEN_14; // @[Mux.scala 27:72]
  wire [7:0] _T_547 = _T_546 | _T_292; // @[Mux.scala 27:72]
  wire [7:0] _T_548 = _T_547 | _T_293; // @[Mux.scala 27:72]
  wire [7:0] _GEN_15 = {{2'd0}, _T_294}; // @[Mux.scala 27:72]
  wire [7:0] _T_549 = _T_548 | _GEN_15; // @[Mux.scala 27:72]
  wire [7:0] _GEN_16 = {{2'd0}, _T_295}; // @[Mux.scala 27:72]
  wire [7:0] _T_550 = _T_549 | _GEN_16; // @[Mux.scala 27:72]
  wire [7:0] _T_551 = _T_550 | _T_296; // @[Mux.scala 27:72]
  wire [7:0] _GEN_17 = {{1'd0}, _T_297}; // @[Mux.scala 27:72]
  wire [7:0] _T_552 = _T_551 | _GEN_17; // @[Mux.scala 27:72]
  wire [7:0] _T_553 = _T_552 | _T_298; // @[Mux.scala 27:72]
  wire [7:0] _GEN_18 = {{4'd0}, _T_299}; // @[Mux.scala 27:72]
  wire [7:0] _T_554 = _T_553 | _GEN_18; // @[Mux.scala 27:72]
  wire [7:0] _GEN_19 = {{1'd0}, _T_300}; // @[Mux.scala 27:72]
  wire [7:0] _T_555 = _T_554 | _GEN_19; // @[Mux.scala 27:72]
  wire [7:0] _T_556 = _T_555 | _T_301; // @[Mux.scala 27:72]
  wire [7:0] _T_557 = _T_556 | _T_302; // @[Mux.scala 27:72]
  wire [7:0] _GEN_20 = {{1'd0}, _T_303}; // @[Mux.scala 27:72]
  wire [7:0] _T_558 = _T_557 | _GEN_20; // @[Mux.scala 27:72]
  wire [7:0] _GEN_21 = {{4'd0}, _T_304}; // @[Mux.scala 27:72]
  wire [7:0] _T_559 = _T_558 | _GEN_21; // @[Mux.scala 27:72]
  wire [7:0] _GEN_22 = {{2'd0}, _T_305}; // @[Mux.scala 27:72]
  wire [7:0] _T_560 = _T_559 | _GEN_22; // @[Mux.scala 27:72]
  wire [7:0] _T_561 = _T_560 | _T_306; // @[Mux.scala 27:72]
  wire [7:0] _GEN_23 = {{1'd0}, _T_307}; // @[Mux.scala 27:72]
  wire [7:0] _T_562 = _T_561 | _GEN_23; // @[Mux.scala 27:72]
  wire [7:0] _GEN_24 = {{2'd0}, _T_308}; // @[Mux.scala 27:72]
  wire [7:0] _T_563 = _T_562 | _GEN_24; // @[Mux.scala 27:72]
  wire [7:0] _T_564 = _T_563 | _T_309; // @[Mux.scala 27:72]
  wire [7:0] _GEN_25 = {{2'd0}, _T_310}; // @[Mux.scala 27:72]
  wire [7:0] _T_565 = _T_564 | _GEN_25; // @[Mux.scala 27:72]
  wire [7:0] _T_566 = _T_565 | _T_311; // @[Mux.scala 27:72]
  wire [7:0] _GEN_26 = {{1'd0}, _T_312}; // @[Mux.scala 27:72]
  wire [7:0] _T_567 = _T_566 | _GEN_26; // @[Mux.scala 27:72]
  wire [7:0] _GEN_27 = {{1'd0}, _T_313}; // @[Mux.scala 27:72]
  wire [7:0] _T_568 = _T_567 | _GEN_27; // @[Mux.scala 27:72]
  wire [7:0] _T_569 = _T_568 | _T_314; // @[Mux.scala 27:72]
  wire [7:0] _GEN_28 = {{1'd0}, _T_315}; // @[Mux.scala 27:72]
  wire [7:0] _T_570 = _T_569 | _GEN_28; // @[Mux.scala 27:72]
  wire [7:0] _GEN_29 = {{1'd0}, _T_316}; // @[Mux.scala 27:72]
  wire [7:0] _T_571 = _T_570 | _GEN_29; // @[Mux.scala 27:72]
  wire [7:0] _T_572 = _T_571 | _T_317; // @[Mux.scala 27:72]
  wire [7:0] _T_573 = _T_572 | _T_318; // @[Mux.scala 27:72]
  wire [7:0] _GEN_30 = {{2'd0}, _T_319}; // @[Mux.scala 27:72]
  wire [7:0] _T_574 = _T_573 | _GEN_30; // @[Mux.scala 27:72]
  wire [7:0] _GEN_31 = {{1'd0}, _T_320}; // @[Mux.scala 27:72]
  wire [7:0] _T_575 = _T_574 | _GEN_31; // @[Mux.scala 27:72]
  wire [7:0] _T_576 = _T_575 | _T_321; // @[Mux.scala 27:72]
  wire [7:0] _T_577 = _T_576 | _T_322; // @[Mux.scala 27:72]
  wire [7:0] _GEN_32 = {{1'd0}, _T_323}; // @[Mux.scala 27:72]
  wire [7:0] _T_578 = _T_577 | _GEN_32; // @[Mux.scala 27:72]
  wire [7:0] _T_579 = _T_578 | _T_324; // @[Mux.scala 27:72]
  wire [7:0] _GEN_33 = {{1'd0}, _T_325}; // @[Mux.scala 27:72]
  wire [7:0] _T_580 = _T_579 | _GEN_33; // @[Mux.scala 27:72]
  wire [7:0] _T_581 = _T_580 | _T_326; // @[Mux.scala 27:72]
  wire [7:0] _GEN_34 = {{3'd0}, _T_327}; // @[Mux.scala 27:72]
  wire [7:0] _T_582 = _T_581 | _GEN_34; // @[Mux.scala 27:72]
  wire [7:0] _T_583 = _T_582 | _T_328; // @[Mux.scala 27:72]
  wire [7:0] _T_584 = _T_583 | _T_329; // @[Mux.scala 27:72]
  wire [7:0] _GEN_35 = {{1'd0}, _T_330}; // @[Mux.scala 27:72]
  wire [7:0] _T_585 = _T_584 | _GEN_35; // @[Mux.scala 27:72]
  wire [7:0] _T_586 = _T_585 | _T_331; // @[Mux.scala 27:72]
  wire [7:0] _GEN_36 = {{1'd0}, _T_332}; // @[Mux.scala 27:72]
  wire [7:0] _T_587 = _T_586 | _GEN_36; // @[Mux.scala 27:72]
  wire [7:0] _GEN_37 = {{1'd0}, _T_333}; // @[Mux.scala 27:72]
  wire [7:0] _T_588 = _T_587 | _GEN_37; // @[Mux.scala 27:72]
  wire [7:0] _T_589 = _T_588 | _T_334; // @[Mux.scala 27:72]
  wire [7:0] _T_590 = _T_589 | _T_335; // @[Mux.scala 27:72]
  wire [7:0] _GEN_38 = {{1'd0}, _T_336}; // @[Mux.scala 27:72]
  wire [7:0] _T_591 = _T_590 | _GEN_38; // @[Mux.scala 27:72]
  wire [7:0] _GEN_39 = {{1'd0}, _T_337}; // @[Mux.scala 27:72]
  wire [7:0] _T_592 = _T_591 | _GEN_39; // @[Mux.scala 27:72]
  wire [7:0] _GEN_40 = {{1'd0}, _T_338}; // @[Mux.scala 27:72]
  wire [7:0] _T_593 = _T_592 | _GEN_40; // @[Mux.scala 27:72]
  wire [7:0] _GEN_41 = {{1'd0}, _T_339}; // @[Mux.scala 27:72]
  wire [7:0] _T_594 = _T_593 | _GEN_41; // @[Mux.scala 27:72]
  wire [7:0] _T_595 = _T_594 | _T_340; // @[Mux.scala 27:72]
  wire [7:0] _T_596 = _T_595 | _T_341; // @[Mux.scala 27:72]
  wire [7:0] _T_597 = _T_596 | _T_342; // @[Mux.scala 27:72]
  wire [7:0] _T_598 = _T_597 | _T_343; // @[Mux.scala 27:72]
  wire [7:0] _GEN_42 = {{1'd0}, _T_344}; // @[Mux.scala 27:72]
  wire [7:0] _T_599 = _T_598 | _GEN_42; // @[Mux.scala 27:72]
  wire [7:0] _GEN_43 = {{3'd0}, _T_345}; // @[Mux.scala 27:72]
  wire [7:0] _T_600 = _T_599 | _GEN_43; // @[Mux.scala 27:72]
  wire [7:0] _GEN_44 = {{1'd0}, _T_346}; // @[Mux.scala 27:72]
  wire [7:0] _T_601 = _T_600 | _GEN_44; // @[Mux.scala 27:72]
  wire [7:0] _GEN_45 = {{1'd0}, _T_347}; // @[Mux.scala 27:72]
  wire [7:0] _T_602 = _T_601 | _GEN_45; // @[Mux.scala 27:72]
  wire [7:0] _T_603 = _T_602 | _T_348; // @[Mux.scala 27:72]
  wire [7:0] _T_604 = _T_603 | _T_349; // @[Mux.scala 27:72]
  wire [7:0] _T_605 = _T_604 | _T_350; // @[Mux.scala 27:72]
  wire [7:0] _T_606 = _T_605 | _T_351; // @[Mux.scala 27:72]
  wire [7:0] _T_607 = _T_606 | _T_352; // @[Mux.scala 27:72]
  wire [7:0] _T_608 = _T_607 | _T_353; // @[Mux.scala 27:72]
  wire [7:0] _T_609 = _T_608 | _T_354; // @[Mux.scala 27:72]
  wire [7:0] _T_611 = _T_609 | _T_356; // @[Mux.scala 27:72]
  wire [7:0] _T_612 = _T_611 | _T_357; // @[Mux.scala 27:72]
  wire [7:0] _T_613 = _T_612 | _T_358; // @[Mux.scala 27:72]
  wire [7:0] _GEN_46 = {{4'd0}, _T_359}; // @[Mux.scala 27:72]
  wire [7:0] _T_614 = _T_613 | _GEN_46; // @[Mux.scala 27:72]
  wire [7:0] _T_615 = _T_614 | _T_360; // @[Mux.scala 27:72]
  wire [7:0] _T_616 = _T_615 | _T_361; // @[Mux.scala 27:72]
  wire [7:0] _GEN_47 = {{1'd0}, _T_362}; // @[Mux.scala 27:72]
  wire [7:0] _T_617 = _T_616 | _GEN_47; // @[Mux.scala 27:72]
  wire [7:0] _GEN_48 = {{5'd0}, _T_363}; // @[Mux.scala 27:72]
  wire [7:0] _T_618 = _T_617 | _GEN_48; // @[Mux.scala 27:72]
  wire [7:0] _T_619 = _T_618 | _T_364; // @[Mux.scala 27:72]
  wire [7:0] _T_620 = _T_619 | _T_365; // @[Mux.scala 27:72]
  wire [7:0] _GEN_49 = {{1'd0}, _T_366}; // @[Mux.scala 27:72]
  wire [7:0] _T_621 = _T_620 | _GEN_49; // @[Mux.scala 27:72]
  wire [7:0] _GEN_50 = {{5'd0}, _T_367}; // @[Mux.scala 27:72]
  wire [7:0] _T_622 = _T_621 | _GEN_50; // @[Mux.scala 27:72]
  wire [7:0] _T_623 = _T_622 | _T_368; // @[Mux.scala 27:72]
  wire [7:0] _GEN_51 = {{2'd0}, _T_369}; // @[Mux.scala 27:72]
  wire [7:0] _T_624 = _T_623 | _GEN_51; // @[Mux.scala 27:72]
  wire [7:0] _GEN_52 = {{3'd0}, _T_370}; // @[Mux.scala 27:72]
  wire [7:0] _T_625 = _T_624 | _GEN_52; // @[Mux.scala 27:72]
  wire [7:0] _T_626 = _T_625 | _T_371; // @[Mux.scala 27:72]
  wire [7:0] _T_627 = _T_626 | _T_372; // @[Mux.scala 27:72]
  wire [7:0] _GEN_53 = {{2'd0}, _T_373}; // @[Mux.scala 27:72]
  wire [7:0] _T_628 = _T_627 | _GEN_53; // @[Mux.scala 27:72]
  wire [7:0] _GEN_54 = {{4'd0}, _T_374}; // @[Mux.scala 27:72]
  wire [7:0] _T_629 = _T_628 | _GEN_54; // @[Mux.scala 27:72]
  wire [7:0] _GEN_55 = {{6'd0}, _T_375}; // @[Mux.scala 27:72]
  wire [7:0] _T_630 = _T_629 | _GEN_55; // @[Mux.scala 27:72]
  wire [7:0] _T_631 = _T_630 | _T_376; // @[Mux.scala 27:72]
  wire [7:0] _T_632 = _T_631 | _T_377; // @[Mux.scala 27:72]
  wire [7:0] _T_633 = _T_632 | _T_378; // @[Mux.scala 27:72]
  wire [7:0] _GEN_56 = {{6'd0}, _T_379}; // @[Mux.scala 27:72]
  wire [7:0] _T_634 = _T_633 | _GEN_56; // @[Mux.scala 27:72]
  wire [7:0] _GEN_57 = {{7'd0}, _T_124}; // @[Mux.scala 27:72]
  wire [7:0] _T_635 = _T_634 | _GEN_57; // @[Mux.scala 27:72]
  wire [7:0] _GEN_58 = {{3'd0}, _T_381}; // @[Mux.scala 27:72]
  wire [7:0] _T_636 = _T_635 | _GEN_58; // @[Mux.scala 27:72]
  wire [7:0] _T_637 = _T_636 | _T_382; // @[Mux.scala 27:72]
  wire [7:0] _GEN_59 = {{1'd0}, _T_383}; // @[Mux.scala 27:72]
  wire [7:0] _T_638 = _T_637 | _GEN_59; // @[Mux.scala 27:72]
  wire [7:0] _GEN_60 = {{2'd0}, _T_384}; // @[Mux.scala 27:72]
  wire [7:0] _T_639 = _T_638 | _GEN_60; // @[Mux.scala 27:72]
  wire [7:0] _T_640 = _T_639 | _T_385; // @[Mux.scala 27:72]
  wire [7:0] _GEN_61 = {{3'd0}, _T_386}; // @[Mux.scala 27:72]
  wire [7:0] _T_641 = _T_640 | _GEN_61; // @[Mux.scala 27:72]
  wire [7:0] _GEN_62 = {{1'd0}, _T_387}; // @[Mux.scala 27:72]
  wire [7:0] _T_642 = _T_641 | _GEN_62; // @[Mux.scala 27:72]
  wire [7:0] _GEN_63 = {{1'd0}, _T_388}; // @[Mux.scala 27:72]
  wire [7:0] _T_643 = _T_642 | _GEN_63; // @[Mux.scala 27:72]
  wire [7:0] _GEN_64 = {{1'd0}, _T_389}; // @[Mux.scala 27:72]
  wire [7:0] _T_644 = _T_643 | _GEN_64; // @[Mux.scala 27:72]
  wire [7:0] _T_645 = _T_644 | _T_390; // @[Mux.scala 27:72]
  wire [7:0] _T_646 = _T_645 | _T_391; // @[Mux.scala 27:72]
  wire [7:0] _T_647 = _T_646 | _T_392; // @[Mux.scala 27:72]
  wire [7:0] _T_648 = _T_647 | _T_393; // @[Mux.scala 27:72]
  wire [7:0] _T_649 = _T_648 | _T_394; // @[Mux.scala 27:72]
  wire [7:0] _T_650 = _T_649 | _T_395; // @[Mux.scala 27:72]
  wire [7:0] _T_651 = _T_650 | _T_396; // @[Mux.scala 27:72]
  wire [7:0] _T_652 = _T_651 | _T_397; // @[Mux.scala 27:72]
  wire [7:0] _T_653 = _T_652 | _T_398; // @[Mux.scala 27:72]
  wire [7:0] _GEN_65 = {{1'd0}, _T_399}; // @[Mux.scala 27:72]
  wire [7:0] _T_654 = _T_653 | _GEN_65; // @[Mux.scala 27:72]
  wire [7:0] _T_655 = _T_654 | _T_400; // @[Mux.scala 27:72]
  wire [7:0] _T_656 = _T_655 | _T_401; // @[Mux.scala 27:72]
  wire [7:0] _GEN_66 = {{1'd0}, _T_402}; // @[Mux.scala 27:72]
  wire [7:0] _T_657 = _T_656 | _GEN_66; // @[Mux.scala 27:72]
  wire [7:0] _GEN_67 = {{2'd0}, _T_403}; // @[Mux.scala 27:72]
  wire [7:0] _T_658 = _T_657 | _GEN_67; // @[Mux.scala 27:72]
  wire [7:0] _T_659 = _T_658 | _T_404; // @[Mux.scala 27:72]
  wire [7:0] _T_660 = _T_659 | _T_405; // @[Mux.scala 27:72]
  wire [7:0] _GEN_68 = {{2'd0}, _T_406}; // @[Mux.scala 27:72]
  wire [7:0] _T_661 = _T_660 | _GEN_68; // @[Mux.scala 27:72]
  wire [7:0] _T_662 = _T_661 | _T_407; // @[Mux.scala 27:72]
  wire [7:0] _T_663 = _T_662 | _T_408; // @[Mux.scala 27:72]
  wire [7:0] _T_664 = _T_663 | _T_409; // @[Mux.scala 27:72]
  wire [7:0] _GEN_69 = {{2'd0}, _T_410}; // @[Mux.scala 27:72]
  wire [7:0] _T_665 = _T_664 | _GEN_69; // @[Mux.scala 27:72]
  wire [7:0] _T_666 = _T_665 | _T_411; // @[Mux.scala 27:72]
  wire [7:0] _GEN_70 = {{3'd0}, _T_412}; // @[Mux.scala 27:72]
  wire [7:0] _T_667 = _T_666 | _GEN_70; // @[Mux.scala 27:72]
  wire [7:0] _GEN_71 = {{1'd0}, _T_413}; // @[Mux.scala 27:72]
  wire [7:0] _T_668 = _T_667 | _GEN_71; // @[Mux.scala 27:72]
  wire [7:0] _T_669 = _T_668 | _T_414; // @[Mux.scala 27:72]
  wire [7:0] _GEN_72 = {{1'd0}, _T_415}; // @[Mux.scala 27:72]
  wire [7:0] _T_670 = _T_669 | _GEN_72; // @[Mux.scala 27:72]
  wire [7:0] _GEN_73 = {{1'd0}, _T_416}; // @[Mux.scala 27:72]
  wire [7:0] _T_671 = _T_670 | _GEN_73; // @[Mux.scala 27:72]
  wire [7:0] _T_672 = _T_671 | _T_417; // @[Mux.scala 27:72]
  wire [7:0] _GEN_74 = {{3'd0}, _T_418}; // @[Mux.scala 27:72]
  wire [7:0] _T_673 = _T_672 | _GEN_74; // @[Mux.scala 27:72]
  wire [7:0] _GEN_75 = {{1'd0}, _T_419}; // @[Mux.scala 27:72]
  wire [7:0] _T_674 = _T_673 | _GEN_75; // @[Mux.scala 27:72]
  wire [7:0] _GEN_76 = {{3'd0}, _T_420}; // @[Mux.scala 27:72]
  wire [7:0] _T_675 = _T_674 | _GEN_76; // @[Mux.scala 27:72]
  wire [7:0] _GEN_77 = {{2'd0}, _T_421}; // @[Mux.scala 27:72]
  wire [7:0] _T_676 = _T_675 | _GEN_77; // @[Mux.scala 27:72]
  wire [7:0] _T_677 = _T_676 | _T_422; // @[Mux.scala 27:72]
  wire [7:0] _T_678 = _T_677 | _T_423; // @[Mux.scala 27:72]
  wire [7:0] _GEN_78 = {{1'd0}, _T_424}; // @[Mux.scala 27:72]
  wire [7:0] _T_679 = _T_678 | _GEN_78; // @[Mux.scala 27:72]
  wire [7:0] _T_680 = _T_679 | _T_425; // @[Mux.scala 27:72]
  wire [7:0] _GEN_79 = {{1'd0}, _T_426}; // @[Mux.scala 27:72]
  wire [7:0] _T_681 = _T_680 | _GEN_79; // @[Mux.scala 27:72]
  wire [7:0] _GEN_80 = {{4'd0}, _T_427}; // @[Mux.scala 27:72]
  wire [7:0] _T_682 = _T_681 | _GEN_80; // @[Mux.scala 27:72]
  wire [7:0] _T_683 = _T_682 | _T_428; // @[Mux.scala 27:72]
  wire [7:0] _GEN_81 = {{3'd0}, _T_429}; // @[Mux.scala 27:72]
  wire [7:0] _T_684 = _T_683 | _GEN_81; // @[Mux.scala 27:72]
  wire [7:0] _T_685 = _T_684 | _T_430; // @[Mux.scala 27:72]
  wire [7:0] _GEN_82 = {{3'd0}, _T_431}; // @[Mux.scala 27:72]
  wire [7:0] _T_686 = _T_685 | _GEN_82; // @[Mux.scala 27:72]
  wire [7:0] _T_687 = _T_686 | _T_432; // @[Mux.scala 27:72]
  wire [7:0] _GEN_83 = {{1'd0}, _T_433}; // @[Mux.scala 27:72]
  wire [7:0] _T_688 = _T_687 | _GEN_83; // @[Mux.scala 27:72]
  wire [7:0] _GEN_84 = {{2'd0}, _T_434}; // @[Mux.scala 27:72]
  wire [7:0] _T_689 = _T_688 | _GEN_84; // @[Mux.scala 27:72]
  wire [7:0] _GEN_85 = {{1'd0}, _T_435}; // @[Mux.scala 27:72]
  wire [7:0] _T_690 = _T_689 | _GEN_85; // @[Mux.scala 27:72]
  wire [7:0] _T_691 = _T_690 | _T_436; // @[Mux.scala 27:72]
  wire [7:0] _T_692 = _T_691 | _T_437; // @[Mux.scala 27:72]
  wire [7:0] _GEN_86 = {{1'd0}, _T_438}; // @[Mux.scala 27:72]
  wire [7:0] _T_693 = _T_692 | _GEN_86; // @[Mux.scala 27:72]
  wire [7:0] _GEN_87 = {{2'd0}, _T_439}; // @[Mux.scala 27:72]
  wire [7:0] _T_694 = _T_693 | _GEN_87; // @[Mux.scala 27:72]
  wire [7:0] _T_695 = _T_694 | _T_440; // @[Mux.scala 27:72]
  wire [7:0] _T_696 = _T_695 | _T_441; // @[Mux.scala 27:72]
  wire [7:0] _T_697 = _T_696 | _T_442; // @[Mux.scala 27:72]
  wire [7:0] _T_698 = _T_697 | _T_443; // @[Mux.scala 27:72]
  wire [7:0] _GEN_88 = {{1'd0}, _T_444}; // @[Mux.scala 27:72]
  wire [7:0] _T_699 = _T_698 | _GEN_88; // @[Mux.scala 27:72]
  wire [7:0] _T_700 = _T_699 | _T_445; // @[Mux.scala 27:72]
  wire [7:0] _GEN_89 = {{1'd0}, _T_446}; // @[Mux.scala 27:72]
  wire [7:0] _T_701 = _T_700 | _GEN_89; // @[Mux.scala 27:72]
  wire [7:0] _T_702 = _T_701 | _T_447; // @[Mux.scala 27:72]
  wire [7:0] _GEN_90 = {{3'd0}, _T_448}; // @[Mux.scala 27:72]
  wire [7:0] _T_703 = _T_702 | _GEN_90; // @[Mux.scala 27:72]
  wire [7:0] _T_704 = _T_703 | _T_449; // @[Mux.scala 27:72]
  wire [7:0] _T_705 = _T_704 | _T_450; // @[Mux.scala 27:72]
  wire [7:0] _GEN_91 = {{2'd0}, _T_451}; // @[Mux.scala 27:72]
  wire [7:0] _T_706 = _T_705 | _GEN_91; // @[Mux.scala 27:72]
  wire [7:0] _T_707 = _T_706 | _T_452; // @[Mux.scala 27:72]
  wire [7:0] _GEN_92 = {{5'd0}, _T_453}; // @[Mux.scala 27:72]
  wire [7:0] _T_708 = _T_707 | _GEN_92; // @[Mux.scala 27:72]
  wire [7:0] _T_709 = _T_708 | _T_454; // @[Mux.scala 27:72]
  wire [7:0] _GEN_93 = {{2'd0}, _T_455}; // @[Mux.scala 27:72]
  wire [7:0] _T_710 = _T_709 | _GEN_93; // @[Mux.scala 27:72]
  wire [7:0] _T_711 = _T_710 | _T_456; // @[Mux.scala 27:72]
  wire [7:0] _GEN_94 = {{3'd0}, _T_457}; // @[Mux.scala 27:72]
  wire [7:0] _T_712 = _T_711 | _GEN_94; // @[Mux.scala 27:72]
  wire [7:0] _GEN_95 = {{3'd0}, _T_458}; // @[Mux.scala 27:72]
  wire [7:0] _T_713 = _T_712 | _GEN_95; // @[Mux.scala 27:72]
  wire [7:0] _GEN_96 = {{1'd0}, _T_459}; // @[Mux.scala 27:72]
  wire [7:0] _T_714 = _T_713 | _GEN_96; // @[Mux.scala 27:72]
  wire [7:0] _GEN_97 = {{2'd0}, _T_460}; // @[Mux.scala 27:72]
  wire [7:0] _T_715 = _T_714 | _GEN_97; // @[Mux.scala 27:72]
  wire [7:0] _T_716 = _T_715 | _T_461; // @[Mux.scala 27:72]
  wire [7:0] _T_717 = _T_716 | _T_462; // @[Mux.scala 27:72]
  wire [7:0] _GEN_98 = {{1'd0}, _T_463}; // @[Mux.scala 27:72]
  wire [7:0] _T_718 = _T_717 | _GEN_98; // @[Mux.scala 27:72]
  wire [7:0] _GEN_99 = {{1'd0}, _T_464}; // @[Mux.scala 27:72]
  wire [7:0] _T_719 = _T_718 | _GEN_99; // @[Mux.scala 27:72]
  wire [7:0] _GEN_100 = {{1'd0}, _T_465}; // @[Mux.scala 27:72]
  wire [7:0] _T_720 = _T_719 | _GEN_100; // @[Mux.scala 27:72]
  wire [7:0] _GEN_101 = {{1'd0}, _T_466}; // @[Mux.scala 27:72]
  wire [7:0] _T_721 = _T_720 | _GEN_101; // @[Mux.scala 27:72]
  wire [7:0] _T_722 = _T_721 | _T_467; // @[Mux.scala 27:72]
  wire [7:0] _GEN_102 = {{3'd0}, _T_468}; // @[Mux.scala 27:72]
  wire [7:0] _T_723 = _T_722 | _GEN_102; // @[Mux.scala 27:72]
  wire [7:0] _T_724 = _T_723 | _T_469; // @[Mux.scala 27:72]
  wire [7:0] _GEN_103 = {{1'd0}, _T_470}; // @[Mux.scala 27:72]
  wire [7:0] _T_725 = _T_724 | _GEN_103; // @[Mux.scala 27:72]
  wire [7:0] _GEN_104 = {{4'd0}, _T_471}; // @[Mux.scala 27:72]
  wire [7:0] _T_726 = _T_725 | _GEN_104; // @[Mux.scala 27:72]
  wire [7:0] _GEN_105 = {{2'd0}, _T_472}; // @[Mux.scala 27:72]
  wire [7:0] _T_727 = _T_726 | _GEN_105; // @[Mux.scala 27:72]
  wire [7:0] _T_728 = _T_727 | _T_473; // @[Mux.scala 27:72]
  wire [7:0] _GEN_106 = {{1'd0}, _T_474}; // @[Mux.scala 27:72]
  wire [7:0] _T_729 = _T_728 | _GEN_106; // @[Mux.scala 27:72]
  wire [7:0] _T_730 = _T_729 | _T_475; // @[Mux.scala 27:72]
  wire [7:0] _T_731 = _T_730 | _T_476; // @[Mux.scala 27:72]
  wire [7:0] _T_732 = _T_731 | _T_477; // @[Mux.scala 27:72]
  wire [7:0] _T_733 = _T_732 | _T_478; // @[Mux.scala 27:72]
  wire [7:0] _T_734 = _T_733 | _T_479; // @[Mux.scala 27:72]
  wire [7:0] _T_735 = _T_734 | _T_480; // @[Mux.scala 27:72]
  wire [7:0] _T_736 = _T_735 | _T_481; // @[Mux.scala 27:72]
  wire [7:0] _GEN_107 = {{2'd0}, _T_482}; // @[Mux.scala 27:72]
  wire [7:0] _T_737 = _T_736 | _GEN_107; // @[Mux.scala 27:72]
  wire [7:0] _GEN_108 = {{1'd0}, _T_483}; // @[Mux.scala 27:72]
  wire [7:0] _T_738 = _T_737 | _GEN_108; // @[Mux.scala 27:72]
  wire [7:0] _T_739 = _T_738 | _T_484; // @[Mux.scala 27:72]
  wire [7:0] _GEN_109 = {{2'd0}, _T_485}; // @[Mux.scala 27:72]
  wire [7:0] _T_740 = _T_739 | _GEN_109; // @[Mux.scala 27:72]
  wire [7:0] _T_741 = _T_740 | _T_486; // @[Mux.scala 27:72]
  wire [7:0] _T_742 = _T_741 | _T_487; // @[Mux.scala 27:72]
  wire [7:0] _T_743 = _T_742 | _T_488; // @[Mux.scala 27:72]
  wire [7:0] _T_744 = _T_743 | _T_489; // @[Mux.scala 27:72]
  wire [7:0] _T_745 = _T_744 | _T_490; // @[Mux.scala 27:72]
  wire [7:0] _GEN_110 = {{2'd0}, _T_491}; // @[Mux.scala 27:72]
  wire [7:0] _T_746 = _T_745 | _GEN_110; // @[Mux.scala 27:72]
  wire [7:0] _T_747 = _T_746 | _T_492; // @[Mux.scala 27:72]
  wire [7:0] _GEN_111 = {{1'd0}, _T_493}; // @[Mux.scala 27:72]
  wire [7:0] _T_748 = _T_747 | _GEN_111; // @[Mux.scala 27:72]
  wire [7:0] _T_749 = _T_748 | _T_494; // @[Mux.scala 27:72]
  wire [7:0] _GEN_112 = {{1'd0}, _T_495}; // @[Mux.scala 27:72]
  wire [7:0] _T_750 = _T_749 | _GEN_112; // @[Mux.scala 27:72]
  wire [7:0] _GEN_113 = {{3'd0}, _T_496}; // @[Mux.scala 27:72]
  wire [7:0] _T_751 = _T_750 | _GEN_113; // @[Mux.scala 27:72]
  wire [7:0] _GEN_114 = {{2'd0}, _T_497}; // @[Mux.scala 27:72]
  wire [7:0] _T_752 = _T_751 | _GEN_114; // @[Mux.scala 27:72]
  wire [7:0] _GEN_115 = {{5'd0}, _T_498}; // @[Mux.scala 27:72]
  wire [7:0] _T_753 = _T_752 | _GEN_115; // @[Mux.scala 27:72]
  wire [7:0] _GEN_116 = {{1'd0}, _T_499}; // @[Mux.scala 27:72]
  wire [7:0] _T_754 = _T_753 | _GEN_116; // @[Mux.scala 27:72]
  wire [7:0] _T_755 = _T_754 | _T_500; // @[Mux.scala 27:72]
  wire [7:0] _GEN_117 = {{1'd0}, _T_501}; // @[Mux.scala 27:72]
  wire [7:0] _T_756 = _T_755 | _GEN_117; // @[Mux.scala 27:72]
  wire [7:0] _T_757 = _T_756 | _T_502; // @[Mux.scala 27:72]
  wire [7:0] _GEN_118 = {{2'd0}, _T_503}; // @[Mux.scala 27:72]
  wire [7:0] _T_758 = _T_757 | _GEN_118; // @[Mux.scala 27:72]
  wire [7:0] _T_759 = _T_758 | _T_504; // @[Mux.scala 27:72]
  wire [7:0] _GEN_119 = {{1'd0}, _T_505}; // @[Mux.scala 27:72]
  wire [7:0] _T_760 = _T_759 | _GEN_119; // @[Mux.scala 27:72]
  wire [7:0] _GEN_120 = {{3'd0}, _T_506}; // @[Mux.scala 27:72]
  wire [7:0] _T_761 = _T_760 | _GEN_120; // @[Mux.scala 27:72]
  wire [7:0] _GEN_121 = {{1'd0}, _T_507}; // @[Mux.scala 27:72]
  wire [7:0] _T_762 = _T_761 | _GEN_121; // @[Mux.scala 27:72]
  wire [7:0] _GEN_122 = {{1'd0}, _T_508}; // @[Mux.scala 27:72]
  wire [7:0] _T_763 = _T_762 | _GEN_122; // @[Mux.scala 27:72]
  wire [7:0] _GEN_123 = {{2'd0}, _T_509}; // @[Mux.scala 27:72]
  wire [7:0] _T_764 = _T_763 | _GEN_123; // @[Mux.scala 27:72]
  wire [7:0] _GEN_124 = {{4'd0}, _T_510}; // @[Mux.scala 27:72]
  wire [7:0] _T_765 = _T_764 | _GEN_124; // @[Mux.scala 27:72]
  wire [7:0] _GEN_125 = {{1'd0}, _T_511}; // @[Mux.scala 27:72]
  assign io_byte_out = _T_765 | _GEN_125; // @[cipher.scala 63:15]
endmodule
