module el2_ifu_compress_ctl(
  input         clock,
  input         reset,
  input  [31:0] io_din,
  output [31:0] io_dout
);
  wire  _T_1 = io_din[1:0] != 2'h3; // @[el2_ifu_compress_ctl.scala 401:27]
  wire  _T_3 = |io_din[12:5]; // @[el2_ifu_compress_ctl.scala 257:29]
  wire [6:0] _T_4 = _T_3 ? 7'h13 : 7'h1f; // @[el2_ifu_compress_ctl.scala 257:20]
  wire [29:0] _T_18 = {io_din[10:7],io_din[12:11],io_din[5],io_din[6],2'h0,5'h2,3'h0,2'h1,io_din[4:2],_T_4}; // @[Cat.scala 29:58]
  wire [7:0] _T_28 = {io_din[6:5],io_din[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_36 = {io_din[6:5],io_din[12:10],3'h0,2'h1,io_din[9:7],3'h3,2'h1,io_din[4:2],7'h7}; // @[Cat.scala 29:58]
  wire [6:0] _T_50 = {io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [26:0] _T_58 = {io_din[5],io_din[12:10],io_din[6],2'h0,2'h1,io_din[9:7],3'h2,2'h1,io_din[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [26:0] _T_80 = {io_din[5],io_din[12:10],io_din[6],2'h0,2'h1,io_din[9:7],3'h2,2'h1,io_din[4:2],7'h7}; // @[Cat.scala 29:58]
  wire [26:0] _T_111 = {_T_50[6:5],2'h1,io_din[4:2],2'h1,io_din[9:7],3'h2,_T_50[4:0],7'h3f}; // @[Cat.scala 29:58]
  wire [27:0] _T_138 = {_T_28[7:5],2'h1,io_din[4:2],2'h1,io_din[9:7],3'h3,_T_28[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [26:0] _T_169 = {_T_50[6:5],2'h1,io_din[4:2],2'h1,io_din[9:7],3'h2,_T_50[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [26:0] _T_200 = {_T_50[6:5],2'h1,io_din[4:2],2'h1,io_din[9:7],3'h2,_T_50[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [6:0] _T_211 = io_din[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_213 = {_T_211,io_din[6:2]}; // @[Cat.scala 29:58]
  wire [31:0] _T_219 = {_T_211,io_din[6:2],io_din[11:7],3'h0,io_din[11:7],7'h13}; // @[Cat.scala 29:58]
  wire [9:0] _T_228 = io_din[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  wire [20:0] _T_243 = {_T_228,io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_306 = {_T_243[20],_T_243[10:1],_T_243[11],_T_243[19:12],5'h1,7'h6f}; // @[Cat.scala 29:58]
  wire [31:0] _T_321 = {_T_211,io_din[6:2],5'h0,3'h0,io_din[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_332 = |_T_213; // @[el2_ifu_compress_ctl.scala 294:29]
  wire [6:0] _T_333 = _T_332 ? 7'h37 : 7'h3f; // @[el2_ifu_compress_ctl.scala 294:20]
  wire [14:0] _T_336 = io_din[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_339 = {_T_336,io_din[6:2],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_343 = {_T_339[31:12],io_din[11:7],_T_333}; // @[Cat.scala 29:58]
  wire  _T_351 = io_din[11:7] == 5'h0; // @[el2_ifu_compress_ctl.scala 296:14]
  wire  _T_353 = io_din[11:7] == 5'h2; // @[el2_ifu_compress_ctl.scala 296:27]
  wire  _T_354 = _T_351 | _T_353; // @[el2_ifu_compress_ctl.scala 296:21]
  wire [6:0] _T_361 = _T_332 ? 7'h13 : 7'h1f; // @[el2_ifu_compress_ctl.scala 290:20]
  wire [2:0] _T_364 = io_din[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_379 = {_T_364,io_din[4:3],io_din[5],io_din[2],io_din[6],4'h0,io_din[11:7],3'h0,io_din[11:7],_T_361}; // @[Cat.scala 29:58]
  wire [31:0] _T_386_bits = _T_354 ? _T_379 : _T_343; // @[el2_ifu_compress_ctl.scala 296:10]
  wire [25:0] _T_397 = {io_din[12],io_din[6:2],2'h1,io_din[9:7],3'h5,2'h1,io_din[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_172 = {{5'd0}, _T_397}; // @[el2_ifu_compress_ctl.scala 303:23]
  wire [30:0] _T_409 = _GEN_172 | 31'h40000000; // @[el2_ifu_compress_ctl.scala 303:23]
  wire [31:0] _T_422 = {_T_211,io_din[6:2],2'h1,io_din[9:7],3'h7,2'h1,io_din[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [2:0] _T_426 = {io_din[12],io_din[6:5]}; // @[Cat.scala 29:58]
  wire  _T_428 = io_din[6:5] == 2'h0; // @[el2_ifu_compress_ctl.scala 307:30]
  wire [30:0] _T_429 = _T_428 ? 31'h40000000 : 31'h0; // @[el2_ifu_compress_ctl.scala 307:22]
  wire [6:0] _T_431 = io_din[12] ? 7'h3b : 7'h33; // @[el2_ifu_compress_ctl.scala 308:22]
  wire [2:0] _GEN_1 = 3'h1 == _T_426 ? 3'h4 : 3'h0; // @[Cat.scala 29:58]
  wire [2:0] _GEN_2 = 3'h2 == _T_426 ? 3'h6 : _GEN_1; // @[Cat.scala 29:58]
  wire [2:0] _GEN_3 = 3'h3 == _T_426 ? 3'h7 : _GEN_2; // @[Cat.scala 29:58]
  wire [2:0] _GEN_4 = 3'h4 == _T_426 ? 3'h0 : _GEN_3; // @[Cat.scala 29:58]
  wire [2:0] _GEN_5 = 3'h5 == _T_426 ? 3'h0 : _GEN_4; // @[Cat.scala 29:58]
  wire [2:0] _GEN_6 = 3'h6 == _T_426 ? 3'h2 : _GEN_5; // @[Cat.scala 29:58]
  wire [2:0] _GEN_7 = 3'h7 == _T_426 ? 3'h3 : _GEN_6; // @[Cat.scala 29:58]
  wire [24:0] _T_441 = {2'h1,io_din[4:2],2'h1,io_din[9:7],_GEN_7,2'h1,io_din[9:7],_T_431}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_173 = {{6'd0}, _T_441}; // @[el2_ifu_compress_ctl.scala 309:43]
  wire [30:0] _T_442 = _GEN_173 | _T_429; // @[el2_ifu_compress_ctl.scala 309:43]
  wire [31:0] _T_443_0 = {{6'd0}, _T_397}; // @[el2_ifu_compress_ctl.scala 311:19 el2_ifu_compress_ctl.scala 311:19]
  wire [31:0] _T_443_1 = {{1'd0}, _T_409}; // @[el2_ifu_compress_ctl.scala 311:19 el2_ifu_compress_ctl.scala 311:19]
  wire [31:0] _GEN_9 = 2'h1 == io_din[11:10] ? _T_443_1 : _T_443_0; // @[el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_10 = 2'h2 == io_din[11:10] ? _T_422 : _GEN_9; // @[el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_443_3 = {{1'd0}, _T_442}; // @[el2_ifu_compress_ctl.scala 311:19 el2_ifu_compress_ctl.scala 311:19]
  wire [31:0] _GEN_11 = 2'h3 == io_din[11:10] ? _T_443_3 : _GEN_10; // @[el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_533 = {_T_243[20],_T_243[10:1],_T_243[11],_T_243[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58]
  wire [4:0] _T_542 = io_din[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [12:0] _T_551 = {_T_542,io_din[6:5],io_din[2],io_din[11:10],io_din[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_600 = {_T_551[12],_T_551[10:5],5'h0,2'h1,io_din[9:7],3'h0,_T_551[4:1],_T_551[11],7'h63}; // @[Cat.scala 29:58]
  wire [31:0] _T_667 = {_T_551[12],_T_551[10:5],5'h0,2'h1,io_din[9:7],3'h1,_T_551[4:1],_T_551[11],7'h63}; // @[Cat.scala 29:58]
  wire  _T_673 = |io_din[11:7]; // @[el2_ifu_compress_ctl.scala 317:27]
  wire [6:0] _T_674 = _T_673 ? 7'h3 : 7'h1f; // @[el2_ifu_compress_ctl.scala 317:23]
  wire [25:0] _T_683 = {io_din[12],io_din[6:2],io_din[11:7],3'h1,io_din[11:7],7'h13}; // @[Cat.scala 29:58]
  wire [28:0] _T_699 = {io_din[4:2],io_din[12],io_din[6:5],3'h0,5'h2,3'h3,io_din[11:7],7'h7}; // @[Cat.scala 29:58]
  wire [27:0] _T_714 = {io_din[3:2],io_din[12],io_din[6:4],2'h0,5'h2,3'h2,io_din[11:7],_T_674}; // @[Cat.scala 29:58]
  wire [27:0] _T_729 = {io_din[3:2],io_din[12],io_din[6:4],2'h0,5'h2,3'h2,io_din[11:7],7'h7}; // @[Cat.scala 29:58]
  wire [24:0] _T_739 = {io_din[6:2],5'h0,3'h0,io_din[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_750 = {io_din[6:2],io_din[11:7],3'h0,io_din[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_761 = {io_din[6:2],io_din[11:7],3'h0,12'h67}; // @[Cat.scala 29:58]
  wire [24:0] _T_763 = {_T_761[24:7],7'h1f}; // @[Cat.scala 29:58]
  wire [24:0] _T_766 = _T_673 ? _T_761 : _T_763; // @[el2_ifu_compress_ctl.scala 338:33]
  wire  _T_772 = |io_din[6:2]; // @[el2_ifu_compress_ctl.scala 339:27]
  wire [31:0] _T_743_bits = {{7'd0}, _T_739}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_770_bits = {{7'd0}, _T_766}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_773_bits = _T_772 ? _T_743_bits : _T_770_bits; // @[el2_ifu_compress_ctl.scala 339:22]
  wire [24:0] _T_779 = {io_din[6:2],io_din[11:7],3'h0,12'he7}; // @[Cat.scala 29:58]
  wire [24:0] _T_781 = {_T_761[24:7],7'h73}; // @[Cat.scala 29:58]
  wire [24:0] _T_782 = _T_781 | 25'h100000; // @[el2_ifu_compress_ctl.scala 341:46]
  wire [24:0] _T_785 = _T_673 ? _T_779 : _T_782; // @[el2_ifu_compress_ctl.scala 342:33]
  wire [31:0] _T_755_bits = {{7'd0}, _T_750}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_789_bits = {{7'd0}, _T_785}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_792_bits = _T_772 ? _T_755_bits : _T_789_bits; // @[el2_ifu_compress_ctl.scala 343:25]
  wire [31:0] _T_794_bits = io_din[12] ? _T_792_bits : _T_773_bits; // @[el2_ifu_compress_ctl.scala 344:10]
  wire [8:0] _T_798 = {io_din[9:7],io_din[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [28:0] _T_810 = {_T_798[8:5],io_din[6:2],5'h2,3'h3,_T_798[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [7:0] _T_818 = {io_din[8:7],io_din[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_830 = {_T_818[7:5],io_din[6:2],5'h2,3'h2,_T_818[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [27:0] _T_850 = {_T_818[7:5],io_din[6:2],5'h2,3'h2,_T_818[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [4:0] _T_898 = {io_din[1:0],io_din[15:13]}; // @[Cat.scala 29:58]
  wire [31:0] _T_24_bits = {{2'd0}, _T_18}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _T_44_bits = {{4'd0}, _T_36}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_17 = 5'h1 == _T_898 ? _T_44_bits : _T_24_bits; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_66_bits = {{5'd0}, _T_58}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_22 = 5'h2 == _T_898 ? _T_66_bits : _GEN_17; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_88_bits = {{5'd0}, _T_80}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_27 = 5'h3 == _T_898 ? _T_88_bits : _GEN_22; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_119_bits = {{5'd0}, _T_111}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_32 = 5'h4 == _T_898 ? _T_119_bits : _GEN_27; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_146_bits = {{4'd0}, _T_138}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_37 = 5'h5 == _T_898 ? _T_146_bits : _GEN_32; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_177_bits = {{5'd0}, _T_169}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_42 = 5'h6 == _T_898 ? _T_177_bits : _GEN_37; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_208_bits = {{5'd0}, _T_200}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_47 = 5'h7 == _T_898 ? _T_208_bits : _GEN_42; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_52 = 5'h8 == _T_898 ? _T_219 : _GEN_47; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_57 = 5'h9 == _T_898 ? _T_306 : _GEN_52; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_62 = 5'ha == _T_898 ? _T_321 : _GEN_57; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_67 = 5'hb == _T_898 ? _T_386_bits : _GEN_62; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_72 = 5'hc == _T_898 ? _GEN_11 : _GEN_67; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_77 = 5'hd == _T_898 ? _T_533 : _GEN_72; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_82 = 5'he == _T_898 ? _T_600 : _GEN_77; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_87 = 5'hf == _T_898 ? _T_667 : _GEN_82; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_688_bits = {{6'd0}, _T_683}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_92 = 5'h10 == _T_898 ? _T_688_bits : _GEN_87; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_703_bits = {{3'd0}, _T_699}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_97 = 5'h11 == _T_898 ? _T_703_bits : _GEN_92; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_718_bits = {{4'd0}, _T_714}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_102 = 5'h12 == _T_898 ? _T_718_bits : _GEN_97; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_733_bits = {{4'd0}, _T_729}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_107 = 5'h13 == _T_898 ? _T_733_bits : _GEN_102; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_112 = 5'h14 == _T_898 ? _T_794_bits : _GEN_107; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_814_bits = {{3'd0}, _T_810}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_117 = 5'h15 == _T_898 ? _T_814_bits : _GEN_112; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_834_bits = {{4'd0}, _T_830}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_122 = 5'h16 == _T_898 ? _T_834_bits : _GEN_117; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _T_854_bits = {{4'd0}, _T_850}; // @[el2_ifu_compress_ctl.scala 225:19 el2_ifu_compress_ctl.scala 226:14]
  wire [31:0] _GEN_127 = 5'h17 == _T_898 ? _T_854_bits : _GEN_122; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_132 = 5'h18 == _T_898 ? io_din : _GEN_127; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_137 = 5'h19 == _T_898 ? io_din : _GEN_132; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_142 = 5'h1a == _T_898 ? io_din : _GEN_137; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_147 = 5'h1b == _T_898 ? io_din : _GEN_142; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_152 = 5'h1c == _T_898 ? io_din : _GEN_147; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_157 = 5'h1d == _T_898 ? io_din : _GEN_152; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_162 = 5'h1e == _T_898 ? io_din : _GEN_157; // @[el2_ifu_compress_ctl.scala 404:19]
  wire [31:0] _GEN_167 = 5'h1f == _T_898 ? io_din : _GEN_162; // @[el2_ifu_compress_ctl.scala 404:19]
  assign io_dout = _T_1 ? 32'h0 : _GEN_167; // @[el2_ifu_compress_ctl.scala 404:13]
endmodule
