module el2_lsu_trigger(
  input         clock,
  input         reset,
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_pkt,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input         io_trigger_pkt_any_0_execute,
  input         io_trigger_pkt_any_0_m,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_pkt,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input         io_trigger_pkt_any_1_execute,
  input         io_trigger_pkt_any_1_m,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_pkt,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input         io_trigger_pkt_any_2_execute,
  input         io_trigger_pkt_any_2_m,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_pkt,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input         io_trigger_pkt_any_3_execute,
  input         io_trigger_pkt_any_3_m,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_lsu_pkt_m_valid,
  input         io_lsu_pkt_m_bits_fast_int,
  input         io_lsu_pkt_m_bits_by,
  input         io_lsu_pkt_m_bits_half,
  input         io_lsu_pkt_m_bits_word,
  input         io_lsu_pkt_m_bits_dword,
  input         io_lsu_pkt_m_bits_load,
  input         io_lsu_pkt_m_bits_store,
  input         io_lsu_pkt_m_bits_unsign,
  input         io_lsu_pkt_m_bits_dma,
  input         io_lsu_pkt_m_bits_store_data_bypass_d,
  input         io_lsu_pkt_m_bits_load_ldst_bypass_d,
  input         io_lsu_pkt_m_bits_store_data_bypass_m,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_store_data_m,
  output [3:0]  io_lsu_trigger_match_m
);
  wire [15:0] _T_1 = io_lsu_pkt_m_bits_word ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_3 = _T_1 & io_store_data_m[31:16]; // @[el2_lsu_trigger.scala 16:66]
  wire  _T_4 = io_lsu_pkt_m_bits_half | io_lsu_pkt_m_bits_word; // @[el2_lsu_trigger.scala 16:124]
  wire [7:0] _T_6 = _T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_8 = _T_6 & io_store_data_m[15:8]; // @[el2_lsu_trigger.scala 16:151]
  wire [31:0] store_data_trigger_m = {_T_3,_T_8,io_store_data_m[7:0]}; // @[Cat.scala 29:58]
  wire  _T_12 = ~io_trigger_pkt_any_0_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_13 = io_trigger_pkt_any_0_select & io_trigger_pkt_any_0_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_15 = _T_12 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_16 = _T_13 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_0 = _T_15 | _T_16; // @[Mux.scala 27:72]
  wire  _T_19 = ~io_trigger_pkt_any_1_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_20 = io_trigger_pkt_any_1_select & io_trigger_pkt_any_1_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_22 = _T_19 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_23 = _T_20 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_1 = _T_22 | _T_23; // @[Mux.scala 27:72]
  wire  _T_26 = ~io_trigger_pkt_any_2_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_27 = io_trigger_pkt_any_2_select & io_trigger_pkt_any_2_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_29 = _T_26 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_30 = _T_27 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_2 = _T_29 | _T_30; // @[Mux.scala 27:72]
  wire  _T_33 = ~io_trigger_pkt_any_3_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_34 = io_trigger_pkt_any_3_select & io_trigger_pkt_any_3_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_36 = _T_33 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_37 = _T_34 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_3 = _T_36 | _T_37; // @[Mux.scala 27:72]
  wire  _T_39 = ~io_lsu_pkt_m_bits_dma; // @[el2_lsu_trigger.scala 18:71]
  wire  _T_40 = io_lsu_pkt_m_valid & _T_39; // @[el2_lsu_trigger.scala 18:69]
  wire  _T_41 = io_trigger_pkt_any_0_store & io_lsu_pkt_m_bits_store; // @[el2_lsu_trigger.scala 18:126]
  wire  _T_42 = io_trigger_pkt_any_0_load & io_lsu_pkt_m_bits_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_44 = _T_42 & _T_12; // @[el2_lsu_trigger.scala 19:58]
  wire  _T_45 = _T_41 | _T_44; // @[el2_lsu_trigger.scala 18:152]
  wire  _T_46 = _T_40 & _T_45; // @[el2_lsu_trigger.scala 18:94]
  wire  _T_49 = &io_trigger_pkt_any_0_tdata2; // @[el2_lib.scala 241:45]
  wire  _T_50 = ~_T_49; // @[el2_lib.scala 241:39]
  wire  _T_51 = io_trigger_pkt_any_0_match_pkt & _T_50; // @[el2_lib.scala 241:37]
  wire  _T_54 = io_trigger_pkt_any_0_tdata2[0] == lsu_match_data_0[0]; // @[el2_lib.scala 242:52]
  wire  _T_55 = _T_51 | _T_54; // @[el2_lib.scala 242:41]
  wire  _T_57 = &io_trigger_pkt_any_0_tdata2[0]; // @[el2_lib.scala 244:36]
  wire  _T_58 = _T_57 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_61 = io_trigger_pkt_any_0_tdata2[1] == lsu_match_data_0[1]; // @[el2_lib.scala 244:78]
  wire  _T_62 = _T_58 | _T_61; // @[el2_lib.scala 244:23]
  wire  _T_64 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[el2_lib.scala 244:36]
  wire  _T_65 = _T_64 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_68 = io_trigger_pkt_any_0_tdata2[2] == lsu_match_data_0[2]; // @[el2_lib.scala 244:78]
  wire  _T_69 = _T_65 | _T_68; // @[el2_lib.scala 244:23]
  wire  _T_71 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[el2_lib.scala 244:36]
  wire  _T_72 = _T_71 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_75 = io_trigger_pkt_any_0_tdata2[3] == lsu_match_data_0[3]; // @[el2_lib.scala 244:78]
  wire  _T_76 = _T_72 | _T_75; // @[el2_lib.scala 244:23]
  wire  _T_78 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[el2_lib.scala 244:36]
  wire  _T_79 = _T_78 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_82 = io_trigger_pkt_any_0_tdata2[4] == lsu_match_data_0[4]; // @[el2_lib.scala 244:78]
  wire  _T_83 = _T_79 | _T_82; // @[el2_lib.scala 244:23]
  wire  _T_85 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[el2_lib.scala 244:36]
  wire  _T_86 = _T_85 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_89 = io_trigger_pkt_any_0_tdata2[5] == lsu_match_data_0[5]; // @[el2_lib.scala 244:78]
  wire  _T_90 = _T_86 | _T_89; // @[el2_lib.scala 244:23]
  wire  _T_92 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[el2_lib.scala 244:36]
  wire  _T_93 = _T_92 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_96 = io_trigger_pkt_any_0_tdata2[6] == lsu_match_data_0[6]; // @[el2_lib.scala 244:78]
  wire  _T_97 = _T_93 | _T_96; // @[el2_lib.scala 244:23]
  wire  _T_99 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[el2_lib.scala 244:36]
  wire  _T_100 = _T_99 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_103 = io_trigger_pkt_any_0_tdata2[7] == lsu_match_data_0[7]; // @[el2_lib.scala 244:78]
  wire  _T_104 = _T_100 | _T_103; // @[el2_lib.scala 244:23]
  wire  _T_106 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[el2_lib.scala 244:36]
  wire  _T_107 = _T_106 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_110 = io_trigger_pkt_any_0_tdata2[8] == lsu_match_data_0[8]; // @[el2_lib.scala 244:78]
  wire  _T_111 = _T_107 | _T_110; // @[el2_lib.scala 244:23]
  wire  _T_113 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[el2_lib.scala 244:36]
  wire  _T_114 = _T_113 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_117 = io_trigger_pkt_any_0_tdata2[9] == lsu_match_data_0[9]; // @[el2_lib.scala 244:78]
  wire  _T_118 = _T_114 | _T_117; // @[el2_lib.scala 244:23]
  wire  _T_120 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[el2_lib.scala 244:36]
  wire  _T_121 = _T_120 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_124 = io_trigger_pkt_any_0_tdata2[10] == lsu_match_data_0[10]; // @[el2_lib.scala 244:78]
  wire  _T_125 = _T_121 | _T_124; // @[el2_lib.scala 244:23]
  wire  _T_127 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[el2_lib.scala 244:36]
  wire  _T_128 = _T_127 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_131 = io_trigger_pkt_any_0_tdata2[11] == lsu_match_data_0[11]; // @[el2_lib.scala 244:78]
  wire  _T_132 = _T_128 | _T_131; // @[el2_lib.scala 244:23]
  wire  _T_134 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[el2_lib.scala 244:36]
  wire  _T_135 = _T_134 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_138 = io_trigger_pkt_any_0_tdata2[12] == lsu_match_data_0[12]; // @[el2_lib.scala 244:78]
  wire  _T_139 = _T_135 | _T_138; // @[el2_lib.scala 244:23]
  wire  _T_141 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[el2_lib.scala 244:36]
  wire  _T_142 = _T_141 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_145 = io_trigger_pkt_any_0_tdata2[13] == lsu_match_data_0[13]; // @[el2_lib.scala 244:78]
  wire  _T_146 = _T_142 | _T_145; // @[el2_lib.scala 244:23]
  wire  _T_148 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[el2_lib.scala 244:36]
  wire  _T_149 = _T_148 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_152 = io_trigger_pkt_any_0_tdata2[14] == lsu_match_data_0[14]; // @[el2_lib.scala 244:78]
  wire  _T_153 = _T_149 | _T_152; // @[el2_lib.scala 244:23]
  wire  _T_155 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[el2_lib.scala 244:36]
  wire  _T_156 = _T_155 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_159 = io_trigger_pkt_any_0_tdata2[15] == lsu_match_data_0[15]; // @[el2_lib.scala 244:78]
  wire  _T_160 = _T_156 | _T_159; // @[el2_lib.scala 244:23]
  wire  _T_162 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[el2_lib.scala 244:36]
  wire  _T_163 = _T_162 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_166 = io_trigger_pkt_any_0_tdata2[16] == lsu_match_data_0[16]; // @[el2_lib.scala 244:78]
  wire  _T_167 = _T_163 | _T_166; // @[el2_lib.scala 244:23]
  wire  _T_169 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[el2_lib.scala 244:36]
  wire  _T_170 = _T_169 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_173 = io_trigger_pkt_any_0_tdata2[17] == lsu_match_data_0[17]; // @[el2_lib.scala 244:78]
  wire  _T_174 = _T_170 | _T_173; // @[el2_lib.scala 244:23]
  wire  _T_176 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[el2_lib.scala 244:36]
  wire  _T_177 = _T_176 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_180 = io_trigger_pkt_any_0_tdata2[18] == lsu_match_data_0[18]; // @[el2_lib.scala 244:78]
  wire  _T_181 = _T_177 | _T_180; // @[el2_lib.scala 244:23]
  wire  _T_183 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[el2_lib.scala 244:36]
  wire  _T_184 = _T_183 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_187 = io_trigger_pkt_any_0_tdata2[19] == lsu_match_data_0[19]; // @[el2_lib.scala 244:78]
  wire  _T_188 = _T_184 | _T_187; // @[el2_lib.scala 244:23]
  wire  _T_190 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[el2_lib.scala 244:36]
  wire  _T_191 = _T_190 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_194 = io_trigger_pkt_any_0_tdata2[20] == lsu_match_data_0[20]; // @[el2_lib.scala 244:78]
  wire  _T_195 = _T_191 | _T_194; // @[el2_lib.scala 244:23]
  wire  _T_197 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[el2_lib.scala 244:36]
  wire  _T_198 = _T_197 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_201 = io_trigger_pkt_any_0_tdata2[21] == lsu_match_data_0[21]; // @[el2_lib.scala 244:78]
  wire  _T_202 = _T_198 | _T_201; // @[el2_lib.scala 244:23]
  wire  _T_204 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[el2_lib.scala 244:36]
  wire  _T_205 = _T_204 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_208 = io_trigger_pkt_any_0_tdata2[22] == lsu_match_data_0[22]; // @[el2_lib.scala 244:78]
  wire  _T_209 = _T_205 | _T_208; // @[el2_lib.scala 244:23]
  wire  _T_211 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[el2_lib.scala 244:36]
  wire  _T_212 = _T_211 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_215 = io_trigger_pkt_any_0_tdata2[23] == lsu_match_data_0[23]; // @[el2_lib.scala 244:78]
  wire  _T_216 = _T_212 | _T_215; // @[el2_lib.scala 244:23]
  wire  _T_218 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[el2_lib.scala 244:36]
  wire  _T_219 = _T_218 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_222 = io_trigger_pkt_any_0_tdata2[24] == lsu_match_data_0[24]; // @[el2_lib.scala 244:78]
  wire  _T_223 = _T_219 | _T_222; // @[el2_lib.scala 244:23]
  wire  _T_225 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[el2_lib.scala 244:36]
  wire  _T_226 = _T_225 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_229 = io_trigger_pkt_any_0_tdata2[25] == lsu_match_data_0[25]; // @[el2_lib.scala 244:78]
  wire  _T_230 = _T_226 | _T_229; // @[el2_lib.scala 244:23]
  wire  _T_232 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[el2_lib.scala 244:36]
  wire  _T_233 = _T_232 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_236 = io_trigger_pkt_any_0_tdata2[26] == lsu_match_data_0[26]; // @[el2_lib.scala 244:78]
  wire  _T_237 = _T_233 | _T_236; // @[el2_lib.scala 244:23]
  wire  _T_239 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[el2_lib.scala 244:36]
  wire  _T_240 = _T_239 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_243 = io_trigger_pkt_any_0_tdata2[27] == lsu_match_data_0[27]; // @[el2_lib.scala 244:78]
  wire  _T_244 = _T_240 | _T_243; // @[el2_lib.scala 244:23]
  wire  _T_246 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[el2_lib.scala 244:36]
  wire  _T_247 = _T_246 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_250 = io_trigger_pkt_any_0_tdata2[28] == lsu_match_data_0[28]; // @[el2_lib.scala 244:78]
  wire  _T_251 = _T_247 | _T_250; // @[el2_lib.scala 244:23]
  wire  _T_253 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[el2_lib.scala 244:36]
  wire  _T_254 = _T_253 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_257 = io_trigger_pkt_any_0_tdata2[29] == lsu_match_data_0[29]; // @[el2_lib.scala 244:78]
  wire  _T_258 = _T_254 | _T_257; // @[el2_lib.scala 244:23]
  wire  _T_260 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[el2_lib.scala 244:36]
  wire  _T_261 = _T_260 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_264 = io_trigger_pkt_any_0_tdata2[30] == lsu_match_data_0[30]; // @[el2_lib.scala 244:78]
  wire  _T_265 = _T_261 | _T_264; // @[el2_lib.scala 244:23]
  wire  _T_267 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[el2_lib.scala 244:36]
  wire  _T_268 = _T_267 & _T_51; // @[el2_lib.scala 244:41]
  wire  _T_271 = io_trigger_pkt_any_0_tdata2[31] == lsu_match_data_0[31]; // @[el2_lib.scala 244:78]
  wire  _T_272 = _T_268 | _T_271; // @[el2_lib.scala 244:23]
  wire [7:0] _T_279 = {_T_104,_T_97,_T_90,_T_83,_T_76,_T_69,_T_62,_T_55}; // @[el2_lib.scala 245:14]
  wire [15:0] _T_287 = {_T_160,_T_153,_T_146,_T_139,_T_132,_T_125,_T_118,_T_111,_T_279}; // @[el2_lib.scala 245:14]
  wire [7:0] _T_294 = {_T_216,_T_209,_T_202,_T_195,_T_188,_T_181,_T_174,_T_167}; // @[el2_lib.scala 245:14]
  wire [31:0] _T_303 = {_T_272,_T_265,_T_258,_T_251,_T_244,_T_237,_T_230,_T_223,_T_294,_T_287}; // @[el2_lib.scala 245:14]
  wire [31:0] _GEN_0 = {{31'd0}, _T_46}; // @[el2_lsu_trigger.scala 19:92]
  wire [31:0] _T_304 = _GEN_0 & _T_303; // @[el2_lsu_trigger.scala 19:92]
  wire  _T_307 = io_trigger_pkt_any_1_store & io_lsu_pkt_m_bits_store; // @[el2_lsu_trigger.scala 18:126]
  wire  _T_308 = io_trigger_pkt_any_1_load & io_lsu_pkt_m_bits_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_310 = _T_308 & _T_19; // @[el2_lsu_trigger.scala 19:58]
  wire  _T_311 = _T_307 | _T_310; // @[el2_lsu_trigger.scala 18:152]
  wire  _T_312 = _T_40 & _T_311; // @[el2_lsu_trigger.scala 18:94]
  wire  _T_315 = &io_trigger_pkt_any_1_tdata2; // @[el2_lib.scala 241:45]
  wire  _T_316 = ~_T_315; // @[el2_lib.scala 241:39]
  wire  _T_317 = io_trigger_pkt_any_1_match_pkt & _T_316; // @[el2_lib.scala 241:37]
  wire  _T_320 = io_trigger_pkt_any_1_tdata2[0] == lsu_match_data_1[0]; // @[el2_lib.scala 242:52]
  wire  _T_321 = _T_317 | _T_320; // @[el2_lib.scala 242:41]
  wire  _T_323 = &io_trigger_pkt_any_1_tdata2[0]; // @[el2_lib.scala 244:36]
  wire  _T_324 = _T_323 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_327 = io_trigger_pkt_any_1_tdata2[1] == lsu_match_data_1[1]; // @[el2_lib.scala 244:78]
  wire  _T_328 = _T_324 | _T_327; // @[el2_lib.scala 244:23]
  wire  _T_330 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[el2_lib.scala 244:36]
  wire  _T_331 = _T_330 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_334 = io_trigger_pkt_any_1_tdata2[2] == lsu_match_data_1[2]; // @[el2_lib.scala 244:78]
  wire  _T_335 = _T_331 | _T_334; // @[el2_lib.scala 244:23]
  wire  _T_337 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[el2_lib.scala 244:36]
  wire  _T_338 = _T_337 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_341 = io_trigger_pkt_any_1_tdata2[3] == lsu_match_data_1[3]; // @[el2_lib.scala 244:78]
  wire  _T_342 = _T_338 | _T_341; // @[el2_lib.scala 244:23]
  wire  _T_344 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[el2_lib.scala 244:36]
  wire  _T_345 = _T_344 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_348 = io_trigger_pkt_any_1_tdata2[4] == lsu_match_data_1[4]; // @[el2_lib.scala 244:78]
  wire  _T_349 = _T_345 | _T_348; // @[el2_lib.scala 244:23]
  wire  _T_351 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[el2_lib.scala 244:36]
  wire  _T_352 = _T_351 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_355 = io_trigger_pkt_any_1_tdata2[5] == lsu_match_data_1[5]; // @[el2_lib.scala 244:78]
  wire  _T_356 = _T_352 | _T_355; // @[el2_lib.scala 244:23]
  wire  _T_358 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[el2_lib.scala 244:36]
  wire  _T_359 = _T_358 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_362 = io_trigger_pkt_any_1_tdata2[6] == lsu_match_data_1[6]; // @[el2_lib.scala 244:78]
  wire  _T_363 = _T_359 | _T_362; // @[el2_lib.scala 244:23]
  wire  _T_365 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[el2_lib.scala 244:36]
  wire  _T_366 = _T_365 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_369 = io_trigger_pkt_any_1_tdata2[7] == lsu_match_data_1[7]; // @[el2_lib.scala 244:78]
  wire  _T_370 = _T_366 | _T_369; // @[el2_lib.scala 244:23]
  wire  _T_372 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[el2_lib.scala 244:36]
  wire  _T_373 = _T_372 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_376 = io_trigger_pkt_any_1_tdata2[8] == lsu_match_data_1[8]; // @[el2_lib.scala 244:78]
  wire  _T_377 = _T_373 | _T_376; // @[el2_lib.scala 244:23]
  wire  _T_379 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[el2_lib.scala 244:36]
  wire  _T_380 = _T_379 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_383 = io_trigger_pkt_any_1_tdata2[9] == lsu_match_data_1[9]; // @[el2_lib.scala 244:78]
  wire  _T_384 = _T_380 | _T_383; // @[el2_lib.scala 244:23]
  wire  _T_386 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[el2_lib.scala 244:36]
  wire  _T_387 = _T_386 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_390 = io_trigger_pkt_any_1_tdata2[10] == lsu_match_data_1[10]; // @[el2_lib.scala 244:78]
  wire  _T_391 = _T_387 | _T_390; // @[el2_lib.scala 244:23]
  wire  _T_393 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[el2_lib.scala 244:36]
  wire  _T_394 = _T_393 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_397 = io_trigger_pkt_any_1_tdata2[11] == lsu_match_data_1[11]; // @[el2_lib.scala 244:78]
  wire  _T_398 = _T_394 | _T_397; // @[el2_lib.scala 244:23]
  wire  _T_400 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[el2_lib.scala 244:36]
  wire  _T_401 = _T_400 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_404 = io_trigger_pkt_any_1_tdata2[12] == lsu_match_data_1[12]; // @[el2_lib.scala 244:78]
  wire  _T_405 = _T_401 | _T_404; // @[el2_lib.scala 244:23]
  wire  _T_407 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[el2_lib.scala 244:36]
  wire  _T_408 = _T_407 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_411 = io_trigger_pkt_any_1_tdata2[13] == lsu_match_data_1[13]; // @[el2_lib.scala 244:78]
  wire  _T_412 = _T_408 | _T_411; // @[el2_lib.scala 244:23]
  wire  _T_414 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[el2_lib.scala 244:36]
  wire  _T_415 = _T_414 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_418 = io_trigger_pkt_any_1_tdata2[14] == lsu_match_data_1[14]; // @[el2_lib.scala 244:78]
  wire  _T_419 = _T_415 | _T_418; // @[el2_lib.scala 244:23]
  wire  _T_421 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[el2_lib.scala 244:36]
  wire  _T_422 = _T_421 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_425 = io_trigger_pkt_any_1_tdata2[15] == lsu_match_data_1[15]; // @[el2_lib.scala 244:78]
  wire  _T_426 = _T_422 | _T_425; // @[el2_lib.scala 244:23]
  wire  _T_428 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[el2_lib.scala 244:36]
  wire  _T_429 = _T_428 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_432 = io_trigger_pkt_any_1_tdata2[16] == lsu_match_data_1[16]; // @[el2_lib.scala 244:78]
  wire  _T_433 = _T_429 | _T_432; // @[el2_lib.scala 244:23]
  wire  _T_435 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[el2_lib.scala 244:36]
  wire  _T_436 = _T_435 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_439 = io_trigger_pkt_any_1_tdata2[17] == lsu_match_data_1[17]; // @[el2_lib.scala 244:78]
  wire  _T_440 = _T_436 | _T_439; // @[el2_lib.scala 244:23]
  wire  _T_442 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[el2_lib.scala 244:36]
  wire  _T_443 = _T_442 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_446 = io_trigger_pkt_any_1_tdata2[18] == lsu_match_data_1[18]; // @[el2_lib.scala 244:78]
  wire  _T_447 = _T_443 | _T_446; // @[el2_lib.scala 244:23]
  wire  _T_449 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[el2_lib.scala 244:36]
  wire  _T_450 = _T_449 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_453 = io_trigger_pkt_any_1_tdata2[19] == lsu_match_data_1[19]; // @[el2_lib.scala 244:78]
  wire  _T_454 = _T_450 | _T_453; // @[el2_lib.scala 244:23]
  wire  _T_456 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[el2_lib.scala 244:36]
  wire  _T_457 = _T_456 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_460 = io_trigger_pkt_any_1_tdata2[20] == lsu_match_data_1[20]; // @[el2_lib.scala 244:78]
  wire  _T_461 = _T_457 | _T_460; // @[el2_lib.scala 244:23]
  wire  _T_463 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[el2_lib.scala 244:36]
  wire  _T_464 = _T_463 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_467 = io_trigger_pkt_any_1_tdata2[21] == lsu_match_data_1[21]; // @[el2_lib.scala 244:78]
  wire  _T_468 = _T_464 | _T_467; // @[el2_lib.scala 244:23]
  wire  _T_470 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[el2_lib.scala 244:36]
  wire  _T_471 = _T_470 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_474 = io_trigger_pkt_any_1_tdata2[22] == lsu_match_data_1[22]; // @[el2_lib.scala 244:78]
  wire  _T_475 = _T_471 | _T_474; // @[el2_lib.scala 244:23]
  wire  _T_477 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[el2_lib.scala 244:36]
  wire  _T_478 = _T_477 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_481 = io_trigger_pkt_any_1_tdata2[23] == lsu_match_data_1[23]; // @[el2_lib.scala 244:78]
  wire  _T_482 = _T_478 | _T_481; // @[el2_lib.scala 244:23]
  wire  _T_484 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[el2_lib.scala 244:36]
  wire  _T_485 = _T_484 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_488 = io_trigger_pkt_any_1_tdata2[24] == lsu_match_data_1[24]; // @[el2_lib.scala 244:78]
  wire  _T_489 = _T_485 | _T_488; // @[el2_lib.scala 244:23]
  wire  _T_491 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[el2_lib.scala 244:36]
  wire  _T_492 = _T_491 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_495 = io_trigger_pkt_any_1_tdata2[25] == lsu_match_data_1[25]; // @[el2_lib.scala 244:78]
  wire  _T_496 = _T_492 | _T_495; // @[el2_lib.scala 244:23]
  wire  _T_498 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[el2_lib.scala 244:36]
  wire  _T_499 = _T_498 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_502 = io_trigger_pkt_any_1_tdata2[26] == lsu_match_data_1[26]; // @[el2_lib.scala 244:78]
  wire  _T_503 = _T_499 | _T_502; // @[el2_lib.scala 244:23]
  wire  _T_505 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[el2_lib.scala 244:36]
  wire  _T_506 = _T_505 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_509 = io_trigger_pkt_any_1_tdata2[27] == lsu_match_data_1[27]; // @[el2_lib.scala 244:78]
  wire  _T_510 = _T_506 | _T_509; // @[el2_lib.scala 244:23]
  wire  _T_512 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[el2_lib.scala 244:36]
  wire  _T_513 = _T_512 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_516 = io_trigger_pkt_any_1_tdata2[28] == lsu_match_data_1[28]; // @[el2_lib.scala 244:78]
  wire  _T_517 = _T_513 | _T_516; // @[el2_lib.scala 244:23]
  wire  _T_519 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[el2_lib.scala 244:36]
  wire  _T_520 = _T_519 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_523 = io_trigger_pkt_any_1_tdata2[29] == lsu_match_data_1[29]; // @[el2_lib.scala 244:78]
  wire  _T_524 = _T_520 | _T_523; // @[el2_lib.scala 244:23]
  wire  _T_526 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[el2_lib.scala 244:36]
  wire  _T_527 = _T_526 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_530 = io_trigger_pkt_any_1_tdata2[30] == lsu_match_data_1[30]; // @[el2_lib.scala 244:78]
  wire  _T_531 = _T_527 | _T_530; // @[el2_lib.scala 244:23]
  wire  _T_533 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[el2_lib.scala 244:36]
  wire  _T_534 = _T_533 & _T_317; // @[el2_lib.scala 244:41]
  wire  _T_537 = io_trigger_pkt_any_1_tdata2[31] == lsu_match_data_1[31]; // @[el2_lib.scala 244:78]
  wire  _T_538 = _T_534 | _T_537; // @[el2_lib.scala 244:23]
  wire [7:0] _T_545 = {_T_370,_T_363,_T_356,_T_349,_T_342,_T_335,_T_328,_T_321}; // @[el2_lib.scala 245:14]
  wire [15:0] _T_553 = {_T_426,_T_419,_T_412,_T_405,_T_398,_T_391,_T_384,_T_377,_T_545}; // @[el2_lib.scala 245:14]
  wire [7:0] _T_560 = {_T_482,_T_475,_T_468,_T_461,_T_454,_T_447,_T_440,_T_433}; // @[el2_lib.scala 245:14]
  wire [31:0] _T_569 = {_T_538,_T_531,_T_524,_T_517,_T_510,_T_503,_T_496,_T_489,_T_560,_T_553}; // @[el2_lib.scala 245:14]
  wire [31:0] _GEN_1 = {{31'd0}, _T_312}; // @[el2_lsu_trigger.scala 19:92]
  wire [31:0] _T_570 = _GEN_1 & _T_569; // @[el2_lsu_trigger.scala 19:92]
  wire  _T_573 = io_trigger_pkt_any_2_store & io_lsu_pkt_m_bits_store; // @[el2_lsu_trigger.scala 18:126]
  wire  _T_574 = io_trigger_pkt_any_2_load & io_lsu_pkt_m_bits_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_576 = _T_574 & _T_26; // @[el2_lsu_trigger.scala 19:58]
  wire  _T_577 = _T_573 | _T_576; // @[el2_lsu_trigger.scala 18:152]
  wire  _T_578 = _T_40 & _T_577; // @[el2_lsu_trigger.scala 18:94]
  wire  _T_581 = &io_trigger_pkt_any_2_tdata2; // @[el2_lib.scala 241:45]
  wire  _T_582 = ~_T_581; // @[el2_lib.scala 241:39]
  wire  _T_583 = io_trigger_pkt_any_2_match_pkt & _T_582; // @[el2_lib.scala 241:37]
  wire  _T_586 = io_trigger_pkt_any_2_tdata2[0] == lsu_match_data_2[0]; // @[el2_lib.scala 242:52]
  wire  _T_587 = _T_583 | _T_586; // @[el2_lib.scala 242:41]
  wire  _T_589 = &io_trigger_pkt_any_2_tdata2[0]; // @[el2_lib.scala 244:36]
  wire  _T_590 = _T_589 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_593 = io_trigger_pkt_any_2_tdata2[1] == lsu_match_data_2[1]; // @[el2_lib.scala 244:78]
  wire  _T_594 = _T_590 | _T_593; // @[el2_lib.scala 244:23]
  wire  _T_596 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[el2_lib.scala 244:36]
  wire  _T_597 = _T_596 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_600 = io_trigger_pkt_any_2_tdata2[2] == lsu_match_data_2[2]; // @[el2_lib.scala 244:78]
  wire  _T_601 = _T_597 | _T_600; // @[el2_lib.scala 244:23]
  wire  _T_603 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[el2_lib.scala 244:36]
  wire  _T_604 = _T_603 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_607 = io_trigger_pkt_any_2_tdata2[3] == lsu_match_data_2[3]; // @[el2_lib.scala 244:78]
  wire  _T_608 = _T_604 | _T_607; // @[el2_lib.scala 244:23]
  wire  _T_610 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[el2_lib.scala 244:36]
  wire  _T_611 = _T_610 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_614 = io_trigger_pkt_any_2_tdata2[4] == lsu_match_data_2[4]; // @[el2_lib.scala 244:78]
  wire  _T_615 = _T_611 | _T_614; // @[el2_lib.scala 244:23]
  wire  _T_617 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[el2_lib.scala 244:36]
  wire  _T_618 = _T_617 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_621 = io_trigger_pkt_any_2_tdata2[5] == lsu_match_data_2[5]; // @[el2_lib.scala 244:78]
  wire  _T_622 = _T_618 | _T_621; // @[el2_lib.scala 244:23]
  wire  _T_624 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[el2_lib.scala 244:36]
  wire  _T_625 = _T_624 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_628 = io_trigger_pkt_any_2_tdata2[6] == lsu_match_data_2[6]; // @[el2_lib.scala 244:78]
  wire  _T_629 = _T_625 | _T_628; // @[el2_lib.scala 244:23]
  wire  _T_631 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[el2_lib.scala 244:36]
  wire  _T_632 = _T_631 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_635 = io_trigger_pkt_any_2_tdata2[7] == lsu_match_data_2[7]; // @[el2_lib.scala 244:78]
  wire  _T_636 = _T_632 | _T_635; // @[el2_lib.scala 244:23]
  wire  _T_638 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[el2_lib.scala 244:36]
  wire  _T_639 = _T_638 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_642 = io_trigger_pkt_any_2_tdata2[8] == lsu_match_data_2[8]; // @[el2_lib.scala 244:78]
  wire  _T_643 = _T_639 | _T_642; // @[el2_lib.scala 244:23]
  wire  _T_645 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[el2_lib.scala 244:36]
  wire  _T_646 = _T_645 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_649 = io_trigger_pkt_any_2_tdata2[9] == lsu_match_data_2[9]; // @[el2_lib.scala 244:78]
  wire  _T_650 = _T_646 | _T_649; // @[el2_lib.scala 244:23]
  wire  _T_652 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[el2_lib.scala 244:36]
  wire  _T_653 = _T_652 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_656 = io_trigger_pkt_any_2_tdata2[10] == lsu_match_data_2[10]; // @[el2_lib.scala 244:78]
  wire  _T_657 = _T_653 | _T_656; // @[el2_lib.scala 244:23]
  wire  _T_659 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[el2_lib.scala 244:36]
  wire  _T_660 = _T_659 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_663 = io_trigger_pkt_any_2_tdata2[11] == lsu_match_data_2[11]; // @[el2_lib.scala 244:78]
  wire  _T_664 = _T_660 | _T_663; // @[el2_lib.scala 244:23]
  wire  _T_666 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[el2_lib.scala 244:36]
  wire  _T_667 = _T_666 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_670 = io_trigger_pkt_any_2_tdata2[12] == lsu_match_data_2[12]; // @[el2_lib.scala 244:78]
  wire  _T_671 = _T_667 | _T_670; // @[el2_lib.scala 244:23]
  wire  _T_673 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[el2_lib.scala 244:36]
  wire  _T_674 = _T_673 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_677 = io_trigger_pkt_any_2_tdata2[13] == lsu_match_data_2[13]; // @[el2_lib.scala 244:78]
  wire  _T_678 = _T_674 | _T_677; // @[el2_lib.scala 244:23]
  wire  _T_680 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[el2_lib.scala 244:36]
  wire  _T_681 = _T_680 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_684 = io_trigger_pkt_any_2_tdata2[14] == lsu_match_data_2[14]; // @[el2_lib.scala 244:78]
  wire  _T_685 = _T_681 | _T_684; // @[el2_lib.scala 244:23]
  wire  _T_687 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[el2_lib.scala 244:36]
  wire  _T_688 = _T_687 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_691 = io_trigger_pkt_any_2_tdata2[15] == lsu_match_data_2[15]; // @[el2_lib.scala 244:78]
  wire  _T_692 = _T_688 | _T_691; // @[el2_lib.scala 244:23]
  wire  _T_694 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[el2_lib.scala 244:36]
  wire  _T_695 = _T_694 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_698 = io_trigger_pkt_any_2_tdata2[16] == lsu_match_data_2[16]; // @[el2_lib.scala 244:78]
  wire  _T_699 = _T_695 | _T_698; // @[el2_lib.scala 244:23]
  wire  _T_701 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[el2_lib.scala 244:36]
  wire  _T_702 = _T_701 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_705 = io_trigger_pkt_any_2_tdata2[17] == lsu_match_data_2[17]; // @[el2_lib.scala 244:78]
  wire  _T_706 = _T_702 | _T_705; // @[el2_lib.scala 244:23]
  wire  _T_708 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[el2_lib.scala 244:36]
  wire  _T_709 = _T_708 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_712 = io_trigger_pkt_any_2_tdata2[18] == lsu_match_data_2[18]; // @[el2_lib.scala 244:78]
  wire  _T_713 = _T_709 | _T_712; // @[el2_lib.scala 244:23]
  wire  _T_715 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[el2_lib.scala 244:36]
  wire  _T_716 = _T_715 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_719 = io_trigger_pkt_any_2_tdata2[19] == lsu_match_data_2[19]; // @[el2_lib.scala 244:78]
  wire  _T_720 = _T_716 | _T_719; // @[el2_lib.scala 244:23]
  wire  _T_722 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[el2_lib.scala 244:36]
  wire  _T_723 = _T_722 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_726 = io_trigger_pkt_any_2_tdata2[20] == lsu_match_data_2[20]; // @[el2_lib.scala 244:78]
  wire  _T_727 = _T_723 | _T_726; // @[el2_lib.scala 244:23]
  wire  _T_729 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[el2_lib.scala 244:36]
  wire  _T_730 = _T_729 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_733 = io_trigger_pkt_any_2_tdata2[21] == lsu_match_data_2[21]; // @[el2_lib.scala 244:78]
  wire  _T_734 = _T_730 | _T_733; // @[el2_lib.scala 244:23]
  wire  _T_736 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[el2_lib.scala 244:36]
  wire  _T_737 = _T_736 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_740 = io_trigger_pkt_any_2_tdata2[22] == lsu_match_data_2[22]; // @[el2_lib.scala 244:78]
  wire  _T_741 = _T_737 | _T_740; // @[el2_lib.scala 244:23]
  wire  _T_743 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[el2_lib.scala 244:36]
  wire  _T_744 = _T_743 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_747 = io_trigger_pkt_any_2_tdata2[23] == lsu_match_data_2[23]; // @[el2_lib.scala 244:78]
  wire  _T_748 = _T_744 | _T_747; // @[el2_lib.scala 244:23]
  wire  _T_750 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[el2_lib.scala 244:36]
  wire  _T_751 = _T_750 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_754 = io_trigger_pkt_any_2_tdata2[24] == lsu_match_data_2[24]; // @[el2_lib.scala 244:78]
  wire  _T_755 = _T_751 | _T_754; // @[el2_lib.scala 244:23]
  wire  _T_757 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[el2_lib.scala 244:36]
  wire  _T_758 = _T_757 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_761 = io_trigger_pkt_any_2_tdata2[25] == lsu_match_data_2[25]; // @[el2_lib.scala 244:78]
  wire  _T_762 = _T_758 | _T_761; // @[el2_lib.scala 244:23]
  wire  _T_764 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[el2_lib.scala 244:36]
  wire  _T_765 = _T_764 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_768 = io_trigger_pkt_any_2_tdata2[26] == lsu_match_data_2[26]; // @[el2_lib.scala 244:78]
  wire  _T_769 = _T_765 | _T_768; // @[el2_lib.scala 244:23]
  wire  _T_771 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[el2_lib.scala 244:36]
  wire  _T_772 = _T_771 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_775 = io_trigger_pkt_any_2_tdata2[27] == lsu_match_data_2[27]; // @[el2_lib.scala 244:78]
  wire  _T_776 = _T_772 | _T_775; // @[el2_lib.scala 244:23]
  wire  _T_778 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[el2_lib.scala 244:36]
  wire  _T_779 = _T_778 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_782 = io_trigger_pkt_any_2_tdata2[28] == lsu_match_data_2[28]; // @[el2_lib.scala 244:78]
  wire  _T_783 = _T_779 | _T_782; // @[el2_lib.scala 244:23]
  wire  _T_785 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[el2_lib.scala 244:36]
  wire  _T_786 = _T_785 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_789 = io_trigger_pkt_any_2_tdata2[29] == lsu_match_data_2[29]; // @[el2_lib.scala 244:78]
  wire  _T_790 = _T_786 | _T_789; // @[el2_lib.scala 244:23]
  wire  _T_792 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[el2_lib.scala 244:36]
  wire  _T_793 = _T_792 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_796 = io_trigger_pkt_any_2_tdata2[30] == lsu_match_data_2[30]; // @[el2_lib.scala 244:78]
  wire  _T_797 = _T_793 | _T_796; // @[el2_lib.scala 244:23]
  wire  _T_799 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[el2_lib.scala 244:36]
  wire  _T_800 = _T_799 & _T_583; // @[el2_lib.scala 244:41]
  wire  _T_803 = io_trigger_pkt_any_2_tdata2[31] == lsu_match_data_2[31]; // @[el2_lib.scala 244:78]
  wire  _T_804 = _T_800 | _T_803; // @[el2_lib.scala 244:23]
  wire [7:0] _T_811 = {_T_636,_T_629,_T_622,_T_615,_T_608,_T_601,_T_594,_T_587}; // @[el2_lib.scala 245:14]
  wire [15:0] _T_819 = {_T_692,_T_685,_T_678,_T_671,_T_664,_T_657,_T_650,_T_643,_T_811}; // @[el2_lib.scala 245:14]
  wire [7:0] _T_826 = {_T_748,_T_741,_T_734,_T_727,_T_720,_T_713,_T_706,_T_699}; // @[el2_lib.scala 245:14]
  wire [31:0] _T_835 = {_T_804,_T_797,_T_790,_T_783,_T_776,_T_769,_T_762,_T_755,_T_826,_T_819}; // @[el2_lib.scala 245:14]
  wire [31:0] _GEN_2 = {{31'd0}, _T_578}; // @[el2_lsu_trigger.scala 19:92]
  wire [31:0] _T_836 = _GEN_2 & _T_835; // @[el2_lsu_trigger.scala 19:92]
  wire  _T_839 = io_trigger_pkt_any_3_store & io_lsu_pkt_m_bits_store; // @[el2_lsu_trigger.scala 18:126]
  wire  _T_840 = io_trigger_pkt_any_3_load & io_lsu_pkt_m_bits_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_842 = _T_840 & _T_33; // @[el2_lsu_trigger.scala 19:58]
  wire  _T_843 = _T_839 | _T_842; // @[el2_lsu_trigger.scala 18:152]
  wire  _T_844 = _T_40 & _T_843; // @[el2_lsu_trigger.scala 18:94]
  wire  _T_847 = &io_trigger_pkt_any_3_tdata2; // @[el2_lib.scala 241:45]
  wire  _T_848 = ~_T_847; // @[el2_lib.scala 241:39]
  wire  _T_849 = io_trigger_pkt_any_3_match_pkt & _T_848; // @[el2_lib.scala 241:37]
  wire  _T_852 = io_trigger_pkt_any_3_tdata2[0] == lsu_match_data_3[0]; // @[el2_lib.scala 242:52]
  wire  _T_853 = _T_849 | _T_852; // @[el2_lib.scala 242:41]
  wire  _T_855 = &io_trigger_pkt_any_3_tdata2[0]; // @[el2_lib.scala 244:36]
  wire  _T_856 = _T_855 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_859 = io_trigger_pkt_any_3_tdata2[1] == lsu_match_data_3[1]; // @[el2_lib.scala 244:78]
  wire  _T_860 = _T_856 | _T_859; // @[el2_lib.scala 244:23]
  wire  _T_862 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[el2_lib.scala 244:36]
  wire  _T_863 = _T_862 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_866 = io_trigger_pkt_any_3_tdata2[2] == lsu_match_data_3[2]; // @[el2_lib.scala 244:78]
  wire  _T_867 = _T_863 | _T_866; // @[el2_lib.scala 244:23]
  wire  _T_869 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[el2_lib.scala 244:36]
  wire  _T_870 = _T_869 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_873 = io_trigger_pkt_any_3_tdata2[3] == lsu_match_data_3[3]; // @[el2_lib.scala 244:78]
  wire  _T_874 = _T_870 | _T_873; // @[el2_lib.scala 244:23]
  wire  _T_876 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[el2_lib.scala 244:36]
  wire  _T_877 = _T_876 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_880 = io_trigger_pkt_any_3_tdata2[4] == lsu_match_data_3[4]; // @[el2_lib.scala 244:78]
  wire  _T_881 = _T_877 | _T_880; // @[el2_lib.scala 244:23]
  wire  _T_883 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[el2_lib.scala 244:36]
  wire  _T_884 = _T_883 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_887 = io_trigger_pkt_any_3_tdata2[5] == lsu_match_data_3[5]; // @[el2_lib.scala 244:78]
  wire  _T_888 = _T_884 | _T_887; // @[el2_lib.scala 244:23]
  wire  _T_890 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[el2_lib.scala 244:36]
  wire  _T_891 = _T_890 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_894 = io_trigger_pkt_any_3_tdata2[6] == lsu_match_data_3[6]; // @[el2_lib.scala 244:78]
  wire  _T_895 = _T_891 | _T_894; // @[el2_lib.scala 244:23]
  wire  _T_897 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[el2_lib.scala 244:36]
  wire  _T_898 = _T_897 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_901 = io_trigger_pkt_any_3_tdata2[7] == lsu_match_data_3[7]; // @[el2_lib.scala 244:78]
  wire  _T_902 = _T_898 | _T_901; // @[el2_lib.scala 244:23]
  wire  _T_904 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[el2_lib.scala 244:36]
  wire  _T_905 = _T_904 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_908 = io_trigger_pkt_any_3_tdata2[8] == lsu_match_data_3[8]; // @[el2_lib.scala 244:78]
  wire  _T_909 = _T_905 | _T_908; // @[el2_lib.scala 244:23]
  wire  _T_911 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[el2_lib.scala 244:36]
  wire  _T_912 = _T_911 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_915 = io_trigger_pkt_any_3_tdata2[9] == lsu_match_data_3[9]; // @[el2_lib.scala 244:78]
  wire  _T_916 = _T_912 | _T_915; // @[el2_lib.scala 244:23]
  wire  _T_918 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[el2_lib.scala 244:36]
  wire  _T_919 = _T_918 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_922 = io_trigger_pkt_any_3_tdata2[10] == lsu_match_data_3[10]; // @[el2_lib.scala 244:78]
  wire  _T_923 = _T_919 | _T_922; // @[el2_lib.scala 244:23]
  wire  _T_925 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[el2_lib.scala 244:36]
  wire  _T_926 = _T_925 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_929 = io_trigger_pkt_any_3_tdata2[11] == lsu_match_data_3[11]; // @[el2_lib.scala 244:78]
  wire  _T_930 = _T_926 | _T_929; // @[el2_lib.scala 244:23]
  wire  _T_932 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[el2_lib.scala 244:36]
  wire  _T_933 = _T_932 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_936 = io_trigger_pkt_any_3_tdata2[12] == lsu_match_data_3[12]; // @[el2_lib.scala 244:78]
  wire  _T_937 = _T_933 | _T_936; // @[el2_lib.scala 244:23]
  wire  _T_939 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[el2_lib.scala 244:36]
  wire  _T_940 = _T_939 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_943 = io_trigger_pkt_any_3_tdata2[13] == lsu_match_data_3[13]; // @[el2_lib.scala 244:78]
  wire  _T_944 = _T_940 | _T_943; // @[el2_lib.scala 244:23]
  wire  _T_946 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[el2_lib.scala 244:36]
  wire  _T_947 = _T_946 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_950 = io_trigger_pkt_any_3_tdata2[14] == lsu_match_data_3[14]; // @[el2_lib.scala 244:78]
  wire  _T_951 = _T_947 | _T_950; // @[el2_lib.scala 244:23]
  wire  _T_953 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[el2_lib.scala 244:36]
  wire  _T_954 = _T_953 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_957 = io_trigger_pkt_any_3_tdata2[15] == lsu_match_data_3[15]; // @[el2_lib.scala 244:78]
  wire  _T_958 = _T_954 | _T_957; // @[el2_lib.scala 244:23]
  wire  _T_960 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[el2_lib.scala 244:36]
  wire  _T_961 = _T_960 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_964 = io_trigger_pkt_any_3_tdata2[16] == lsu_match_data_3[16]; // @[el2_lib.scala 244:78]
  wire  _T_965 = _T_961 | _T_964; // @[el2_lib.scala 244:23]
  wire  _T_967 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[el2_lib.scala 244:36]
  wire  _T_968 = _T_967 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_971 = io_trigger_pkt_any_3_tdata2[17] == lsu_match_data_3[17]; // @[el2_lib.scala 244:78]
  wire  _T_972 = _T_968 | _T_971; // @[el2_lib.scala 244:23]
  wire  _T_974 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[el2_lib.scala 244:36]
  wire  _T_975 = _T_974 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_978 = io_trigger_pkt_any_3_tdata2[18] == lsu_match_data_3[18]; // @[el2_lib.scala 244:78]
  wire  _T_979 = _T_975 | _T_978; // @[el2_lib.scala 244:23]
  wire  _T_981 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[el2_lib.scala 244:36]
  wire  _T_982 = _T_981 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_985 = io_trigger_pkt_any_3_tdata2[19] == lsu_match_data_3[19]; // @[el2_lib.scala 244:78]
  wire  _T_986 = _T_982 | _T_985; // @[el2_lib.scala 244:23]
  wire  _T_988 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[el2_lib.scala 244:36]
  wire  _T_989 = _T_988 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_992 = io_trigger_pkt_any_3_tdata2[20] == lsu_match_data_3[20]; // @[el2_lib.scala 244:78]
  wire  _T_993 = _T_989 | _T_992; // @[el2_lib.scala 244:23]
  wire  _T_995 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[el2_lib.scala 244:36]
  wire  _T_996 = _T_995 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_999 = io_trigger_pkt_any_3_tdata2[21] == lsu_match_data_3[21]; // @[el2_lib.scala 244:78]
  wire  _T_1000 = _T_996 | _T_999; // @[el2_lib.scala 244:23]
  wire  _T_1002 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[el2_lib.scala 244:36]
  wire  _T_1003 = _T_1002 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1006 = io_trigger_pkt_any_3_tdata2[22] == lsu_match_data_3[22]; // @[el2_lib.scala 244:78]
  wire  _T_1007 = _T_1003 | _T_1006; // @[el2_lib.scala 244:23]
  wire  _T_1009 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[el2_lib.scala 244:36]
  wire  _T_1010 = _T_1009 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1013 = io_trigger_pkt_any_3_tdata2[23] == lsu_match_data_3[23]; // @[el2_lib.scala 244:78]
  wire  _T_1014 = _T_1010 | _T_1013; // @[el2_lib.scala 244:23]
  wire  _T_1016 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[el2_lib.scala 244:36]
  wire  _T_1017 = _T_1016 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1020 = io_trigger_pkt_any_3_tdata2[24] == lsu_match_data_3[24]; // @[el2_lib.scala 244:78]
  wire  _T_1021 = _T_1017 | _T_1020; // @[el2_lib.scala 244:23]
  wire  _T_1023 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[el2_lib.scala 244:36]
  wire  _T_1024 = _T_1023 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1027 = io_trigger_pkt_any_3_tdata2[25] == lsu_match_data_3[25]; // @[el2_lib.scala 244:78]
  wire  _T_1028 = _T_1024 | _T_1027; // @[el2_lib.scala 244:23]
  wire  _T_1030 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[el2_lib.scala 244:36]
  wire  _T_1031 = _T_1030 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1034 = io_trigger_pkt_any_3_tdata2[26] == lsu_match_data_3[26]; // @[el2_lib.scala 244:78]
  wire  _T_1035 = _T_1031 | _T_1034; // @[el2_lib.scala 244:23]
  wire  _T_1037 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[el2_lib.scala 244:36]
  wire  _T_1038 = _T_1037 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1041 = io_trigger_pkt_any_3_tdata2[27] == lsu_match_data_3[27]; // @[el2_lib.scala 244:78]
  wire  _T_1042 = _T_1038 | _T_1041; // @[el2_lib.scala 244:23]
  wire  _T_1044 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[el2_lib.scala 244:36]
  wire  _T_1045 = _T_1044 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1048 = io_trigger_pkt_any_3_tdata2[28] == lsu_match_data_3[28]; // @[el2_lib.scala 244:78]
  wire  _T_1049 = _T_1045 | _T_1048; // @[el2_lib.scala 244:23]
  wire  _T_1051 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[el2_lib.scala 244:36]
  wire  _T_1052 = _T_1051 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1055 = io_trigger_pkt_any_3_tdata2[29] == lsu_match_data_3[29]; // @[el2_lib.scala 244:78]
  wire  _T_1056 = _T_1052 | _T_1055; // @[el2_lib.scala 244:23]
  wire  _T_1058 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[el2_lib.scala 244:36]
  wire  _T_1059 = _T_1058 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1062 = io_trigger_pkt_any_3_tdata2[30] == lsu_match_data_3[30]; // @[el2_lib.scala 244:78]
  wire  _T_1063 = _T_1059 | _T_1062; // @[el2_lib.scala 244:23]
  wire  _T_1065 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[el2_lib.scala 244:36]
  wire  _T_1066 = _T_1065 & _T_849; // @[el2_lib.scala 244:41]
  wire  _T_1069 = io_trigger_pkt_any_3_tdata2[31] == lsu_match_data_3[31]; // @[el2_lib.scala 244:78]
  wire  _T_1070 = _T_1066 | _T_1069; // @[el2_lib.scala 244:23]
  wire [7:0] _T_1077 = {_T_902,_T_895,_T_888,_T_881,_T_874,_T_867,_T_860,_T_853}; // @[el2_lib.scala 245:14]
  wire [15:0] _T_1085 = {_T_958,_T_951,_T_944,_T_937,_T_930,_T_923,_T_916,_T_909,_T_1077}; // @[el2_lib.scala 245:14]
  wire [7:0] _T_1092 = {_T_1014,_T_1007,_T_1000,_T_993,_T_986,_T_979,_T_972,_T_965}; // @[el2_lib.scala 245:14]
  wire [31:0] _T_1101 = {_T_1070,_T_1063,_T_1056,_T_1049,_T_1042,_T_1035,_T_1028,_T_1021,_T_1092,_T_1085}; // @[el2_lib.scala 245:14]
  wire [31:0] _GEN_3 = {{31'd0}, _T_844}; // @[el2_lsu_trigger.scala 19:92]
  wire [31:0] _T_1102 = _GEN_3 & _T_1101; // @[el2_lsu_trigger.scala 19:92]
  wire [127:0] _T_1105 = {_T_1102,_T_836,_T_570,_T_304}; // @[Cat.scala 29:58]
  assign io_lsu_trigger_match_m = _T_1105[3:0]; // @[el2_lsu_trigger.scala 18:26]
endmodule
