module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [63:0] _RAND_176;
  reg [63:0] _RAND_177;
  reg [63:0] _RAND_178;
  reg [63:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 180:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 316:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 317:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 317:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 249:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 541:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 543:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 182:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 304:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 658:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 658:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 661:91]
  wire [1:0] _T_3069 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 661:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 318:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 271:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 661:113]
  wire [1:0] _T_3070 = _T_3069 & _GEN_465; // @[el2_ifu_mem_ctl.scala 661:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 647:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 661:130]
  wire [1:0] _T_3071 = _T_3070 | _GEN_466; // @[el2_ifu_mem_ctl.scala 661:130]
  wire  _T_3072 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 661:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_3072}; // @[el2_ifu_mem_ctl.scala 661:152]
  wire [1:0] _T_3073 = _T_3071 & _GEN_467; // @[el2_ifu_mem_ctl.scala 661:152]
  wire [1:0] _T_3062 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 661:91]
  wire [1:0] _T_3063 = _T_3062 & _GEN_465; // @[el2_ifu_mem_ctl.scala 661:113]
  wire [1:0] _T_3064 = _T_3063 | _GEN_466; // @[el2_ifu_mem_ctl.scala 661:130]
  wire [1:0] _T_3066 = _T_3064 & _GEN_467; // @[el2_ifu_mem_ctl.scala 661:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3073,_T_3066}; // @[Cat.scala 29:58]
  wire  _T_3173 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3174 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3175 = _T_3173 ^ _T_3174; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3183 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3184 = ^_T_3183; // @[el2_lib.scala 301:83]
  wire  _T_3185 = io_iccm_rd_data_ecc[37] ^ _T_3184; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3192 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3200 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3192}; // @[el2_lib.scala 301:103]
  wire  _T_3201 = ^_T_3200; // @[el2_lib.scala 301:110]
  wire  _T_3202 = io_iccm_rd_data_ecc[36] ^ _T_3201; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3209 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3217 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3209}; // @[el2_lib.scala 301:130]
  wire  _T_3218 = ^_T_3217; // @[el2_lib.scala 301:137]
  wire  _T_3219 = io_iccm_rd_data_ecc[35] ^ _T_3218; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3228 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3237 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3228}; // @[el2_lib.scala 301:157]
  wire  _T_3238 = ^_T_3237; // @[el2_lib.scala 301:164]
  wire  _T_3239 = io_iccm_rd_data_ecc[34] ^ _T_3238; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3248 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3257 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3248}; // @[el2_lib.scala 301:184]
  wire  _T_3258 = ^_T_3257; // @[el2_lib.scala 301:191]
  wire  _T_3259 = io_iccm_rd_data_ecc[33] ^ _T_3258; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3268 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3277 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3268}; // @[el2_lib.scala 301:211]
  wire  _T_3278 = ^_T_3277; // @[el2_lib.scala 301:218]
  wire  _T_3279 = io_iccm_rd_data_ecc[32] ^ _T_3278; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3285 = {_T_3175,_T_3185,_T_3202,_T_3219,_T_3239,_T_3259,_T_3279}; // @[Cat.scala 29:58]
  wire  _T_3286 = _T_3285 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3287 = iccm_ecc_word_enable[0] & _T_3286; // @[el2_lib.scala 302:32]
  wire  _T_3289 = _T_3287 & _T_3285[6]; // @[el2_lib.scala 302:53]
  wire  _T_3558 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3559 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3560 = _T_3558 ^ _T_3559; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3568 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3569 = ^_T_3568; // @[el2_lib.scala 301:83]
  wire  _T_3570 = io_iccm_rd_data_ecc[76] ^ _T_3569; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3577 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3585 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3577}; // @[el2_lib.scala 301:103]
  wire  _T_3586 = ^_T_3585; // @[el2_lib.scala 301:110]
  wire  _T_3587 = io_iccm_rd_data_ecc[75] ^ _T_3586; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3594 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3602 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3594}; // @[el2_lib.scala 301:130]
  wire  _T_3603 = ^_T_3602; // @[el2_lib.scala 301:137]
  wire  _T_3604 = io_iccm_rd_data_ecc[74] ^ _T_3603; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3613 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3622 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3613}; // @[el2_lib.scala 301:157]
  wire  _T_3623 = ^_T_3622; // @[el2_lib.scala 301:164]
  wire  _T_3624 = io_iccm_rd_data_ecc[73] ^ _T_3623; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3633 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3642 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3633}; // @[el2_lib.scala 301:184]
  wire  _T_3643 = ^_T_3642; // @[el2_lib.scala 301:191]
  wire  _T_3644 = io_iccm_rd_data_ecc[72] ^ _T_3643; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3653 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3662 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3653}; // @[el2_lib.scala 301:211]
  wire  _T_3663 = ^_T_3662; // @[el2_lib.scala 301:218]
  wire  _T_3664 = io_iccm_rd_data_ecc[71] ^ _T_3663; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3670 = {_T_3560,_T_3570,_T_3587,_T_3604,_T_3624,_T_3644,_T_3664}; // @[Cat.scala 29:58]
  wire  _T_3671 = _T_3670 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3672 = iccm_ecc_word_enable[1] & _T_3671; // @[el2_lib.scala 302:32]
  wire  _T_3674 = _T_3672 & _T_3670[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3289,_T_3674}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 185:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 625:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 186:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 187:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 470:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 187:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 187:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 187:72]
  wire  _T_2438 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2443 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2463 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 520:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 386:42]
  wire  _T_2465 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 520:79]
  wire  _T_2466 = _T_2463 | _T_2465; // @[el2_ifu_mem_ctl.scala 520:56]
  wire  _T_2467 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 520:122]
  wire  _T_2468 = ~_T_2467; // @[el2_ifu_mem_ctl.scala 520:101]
  wire  _T_2469 = _T_2466 & _T_2468; // @[el2_ifu_mem_ctl.scala 520:99]
  wire  _T_2470 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2484 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 527:45]
  wire  _T_2485 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 527:69]
  wire  _T_2486 = _T_2484 & _T_2485; // @[el2_ifu_mem_ctl.scala 527:67]
  wire  _T_2487 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_2470 ? _T_2486 : _T_2487; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2443 ? _T_2469 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2438 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 187:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 189:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 189:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 279:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 279:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 693:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 279:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 270:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 270:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 320:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 270:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 270:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 279:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 279:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 279:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 279:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 540:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 582:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 609:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 306:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 590:56]
  wire  _T_2589 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 607:69]
  wire  _T_2590 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 607:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2589 : _T_2590; // @[el2_ifu_mem_ctl.scala 607:28]
  wire  _T_2536 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 586:68]
  wire  _T_2537 = ic_act_miss_f | _T_2536; // @[el2_ifu_mem_ctl.scala 586:48]
  wire  bus_reset_data_beat_cnt = _T_2537 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 586:91]
  wire  _T_2533 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 585:50]
  wire  _T_2534 = bus_ifu_wr_en_ff & _T_2533; // @[el2_ifu_mem_ctl.scala 585:48]
  wire  _T_2535 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 585:72]
  wire  bus_inc_data_beat_cnt = _T_2534 & _T_2535; // @[el2_ifu_mem_ctl.scala 585:70]
  wire [2:0] _T_2541 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 589:115]
  wire [2:0] _T_2543 = bus_inc_data_beat_cnt ? _T_2541 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2538 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 587:32]
  wire  _T_2539 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 587:57]
  wire  bus_hold_data_beat_cnt = _T_2538 & _T_2539; // @[el2_ifu_mem_ctl.scala 587:55]
  wire [2:0] _T_2544 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2543 | _T_2544; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 189:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 189:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 190:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 189:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 190:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 196:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 196:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 422:45]
  wire  _T_2108 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 443:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 399:60]
  wire  _T_2139 = _T_2108 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2112 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 443:127]
  wire  _T_2140 = _T_2112 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2147 = _T_2139 | _T_2140; // @[Mux.scala 27:72]
  wire  _T_2116 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 443:127]
  wire  _T_2141 = _T_2116 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2148 = _T_2147 | _T_2141; // @[Mux.scala 27:72]
  wire  _T_2120 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 443:127]
  wire  _T_2142 = _T_2120 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2149 = _T_2148 | _T_2142; // @[Mux.scala 27:72]
  wire  _T_2124 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 443:127]
  wire  _T_2143 = _T_2124 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2150 = _T_2149 | _T_2143; // @[Mux.scala 27:72]
  wire  _T_2128 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 443:127]
  wire  _T_2144 = _T_2128 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2151 = _T_2150 | _T_2144; // @[Mux.scala 27:72]
  wire  _T_2132 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 443:127]
  wire  _T_2145 = _T_2132 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2152 = _T_2151 | _T_2145; // @[Mux.scala 27:72]
  wire  _T_2136 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 443:127]
  wire  _T_2146 = _T_2136 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2152 | _T_2146; // @[Mux.scala 27:72]
  wire  _T_2194 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 445:69]
  wire  _T_2195 = ic_miss_buff_data_valid_bypass_index & _T_2194; // @[el2_ifu_mem_ctl.scala 445:67]
  wire  _T_2197 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 445:91]
  wire  _T_2198 = _T_2195 & _T_2197; // @[el2_ifu_mem_ctl.scala 445:89]
  wire  _T_2203 = _T_2195 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 446:65]
  wire  _T_2204 = _T_2198 | _T_2203; // @[el2_ifu_mem_ctl.scala 445:112]
  wire  _T_2206 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 447:43]
  wire  _T_2209 = _T_2206 & _T_2197; // @[el2_ifu_mem_ctl.scala 447:65]
  wire  _T_2210 = _T_2204 | _T_2209; // @[el2_ifu_mem_ctl.scala 446:88]
  wire  _T_2214 = _T_2206 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 448:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 425:75]
  wire  _T_2154 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2178 = _T_2154 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2157 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2179 = _T_2157 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2186 = _T_2178 | _T_2179; // @[Mux.scala 27:72]
  wire  _T_2160 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2180 = _T_2160 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2187 = _T_2186 | _T_2180; // @[Mux.scala 27:72]
  wire  _T_2163 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2181 = _T_2163 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2188 = _T_2187 | _T_2181; // @[Mux.scala 27:72]
  wire  _T_2166 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2182 = _T_2166 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2189 = _T_2188 | _T_2182; // @[Mux.scala 27:72]
  wire  _T_2169 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2183 = _T_2169 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2190 = _T_2189 | _T_2183; // @[Mux.scala 27:72]
  wire  _T_2172 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2184 = _T_2172 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2191 = _T_2190 | _T_2184; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 444:110]
  wire  _T_2185 = _T_2175 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2191 | _T_2185; // @[Mux.scala 27:72]
  wire  _T_2215 = _T_2214 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 448:87]
  wire  _T_2216 = _T_2210 | _T_2215; // @[el2_ifu_mem_ctl.scala 447:88]
  wire  _T_2220 = ic_miss_buff_data_valid_bypass_index & _T_2136; // @[el2_ifu_mem_ctl.scala 449:43]
  wire  miss_buff_hit_unq_f = _T_2216 | _T_2220; // @[el2_ifu_mem_ctl.scala 448:131]
  wire  _T_2236 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 454:55]
  wire  _T_2237 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 454:87]
  wire  _T_2238 = _T_2236 | _T_2237; // @[el2_ifu_mem_ctl.scala 454:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2238; // @[el2_ifu_mem_ctl.scala 454:41]
  wire  _T_2221 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 451:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 307:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 442:51]
  wire  _T_2222 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 451:68]
  wire  _T_2223 = miss_buff_hit_unq_f & _T_2222; // @[el2_ifu_mem_ctl.scala 451:66]
  wire  stream_hit_f = _T_2221 & _T_2223; // @[el2_ifu_mem_ctl.scala 451:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 274:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 274:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 274:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 592:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 619:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 200:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 200:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 200:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 200:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 200:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 201:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 201:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 202:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 202:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 202:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 202:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 203:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 204:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 204:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 204:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 192:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 204:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 204:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 204:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 205:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 205:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 205:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 205:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 206:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 207:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 207:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 207:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 206:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 205:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 204:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 203:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 202:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 201:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 200:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2233 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 453:60]
  wire  _T_2234 = _T_2233 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 453:92]
  wire  stream_eol_f = _T_2234 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 453:110]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 215:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 215:87]
  wire  _T_113 = _T_111 & _T_2535; // @[el2_ifu_mem_ctl.scala 215:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 215:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 219:48]
  wire  _T_126 = _T_124 & _T_2535; // @[el2_ifu_mem_ctl.scala 219:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 219:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 280:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 280:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 280:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 280:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 280:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 281:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 280:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 281:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 334:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 281:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 281:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 281:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 223:50]
  wire  _T_137 = _T_135 & _T_2535; // @[el2_ifu_mem_ctl.scala 223:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 282:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 283:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 283:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 282:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 224:35]
  wire  _T_143 = _T_141 & _T_2535; // @[el2_ifu_mem_ctl.scala 224:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 223:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 228:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 233:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 190:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 190:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 190:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 190:91]
  wire  _T_30 = ic_act_miss_f & _T_2535; // @[el2_ifu_mem_ctl.scala 197:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 208:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 208:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 208:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 208:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 208:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 208:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 212:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 212:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 212:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 216:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 216:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 220:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 220:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 225:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 225:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 250:95]
  wire  _T_175 = _T_2236 & _T_174; // @[el2_ifu_mem_ctl.scala 250:93]
  wire  crit_wd_byp_ok_ff = _T_2237 | _T_175; // @[el2_ifu_mem_ctl.scala 250:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 251:36]
  wire  _T_180 = _T_2236 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 251:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 251:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 251:70]
  wire  _T_184 = _T_2236 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 252:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 252:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 251:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 252:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 253:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 253:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 252:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 255:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 255:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 263:35]
  reg [6:0] _T_5114; // @[el2_ifu_mem_ctl.scala 721:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_5114[5:0]; // @[el2_ifu_mem_ctl.scala 720:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 717:121]
  wire  _T_4979 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4981 = _T_4979 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4470; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_4470[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4982 = _T_4981 & _GEN_473; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4975 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4977 = _T_4975 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4466; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_4466[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4978 = _T_4977 & _GEN_475; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4971 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4973 = _T_4971 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4462; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_4462[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4974 = _T_4973 & _GEN_477; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4967 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4969 = _T_4967 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4458; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_4458[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4970 = _T_4969 & _GEN_479; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4963 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4965 = _T_4963 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4454; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_4454[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4966 = _T_4965 & _GEN_481; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4959 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4961 = _T_4959 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4450; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_4450[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4962 = _T_4961 & _GEN_483; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4955 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4957 = _T_4955 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4446; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_4446[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4958 = _T_4957 & _GEN_485; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4951 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4953 = _T_4951 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4442; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_4442[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4954 = _T_4953 & _GEN_487; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4947 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4949 = _T_4947 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4438; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_4438[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4950 = _T_4949 & _GEN_489; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4943 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4945 = _T_4943 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4434; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_4434[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4946 = _T_4945 & _GEN_491; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [59:0] _T_4991 = {_T_4982,_T_4978,_T_4974,_T_4970,_T_4966,_T_4962,_T_4958,_T_4954,_T_4950,_T_4946}; // @[Cat.scala 29:58]
  wire  _T_4939 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4941 = _T_4939 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4430; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_4430[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4942 = _T_4941 & _GEN_493; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4935 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4937 = _T_4935 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4426; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_4426[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4938 = _T_4937 & _GEN_495; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4931 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4933 = _T_4931 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4422; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_4422[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4934 = _T_4933 & _GEN_497; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4927 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4929 = _T_4927 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4418; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_4418[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4930 = _T_4929 & _GEN_499; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4923 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4925 = _T_4923 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4414; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_4414[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4926 = _T_4925 & _GEN_501; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4919 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4921 = _T_4919 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4410; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_4410[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4922 = _T_4921 & _GEN_503; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4915 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4917 = _T_4915 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4406; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_4406[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4918 = _T_4917 & _GEN_505; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4911 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4913 = _T_4911 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4402; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_4402[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4914 = _T_4913 & _GEN_507; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4907 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4909 = _T_4907 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4398; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_4398[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4910 = _T_4909 & _GEN_509; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [113:0] _T_5000 = {_T_4991,_T_4942,_T_4938,_T_4934,_T_4930,_T_4926,_T_4922,_T_4918,_T_4914,_T_4910}; // @[Cat.scala 29:58]
  wire  _T_4903 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4905 = _T_4903 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4394; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_4394[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4906 = _T_4905 & _GEN_511; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4899 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4901 = _T_4899 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4390; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_4390[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4902 = _T_4901 & _GEN_513; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4895 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4897 = _T_4895 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4386; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_4386[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4898 = _T_4897 & _GEN_515; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4891 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4893 = _T_4891 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4382; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_4382[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4894 = _T_4893 & _GEN_517; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4887 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4889 = _T_4887 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4378; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_4378[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4890 = _T_4889 & _GEN_519; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4883 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4885 = _T_4883 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4374; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_4374[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4886 = _T_4885 & _GEN_521; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4879 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4881 = _T_4879 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4370; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_4370[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4882 = _T_4881 & _GEN_523; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4875 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4877 = _T_4875 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4366; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_4366[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4878 = _T_4877 & _GEN_525; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4871 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4873 = _T_4871 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4362; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_4362[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4874 = _T_4873 & _GEN_527; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [167:0] _T_5009 = {_T_5000,_T_4906,_T_4902,_T_4898,_T_4894,_T_4890,_T_4886,_T_4882,_T_4878,_T_4874}; // @[Cat.scala 29:58]
  wire  _T_4867 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4869 = _T_4867 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4358; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_4358[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4870 = _T_4869 & _GEN_529; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4863 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4865 = _T_4863 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4354; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_4354[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4866 = _T_4865 & _GEN_531; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4859 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4861 = _T_4859 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4350; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_4350[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4862 = _T_4861 & _GEN_533; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4855 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4857 = _T_4855 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4346; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_4346[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4858 = _T_4857 & _GEN_535; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4851 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4853 = _T_4851 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4342; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_4342[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4854 = _T_4853 & _GEN_537; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4847 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4849 = _T_4847 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4338; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_4338[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4850 = _T_4849 & _GEN_539; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4843 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4845 = _T_4843 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4334; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_4334[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4846 = _T_4845 & _GEN_541; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4839 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4841 = _T_4839 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4330; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_4330[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4842 = _T_4841 & _GEN_543; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4835 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4837 = _T_4835 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4326; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_4326[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4838 = _T_4837 & _GEN_545; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [221:0] _T_5018 = {_T_5009,_T_4870,_T_4866,_T_4862,_T_4858,_T_4854,_T_4850,_T_4846,_T_4842,_T_4838}; // @[Cat.scala 29:58]
  wire  _T_4831 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4833 = _T_4831 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4322; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_4322[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4834 = _T_4833 & _GEN_547; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4827 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4829 = _T_4827 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4318; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_4318[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4830 = _T_4829 & _GEN_549; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4823 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4825 = _T_4823 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4314; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_4314[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4826 = _T_4825 & _GEN_551; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4819 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4821 = _T_4819 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4310; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_4310[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4822 = _T_4821 & _GEN_553; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4815 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4817 = _T_4815 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4306; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_4306[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4818 = _T_4817 & _GEN_555; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4811 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4813 = _T_4811 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4302; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_4302[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4814 = _T_4813 & _GEN_557; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4807 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4809 = _T_4807 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4298; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_4298[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4810 = _T_4809 & _GEN_559; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4803 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4805 = _T_4803 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4294; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_4294[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4806 = _T_4805 & _GEN_561; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4799 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4801 = _T_4799 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4290; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_4290[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4802 = _T_4801 & _GEN_563; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [275:0] _T_5027 = {_T_5018,_T_4834,_T_4830,_T_4826,_T_4822,_T_4818,_T_4814,_T_4810,_T_4806,_T_4802}; // @[Cat.scala 29:58]
  wire  _T_4795 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4797 = _T_4795 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4286; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_4286[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4798 = _T_4797 & _GEN_565; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4791 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4793 = _T_4791 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4282; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_4282[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4794 = _T_4793 & _GEN_567; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4787 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4789 = _T_4787 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4278; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_4278[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4790 = _T_4789 & _GEN_569; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4783 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4785 = _T_4783 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4274; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_4274[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4786 = _T_4785 & _GEN_571; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4779 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4781 = _T_4779 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4270; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_4270[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4782 = _T_4781 & _GEN_573; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4775 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4777 = _T_4775 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4266; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_4266[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4778 = _T_4777 & _GEN_575; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4771 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4773 = _T_4771 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4262; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_4262[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4774 = _T_4773 & _GEN_577; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4767 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4769 = _T_4767 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4258; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_4258[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4770 = _T_4769 & _GEN_579; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4763 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4765 = _T_4763 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4254; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_4254[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4766 = _T_4765 & _GEN_581; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [329:0] _T_5036 = {_T_5027,_T_4798,_T_4794,_T_4790,_T_4786,_T_4782,_T_4778,_T_4774,_T_4770,_T_4766}; // @[Cat.scala 29:58]
  wire  _T_4759 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4761 = _T_4759 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4250; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_4250[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4762 = _T_4761 & _GEN_583; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4755 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4757 = _T_4755 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4246; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_4246[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4758 = _T_4757 & _GEN_585; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4751 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4753 = _T_4751 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4242; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_4242[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4754 = _T_4753 & _GEN_587; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4747 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4749 = _T_4747 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4238; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_4238[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4750 = _T_4749 & _GEN_589; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4743 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4745 = _T_4743 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4234; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_4234[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4746 = _T_4745 & _GEN_591; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4739 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4741 = _T_4739 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4230; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_4230[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4742 = _T_4741 & _GEN_593; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4735 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4737 = _T_4735 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4226; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_4226[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4738 = _T_4737 & _GEN_595; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4731 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4733 = _T_4731 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4222; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_4222[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4734 = _T_4733 & _GEN_597; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4727 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4729 = _T_4727 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4218; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_4218[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4730 = _T_4729 & _GEN_599; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [383:0] _T_5045 = {_T_5036,_T_4762,_T_4758,_T_4754,_T_4750,_T_4746,_T_4742,_T_4738,_T_4734,_T_4730}; // @[Cat.scala 29:58]
  wire  _T_4723 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4725 = _T_4723 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4214; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_4214[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4726 = _T_4725 & _GEN_600; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4719 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4721 = _T_4719 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4210; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_4210[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4722 = _T_4721 & _GEN_601; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4715 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4717 = _T_4715 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4206; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_4206[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4718 = _T_4717 & _GEN_602; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4711 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4713 = _T_4711 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4202; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_4202[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4714 = _T_4713 & _GEN_603; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4707 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4709 = _T_4707 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4198; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_4198[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4710 = _T_4709 & _GEN_604; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4703 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4705 = _T_4703 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4194; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_4194[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4706 = _T_4705 & _GEN_605; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4699 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4701 = _T_4699 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4190; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_4190[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4702 = _T_4701 & _GEN_606; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4695 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4697 = _T_4695 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4186; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_4186[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4698 = _T_4697 & _GEN_607; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4691 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4693 = _T_4691 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4182; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_4182[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4694 = _T_4693 & _GEN_608; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [437:0] _T_5054 = {_T_5045,_T_4726,_T_4722,_T_4718,_T_4714,_T_4710,_T_4706,_T_4702,_T_4698,_T_4694}; // @[Cat.scala 29:58]
  wire  _T_4687 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4689 = _T_4687 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4178; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_4178[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4690 = _T_4689 & _GEN_609; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4683 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4685 = _T_4683 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4174; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_4174[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4686 = _T_4685 & _GEN_610; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4679 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4681 = _T_4679 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4170; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_4170[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4682 = _T_4681 & _GEN_611; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4675 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4677 = _T_4675 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4166; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_4166[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4678 = _T_4677 & _GEN_612; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4671 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4673 = _T_4671 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4162; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_4162[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4674 = _T_4673 & _GEN_613; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4667 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4669 = _T_4667 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4158; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_4158[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4670 = _T_4669 & _GEN_614; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4663 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4665 = _T_4663 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4154; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_4154[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4666 = _T_4665 & _GEN_615; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4659 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4661 = _T_4659 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4150; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_4150[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4662 = _T_4661 & _GEN_616; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4655 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4657 = _T_4655 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4146; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_4146[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4658 = _T_4657 & _GEN_617; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [491:0] _T_5063 = {_T_5054,_T_4690,_T_4686,_T_4682,_T_4678,_T_4674,_T_4670,_T_4666,_T_4662,_T_4658}; // @[Cat.scala 29:58]
  wire  _T_4651 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4653 = _T_4651 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4142; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_4142[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4654 = _T_4653 & _GEN_618; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4647 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4649 = _T_4647 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4138; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_4138[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4650 = _T_4649 & _GEN_619; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4643 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4645 = _T_4643 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4134; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_4134[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4646 = _T_4645 & _GEN_620; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4639 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4641 = _T_4639 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4130; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_4130[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4642 = _T_4641 & _GEN_621; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4635 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4637 = _T_4635 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4126; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_4126[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4638 = _T_4637 & _GEN_622; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4631 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4633 = _T_4631 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4122; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_4122[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4634 = _T_4633 & _GEN_623; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4627 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4629 = _T_4627 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4118; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_4118[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4630 = _T_4629 & _GEN_624; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4623 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4625 = _T_4623 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4114; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_4114[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4626 = _T_4625 & _GEN_625; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4619 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4621 = _T_4619 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4110; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_4110[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4622 = _T_4621 & _GEN_626; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [545:0] _T_5072 = {_T_5063,_T_4654,_T_4650,_T_4646,_T_4642,_T_4638,_T_4634,_T_4630,_T_4626,_T_4622}; // @[Cat.scala 29:58]
  wire  _T_4615 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4617 = _T_4615 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4106; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_4106[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4618 = _T_4617 & _GEN_627; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4611 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4613 = _T_4611 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4102; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_4102[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4614 = _T_4613 & _GEN_628; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4607 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4609 = _T_4607 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4098; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_4098[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4610 = _T_4609 & _GEN_629; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4603 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4605 = _T_4603 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4094; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_4094[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4606 = _T_4605 & _GEN_630; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4599 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4601 = _T_4599 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4090; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_4090[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4602 = _T_4601 & _GEN_631; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4595 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4597 = _T_4595 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4086; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_4086[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4598 = _T_4597 & _GEN_632; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4591 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4593 = _T_4591 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4082; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_4082[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4594 = _T_4593 & _GEN_633; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4587 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4589 = _T_4587 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4078; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_4078[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4590 = _T_4589 & _GEN_634; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4583 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4585 = _T_4583 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4074; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_4074[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4586 = _T_4585 & _GEN_635; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [599:0] _T_5081 = {_T_5072,_T_4618,_T_4614,_T_4610,_T_4606,_T_4602,_T_4598,_T_4594,_T_4590,_T_4586}; // @[Cat.scala 29:58]
  wire  _T_4579 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4581 = _T_4579 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4070; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_4070[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4582 = _T_4581 & _GEN_636; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4575 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4577 = _T_4575 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4066; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_4066[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4578 = _T_4577 & _GEN_637; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4571 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4573 = _T_4571 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4062; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_4062[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4574 = _T_4573 & _GEN_638; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4567 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4569 = _T_4567 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4058; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_4058[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4570 = _T_4569 & _GEN_639; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4563 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4565 = _T_4563 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4054; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_4054[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4566 = _T_4565 & _GEN_640; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4559 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4561 = _T_4559 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4050; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_4050[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4562 = _T_4561 & _GEN_641; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4555 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4557 = _T_4555 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4046; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_4046[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4558 = _T_4557 & _GEN_642; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4551 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4553 = _T_4551 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4042; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_4042[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4554 = _T_4553 & _GEN_643; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4547 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4549 = _T_4547 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4038; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_4038[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4550 = _T_4549 & _GEN_644; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [653:0] _T_5090 = {_T_5081,_T_4582,_T_4578,_T_4574,_T_4570,_T_4566,_T_4562,_T_4558,_T_4554,_T_4550}; // @[Cat.scala 29:58]
  wire  _T_4543 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4545 = _T_4543 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4034; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_4034[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4546 = _T_4545 & _GEN_645; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4539 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4541 = _T_4539 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4030; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_4030[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4542 = _T_4541 & _GEN_646; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4535 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4537 = _T_4535 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4026; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_4026[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4538 = _T_4537 & _GEN_647; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4531 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4533 = _T_4531 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4022; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_4022[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4534 = _T_4533 & _GEN_648; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4527 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4529 = _T_4527 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4018; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_4018[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4530 = _T_4529 & _GEN_649; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4523 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4525 = _T_4523 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4014; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_4014[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4526 = _T_4525 & _GEN_650; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4519 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4521 = _T_4519 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4010; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_4010[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4522 = _T_4521 & _GEN_651; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4515 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4517 = _T_4515 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4006; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_4006[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4518 = _T_4517 & _GEN_652; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4511 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4513 = _T_4511 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4002; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_4002[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4514 = _T_4513 & _GEN_653; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [707:0] _T_5099 = {_T_5090,_T_4546,_T_4542,_T_4538,_T_4534,_T_4530,_T_4526,_T_4522,_T_4518,_T_4514}; // @[Cat.scala 29:58]
  wire  _T_4507 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4509 = _T_4507 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3998; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3998[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4510 = _T_4509 & _GEN_654; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4503 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4505 = _T_4503 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3994; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3994[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4506 = _T_4505 & _GEN_655; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4499 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4501 = _T_4499 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3990; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3990[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4502 = _T_4501 & _GEN_656; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4495 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4497 = _T_4495 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3986; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3986[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4498 = _T_4497 & _GEN_657; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4491 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4493 = _T_4491 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3982; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3982[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4494 = _T_4493 & _GEN_658; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4487 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4489 = _T_4487 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3978; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3978[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4490 = _T_4489 & _GEN_659; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4483 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4485 = _T_4483 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3974; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3974[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4486 = _T_4485 & _GEN_660; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4479 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4481 = _T_4479 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3970; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3970[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4482 = _T_4481 & _GEN_661; // @[el2_ifu_mem_ctl.scala 717:130]
  wire  _T_4475 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4477 = _T_4475 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3966; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3966[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4478 = _T_4477 & _GEN_662; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [761:0] _T_5108 = {_T_5099,_T_4510,_T_4506,_T_4502,_T_4498,_T_4494,_T_4490,_T_4486,_T_4482,_T_4478}; // @[Cat.scala 29:58]
  wire  _T_4471 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 717:121]
  wire [5:0] _T_4473 = _T_4471 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3962; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3962[0]; // @[el2_ifu_mem_ctl.scala 714:30 el2_ifu_mem_ctl.scala 716:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [5:0] _T_4474 = _T_4473 & _GEN_663; // @[el2_ifu_mem_ctl.scala 717:130]
  wire [767:0] _T_5109 = {_T_5108,_T_4474}; // @[Cat.scala 29:58]
  wire  way_status = _T_5109[0]; // @[el2_ifu_mem_ctl.scala 717:16]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 258:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 260:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 262:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 267:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 272:59]
  wire  _T_214 = _T_212 | _T_2221; // @[el2_ifu_mem_ctl.scala 272:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 272:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 278:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 278:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 278:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 278:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 285:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 285:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 285:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 286:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 286:32]
  wire  _T_274 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 289:75]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 289:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2610 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 615:48]
  wire  _T_2611 = _T_2610 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 615:52]
  wire  bus_ifu_wr_data_error_ff = _T_2611 & miss_pending; // @[el2_ifu_mem_ctl.scala 615:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 361:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 360:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 289:145]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 289:143]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 292:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 292:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 293:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 312:30]
  wire  _T_10059 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 770:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 313:24]
  wire  _T_10061 = _T_10059 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 770:51]
  wire  _T_10063 = _T_10061 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 770:67]
  wire  _T_10065 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 770:86]
  wire  replace_way_mb_any_0 = _T_10063 | _T_10065; // @[el2_ifu_mem_ctl.scala 770:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10068 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 771:50]
  wire  _T_10070 = _T_10068 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 771:66]
  wire  _T_10072 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 771:85]
  wire  _T_10074 = _T_10072 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 771:100]
  wire  replace_way_mb_any_1 = _T_10070 | _T_10074; // @[el2_ifu_mem_ctl.scala 771:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 297:110]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 301:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 301:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 302:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 301:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 301:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 303:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 311:23]
  wire  _T_313 = _T_2236 & flush_final_f; // @[el2_ifu_mem_ctl.scala 315:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 315:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 315:53]
  wire  _T_2228 = ~_T_2223; // @[el2_ifu_mem_ctl.scala 452:46]
  wire  _T_2229 = _T_2221 & _T_2228; // @[el2_ifu_mem_ctl.scala 452:44]
  wire  stream_miss_f = _T_2229 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 452:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 315:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 315:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 321:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_2221; // @[el2_ifu_mem_ctl.scala 323:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 323:82]
  wire  _T_2242 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 457:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2242}; // @[Cat.scala 29:58]
  wire  _T_2243 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2267 = _T_2243 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2246 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2268 = _T_2246 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2275 = _T_2267 | _T_2268; // @[Mux.scala 27:72]
  wire  _T_2249 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2269 = _T_2249 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2276 = _T_2275 | _T_2269; // @[Mux.scala 27:72]
  wire  _T_2252 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2270 = _T_2252 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2277 = _T_2276 | _T_2270; // @[Mux.scala 27:72]
  wire  _T_2255 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2271 = _T_2255 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2278 = _T_2277 | _T_2271; // @[Mux.scala 27:72]
  wire  _T_2258 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2272 = _T_2258 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2279 = _T_2278 | _T_2272; // @[Mux.scala 27:72]
  wire  _T_2261 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2273 = _T_2261 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2280 = _T_2279 | _T_2273; // @[Mux.scala 27:72]
  wire  _T_2264 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 458:81]
  wire  _T_2274 = _T_2264 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2280 | _T_2274; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 459:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 327:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 327:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 612:61]
  wire  _T_2604 = ic_act_miss_f_delayed & _T_2237; // @[el2_ifu_mem_ctl.scala 613:53]
  wire  reset_tag_valid_for_miss = _T_2604 & _T_17; // @[el2_ifu_mem_ctl.scala 613:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 327:79]
  wire [30:0] _T_337 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_339 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 329:37]
  wire [30:0] _T_340 = sel_mb_addr ? _T_337 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_341 = _T_339 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_340 | _T_341; // @[Mux.scala 27:72]
  wire  _T_346 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 331:84]
  wire  _T_2598 = ~_T_2610; // @[el2_ifu_mem_ctl.scala 610:84]
  wire  _T_2599 = _T_100 & _T_2598; // @[el2_ifu_mem_ctl.scala 610:82]
  wire  bus_ifu_wr_en_ff_q = _T_2599 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 610:108]
  wire  sel_mb_status_addr = _T_346 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 331:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_337 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 332:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [7:0] _T_570 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_579 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_570}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_587 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_596 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_587}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_597 = {_T_596,_T_579}; // @[el2_lib.scala 348:27]
  wire  _T_598 = ^_T_597; // @[el2_lib.scala 348:34]
  wire [7:0] _T_605 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_614 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_605}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_622 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_631 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_622}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_632 = {_T_631,_T_614}; // @[el2_lib.scala 348:44]
  wire  _T_633 = ^_T_632; // @[el2_lib.scala 348:51]
  wire [7:0] _T_640 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_649 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_640}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_657 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_666 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_657}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_667 = {_T_666,_T_649}; // @[el2_lib.scala 348:61]
  wire  _T_668 = ^_T_667; // @[el2_lib.scala 348:68]
  wire [6:0] _T_674 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_682 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_674}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_689 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_698 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_689,_T_682}; // @[el2_lib.scala 348:78]
  wire  _T_699 = ^_T_698; // @[el2_lib.scala 348:85]
  wire [6:0] _T_705 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_713 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_705}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_720 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_729 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_720,_T_713}; // @[el2_lib.scala 348:95]
  wire  _T_730 = ^_T_729; // @[el2_lib.scala 348:102]
  wire [6:0] _T_736 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_744 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_736}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_760 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_720,_T_744}; // @[el2_lib.scala 348:112]
  wire  _T_761 = ^_T_760; // @[el2_lib.scala 348:119]
  wire [6:0] _T_767 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 348:129]
  wire  _T_768 = ^_T_767; // @[el2_lib.scala 348:136]
  wire [3:0] _T_2283 = {ifu_bus_rid_ff[2:1],_T_2242,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2284 = _T_2283 == 4'h0; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1295; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_0 = _T_1295[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2331 = _T_2284 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2287 = _T_2283 == 4'h1; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1297; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_1 = _T_1297[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2332 = _T_2287 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2347 = _T_2331 | _T_2332; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2283 == 4'h2; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1299; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_2 = _T_1299[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2333 = _T_2290 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2348 = _T_2347 | _T_2333; // @[Mux.scala 27:72]
  wire  _T_2293 = _T_2283 == 4'h3; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1301; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_3 = _T_1301[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2334 = _T_2293 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2349 = _T_2348 | _T_2334; // @[Mux.scala 27:72]
  wire  _T_2296 = _T_2283 == 4'h4; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1303; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_4 = _T_1303[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2335 = _T_2296 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2350 = _T_2349 | _T_2335; // @[Mux.scala 27:72]
  wire  _T_2299 = _T_2283 == 4'h5; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1305; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_5 = _T_1305[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2336 = _T_2299 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2351 = _T_2350 | _T_2336; // @[Mux.scala 27:72]
  wire  _T_2302 = _T_2283 == 4'h6; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1307; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_6 = _T_1307[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2337 = _T_2302 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2352 = _T_2351 | _T_2337; // @[Mux.scala 27:72]
  wire  _T_2305 = _T_2283 == 4'h7; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1309; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_7 = _T_1309[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2338 = _T_2305 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2353 = _T_2352 | _T_2338; // @[Mux.scala 27:72]
  wire  _T_2308 = _T_2283 == 4'h8; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1311; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_8 = _T_1311[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2339 = _T_2308 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2354 = _T_2353 | _T_2339; // @[Mux.scala 27:72]
  wire  _T_2311 = _T_2283 == 4'h9; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1313; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_9 = _T_1313[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2340 = _T_2311 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2355 = _T_2354 | _T_2340; // @[Mux.scala 27:72]
  wire  _T_2314 = _T_2283 == 4'ha; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1315; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_10 = _T_1315[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2341 = _T_2314 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2356 = _T_2355 | _T_2341; // @[Mux.scala 27:72]
  wire  _T_2317 = _T_2283 == 4'hb; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1317; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_11 = _T_1317[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2342 = _T_2317 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2357 = _T_2356 | _T_2342; // @[Mux.scala 27:72]
  wire  _T_2320 = _T_2283 == 4'hc; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1319; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_12 = _T_1319[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2343 = _T_2320 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2358 = _T_2357 | _T_2343; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2283 == 4'hd; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1321; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_13 = _T_1321[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2344 = _T_2323 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2358 | _T_2344; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2283 == 4'he; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1323; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_14 = _T_1323[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 395:26]
  wire [31:0] _T_2345 = _T_2326 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2360 = _T_2359 | _T_2345; // @[Mux.scala 27:72]
  wire  _T_2329 = _T_2283 == 4'hf; // @[el2_ifu_mem_ctl.scala 460:89]
  reg [63:0] _T_1325; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_15 = _T_1325[31:0]; // @[el2_ifu_mem_ctl.scala 393:31 el2_ifu_mem_ctl.scala 396:28]
  wire [31:0] _T_2346 = _T_2329 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2360 | _T_2346; // @[Mux.scala 27:72]
  wire [3:0] _T_2363 = {ifu_bus_rid_ff[2:1],_T_2242,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2364 = _T_2363 == 4'h0; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2387 = _T_2364 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2367 = _T_2363 == 4'h1; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2388 = _T_2367 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2395 = _T_2387 | _T_2388; // @[Mux.scala 27:72]
  wire  _T_2370 = _T_2363 == 4'h2; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2389 = _T_2370 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2396 = _T_2395 | _T_2389; // @[Mux.scala 27:72]
  wire  _T_2373 = _T_2363 == 4'h3; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2390 = _T_2373 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2397 = _T_2396 | _T_2390; // @[Mux.scala 27:72]
  wire  _T_2376 = _T_2363 == 4'h4; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2391 = _T_2376 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2398 = _T_2397 | _T_2391; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2363 == 4'h5; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2392 = _T_2379 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2399 = _T_2398 | _T_2392; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2363 == 4'h6; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2393 = _T_2382 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2400 = _T_2399 | _T_2393; // @[Mux.scala 27:72]
  wire  _T_2385 = _T_2363 == 4'h7; // @[el2_ifu_mem_ctl.scala 461:64]
  wire [31:0] _T_2394 = _T_2385 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2401 = _T_2400 | _T_2394; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2361,_T_2401}; // @[Cat.scala 29:58]
  wire [7:0] _T_992 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_1001 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_992}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_1009 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_1018 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1009}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_1019 = {_T_1018,_T_1001}; // @[el2_lib.scala 348:27]
  wire  _T_1020 = ^_T_1019; // @[el2_lib.scala 348:34]
  wire [7:0] _T_1027 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_1036 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1027}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_1044 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_1053 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1044}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_1054 = {_T_1053,_T_1036}; // @[el2_lib.scala 348:44]
  wire  _T_1055 = ^_T_1054; // @[el2_lib.scala 348:51]
  wire [7:0] _T_1062 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_1071 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1062}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_1079 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_1088 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1079}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_1089 = {_T_1088,_T_1071}; // @[el2_lib.scala 348:61]
  wire  _T_1090 = ^_T_1089; // @[el2_lib.scala 348:68]
  wire [6:0] _T_1096 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_1104 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1096}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_1111 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_1120 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1111,_T_1104}; // @[el2_lib.scala 348:78]
  wire  _T_1121 = ^_T_1120; // @[el2_lib.scala 348:85]
  wire [6:0] _T_1127 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_1135 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1127}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_1142 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_1151 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1142,_T_1135}; // @[el2_lib.scala 348:95]
  wire  _T_1152 = ^_T_1151; // @[el2_lib.scala 348:102]
  wire [6:0] _T_1158 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_1166 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_1158}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_1182 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1142,_T_1166}; // @[el2_lib.scala 348:112]
  wire  _T_1183 = ^_T_1182; // @[el2_lib.scala 348:119]
  wire [6:0] _T_1189 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 348:129]
  wire  _T_1190 = ^_T_1189; // @[el2_lib.scala 348:136]
  wire [70:0] _T_1237 = {_T_598,_T_633,_T_668,_T_699,_T_730,_T_761,_T_768,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1236 = {_T_1020,_T_1055,_T_1090,_T_1121,_T_1152,_T_1183,_T_1190,_T_2361,_T_2401}; // @[Cat.scala 29:58]
  wire [141:0] _T_1238 = {_T_598,_T_633,_T_668,_T_699,_T_730,_T_761,_T_768,ifu_bus_rdata_ff,_T_1236}; // @[Cat.scala 29:58]
  wire [141:0] _T_1241 = {_T_1020,_T_1055,_T_1090,_T_1121,_T_1152,_T_1183,_T_1190,_T_2361,_T_2401,_T_1237}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1238 : _T_1241; // @[el2_ifu_mem_ctl.scala 353:28]
  wire  _T_1198 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 343:56]
  wire  _T_1199 = _T_1198 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 343:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 407:28]
  wire  _T_1401 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 608:35]
  wire  _T_1286 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1327 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 398:118]
  wire  _T_1328 = ic_miss_buff_data_valid[0] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1328; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1424 = _T_1401 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1404 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1331 = ic_miss_buff_data_valid[1] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1331; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1425 = _T_1404 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1432 = _T_1424 | _T_1425; // @[Mux.scala 27:72]
  wire  _T_1407 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1334 = ic_miss_buff_data_valid[2] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1334; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1426 = _T_1407 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1433 = _T_1432 | _T_1426; // @[Mux.scala 27:72]
  wire  _T_1410 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1337 = ic_miss_buff_data_valid[3] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1337; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1427 = _T_1410 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1434 = _T_1433 | _T_1427; // @[Mux.scala 27:72]
  wire  _T_1413 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  _T_1290 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1290; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1340 = ic_miss_buff_data_valid[4] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1340; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1428 = _T_1413 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1435 = _T_1434 | _T_1428; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  _T_1291 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1291; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1343 = ic_miss_buff_data_valid[5] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1343; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1429 = _T_1416 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1436 = _T_1435 | _T_1429; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  _T_1292 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1292; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1346 = ic_miss_buff_data_valid[6] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1346; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1430 = _T_1419 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1437 = _T_1436 | _T_1430; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 409:114]
  wire  _T_1293 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 392:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1293; // @[el2_ifu_mem_ctl.scala 392:73]
  wire  _T_1349 = ic_miss_buff_data_valid[7] & _T_1327; // @[el2_ifu_mem_ctl.scala 398:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1349; // @[el2_ifu_mem_ctl.scala 398:88]
  wire  _T_1431 = _T_1422 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1437 | _T_1431; // @[Mux.scala 27:72]
  wire  _T_1440 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 410:58]
  wire  _T_1441 = bypass_valid_value_check & _T_1440; // @[el2_ifu_mem_ctl.scala 410:56]
  wire  _T_1443 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 410:77]
  wire  _T_1444 = _T_1441 & _T_1443; // @[el2_ifu_mem_ctl.scala 410:75]
  wire  _T_1449 = _T_1441 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 411:75]
  wire  _T_1450 = _T_1444 | _T_1449; // @[el2_ifu_mem_ctl.scala 410:95]
  wire  _T_1452 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 412:56]
  wire  _T_1455 = _T_1452 & _T_1443; // @[el2_ifu_mem_ctl.scala 412:74]
  wire  _T_1456 = _T_1450 | _T_1455; // @[el2_ifu_mem_ctl.scala 411:94]
  wire  _T_1460 = _T_1452 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 413:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 408:70]
  wire  _T_1461 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1477 = _T_1461 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1463 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1478 = _T_1463 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1485 = _T_1477 | _T_1478; // @[Mux.scala 27:72]
  wire  _T_1465 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1479 = _T_1465 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1486 = _T_1485 | _T_1479; // @[Mux.scala 27:72]
  wire  _T_1467 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1480 = _T_1467 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1487 = _T_1486 | _T_1480; // @[Mux.scala 27:72]
  wire  _T_1469 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1481 = _T_1469 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1487 | _T_1481; // @[Mux.scala 27:72]
  wire  _T_1471 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1482 = _T_1471 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1488 | _T_1482; // @[Mux.scala 27:72]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1483 = _T_1473 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1490 = _T_1489 | _T_1483; // @[Mux.scala 27:72]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 413:132]
  wire  _T_1484 = _T_1475 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1490 | _T_1484; // @[Mux.scala 27:72]
  wire  _T_1493 = _T_1460 & _T_1491; // @[el2_ifu_mem_ctl.scala 413:69]
  wire  _T_1494 = _T_1456 | _T_1493; // @[el2_ifu_mem_ctl.scala 412:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 414:95]
  wire  _T_1497 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 414:95]
  wire  _T_1498 = bypass_valid_value_check & _T_1497; // @[el2_ifu_mem_ctl.scala 414:56]
  wire  bypass_data_ready_in = _T_1494 | _T_1498; // @[el2_ifu_mem_ctl.scala 413:181]
  wire  _T_1499 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 418:53]
  wire  _T_1500 = _T_1499 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 418:73]
  wire  _T_1502 = _T_1500 & _T_317; // @[el2_ifu_mem_ctl.scala 418:96]
  wire  _T_1504 = _T_1502 & _T_58; // @[el2_ifu_mem_ctl.scala 418:118]
  wire  _T_1506 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 419:73]
  wire  _T_1508 = _T_1506 & _T_317; // @[el2_ifu_mem_ctl.scala 419:96]
  wire  _T_1510 = _T_1508 & _T_58; // @[el2_ifu_mem_ctl.scala 419:118]
  wire  _T_1511 = _T_1504 | _T_1510; // @[el2_ifu_mem_ctl.scala 418:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 421:58]
  wire  _T_1512 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 420:54]
  wire  _T_1513 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 420:76]
  wire  _T_1514 = _T_1512 & _T_1513; // @[el2_ifu_mem_ctl.scala 420:74]
  wire  _T_1516 = _T_1514 & _T_317; // @[el2_ifu_mem_ctl.scala 420:96]
  wire  ic_crit_wd_rdy_new_in = _T_1511 | _T_1516; // @[el2_ifu_mem_ctl.scala 419:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 618:43]
  wire  _T_1253 = ic_crit_wd_rdy | _T_2221; // @[el2_ifu_mem_ctl.scala 365:38]
  wire  _T_1255 = _T_1253 | _T_2237; // @[el2_ifu_mem_ctl.scala 365:64]
  wire  _T_1256 = ~_T_1255; // @[el2_ifu_mem_ctl.scala 365:21]
  wire  _T_1257 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 365:98]
  wire  sel_ic_data = _T_1256 & _T_1257; // @[el2_ifu_mem_ctl.scala 365:96]
  wire  _T_2404 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 463:44]
  wire  _T_1610 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 432:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 404:60]
  wire  _T_1554 = _T_1401 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1404 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1562 = _T_1554 | _T_1555; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1407 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1563 = _T_1562 | _T_1556; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1410 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1564 = _T_1563 | _T_1557; // @[Mux.scala 27:72]
  wire  _T_1558 = _T_1413 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1565 = _T_1564 | _T_1558; // @[Mux.scala 27:72]
  wire  _T_1559 = _T_1416 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1566 = _T_1565 | _T_1559; // @[Mux.scala 27:72]
  wire  _T_1560 = _T_1419 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1566 | _T_1560; // @[Mux.scala 27:72]
  wire  _T_1561 = _T_1422 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1567 | _T_1561; // @[Mux.scala 27:72]
  wire  _T_1593 = _T_2154 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1594 = _T_2157 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1601 = _T_1593 | _T_1594; // @[Mux.scala 27:72]
  wire  _T_1595 = _T_2160 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1602 = _T_1601 | _T_1595; // @[Mux.scala 27:72]
  wire  _T_1596 = _T_2163 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1603 = _T_1602 | _T_1596; // @[Mux.scala 27:72]
  wire  _T_1597 = _T_2166 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1604 = _T_1603 | _T_1597; // @[Mux.scala 27:72]
  wire  _T_1598 = _T_2169 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1605 = _T_1604 | _T_1598; // @[Mux.scala 27:72]
  wire  _T_1599 = _T_2172 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1606 = _T_1605 | _T_1599; // @[Mux.scala 27:72]
  wire  _T_1600 = _T_2175 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1606 | _T_1600; // @[Mux.scala 27:72]
  wire  _T_1611 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 434:70]
  wire  ifu_byp_data_err_new = _T_1610 ? ic_miss_buff_data_error_bypass : _T_1611; // @[el2_ifu_mem_ctl.scala 432:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 376:42]
  wire  _T_2405 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 463:91]
  wire  _T_2406 = ~_T_2405; // @[el2_ifu_mem_ctl.scala 463:60]
  wire  ic_rd_parity_final_err = _T_2404 & _T_2406; // @[el2_ifu_mem_ctl.scala 463:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9677 = _T_4471 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 745:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9679 = _T_4475 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9932 = _T_9677 | _T_9679; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9681 = _T_4479 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9933 = _T_9932 | _T_9681; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9683 = _T_4483 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9934 = _T_9933 | _T_9683; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9685 = _T_4487 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9935 = _T_9934 | _T_9685; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9687 = _T_4491 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9936 = _T_9935 | _T_9687; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9689 = _T_4495 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9937 = _T_9936 | _T_9689; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9691 = _T_4499 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9938 = _T_9937 | _T_9691; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9693 = _T_4503 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9939 = _T_9938 | _T_9693; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9695 = _T_4507 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9940 = _T_9939 | _T_9695; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9697 = _T_4511 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9941 = _T_9940 | _T_9697; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9699 = _T_4515 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9942 = _T_9941 | _T_9699; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9701 = _T_4519 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9943 = _T_9942 | _T_9701; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9703 = _T_4523 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9944 = _T_9943 | _T_9703; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9705 = _T_4527 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9945 = _T_9944 | _T_9705; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9707 = _T_4531 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9946 = _T_9945 | _T_9707; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9709 = _T_4535 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9947 = _T_9946 | _T_9709; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9711 = _T_4539 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9948 = _T_9947 | _T_9711; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9713 = _T_4543 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9949 = _T_9948 | _T_9713; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9715 = _T_4547 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9950 = _T_9949 | _T_9715; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9717 = _T_4551 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9951 = _T_9950 | _T_9717; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9719 = _T_4555 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9952 = _T_9951 | _T_9719; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9721 = _T_4559 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9953 = _T_9952 | _T_9721; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9723 = _T_4563 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9954 = _T_9953 | _T_9723; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9725 = _T_4567 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9955 = _T_9954 | _T_9725; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9727 = _T_4571 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9956 = _T_9955 | _T_9727; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9729 = _T_4575 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9957 = _T_9956 | _T_9729; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9731 = _T_4579 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9958 = _T_9957 | _T_9731; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9733 = _T_4583 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9959 = _T_9958 | _T_9733; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9735 = _T_4587 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9960 = _T_9959 | _T_9735; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9737 = _T_4591 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9961 = _T_9960 | _T_9737; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9739 = _T_4595 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9962 = _T_9961 | _T_9739; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9741 = _T_4599 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9963 = _T_9962 | _T_9741; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9743 = _T_4603 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9964 = _T_9963 | _T_9743; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9745 = _T_4607 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9965 = _T_9964 | _T_9745; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9747 = _T_4611 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9966 = _T_9965 | _T_9747; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9749 = _T_4615 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9967 = _T_9966 | _T_9749; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9751 = _T_4619 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9968 = _T_9967 | _T_9751; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9753 = _T_4623 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9969 = _T_9968 | _T_9753; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9755 = _T_4627 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9970 = _T_9969 | _T_9755; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9757 = _T_4631 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9971 = _T_9970 | _T_9757; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9759 = _T_4635 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9972 = _T_9971 | _T_9759; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9761 = _T_4639 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9973 = _T_9972 | _T_9761; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9763 = _T_4643 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9974 = _T_9973 | _T_9763; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9765 = _T_4647 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9975 = _T_9974 | _T_9765; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9767 = _T_4651 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9976 = _T_9975 | _T_9767; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9769 = _T_4655 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9977 = _T_9976 | _T_9769; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9771 = _T_4659 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9978 = _T_9977 | _T_9771; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9773 = _T_4663 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9979 = _T_9978 | _T_9773; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9775 = _T_4667 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9980 = _T_9979 | _T_9775; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9777 = _T_4671 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9981 = _T_9980 | _T_9777; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9779 = _T_4675 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9982 = _T_9981 | _T_9779; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9781 = _T_4679 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9983 = _T_9982 | _T_9781; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9783 = _T_4683 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9984 = _T_9983 | _T_9783; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9785 = _T_4687 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9985 = _T_9984 | _T_9785; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9787 = _T_4691 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9986 = _T_9985 | _T_9787; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9789 = _T_4695 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9987 = _T_9986 | _T_9789; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9791 = _T_4699 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9988 = _T_9987 | _T_9791; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9793 = _T_4703 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9989 = _T_9988 | _T_9793; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9795 = _T_4707 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9990 = _T_9989 | _T_9795; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9797 = _T_4711 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9991 = _T_9990 | _T_9797; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9799 = _T_4715 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9992 = _T_9991 | _T_9799; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9801 = _T_4719 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9993 = _T_9992 | _T_9801; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9803 = _T_4723 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9994 = _T_9993 | _T_9803; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9805 = _T_4727 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9995 = _T_9994 | _T_9805; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9807 = _T_4731 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9996 = _T_9995 | _T_9807; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9809 = _T_4735 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9997 = _T_9996 | _T_9809; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9811 = _T_4739 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9998 = _T_9997 | _T_9811; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9813 = _T_4743 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9999 = _T_9998 | _T_9813; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9815 = _T_4747 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10000 = _T_9999 | _T_9815; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9817 = _T_4751 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10001 = _T_10000 | _T_9817; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9819 = _T_4755 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10002 = _T_10001 | _T_9819; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9821 = _T_4759 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10003 = _T_10002 | _T_9821; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9823 = _T_4763 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10004 = _T_10003 | _T_9823; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9825 = _T_4767 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10005 = _T_10004 | _T_9825; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9827 = _T_4771 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10006 = _T_10005 | _T_9827; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9829 = _T_4775 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10007 = _T_10006 | _T_9829; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9831 = _T_4779 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10008 = _T_10007 | _T_9831; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9833 = _T_4783 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10009 = _T_10008 | _T_9833; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9835 = _T_4787 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10010 = _T_10009 | _T_9835; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9837 = _T_4791 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10011 = _T_10010 | _T_9837; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9839 = _T_4795 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10012 = _T_10011 | _T_9839; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9841 = _T_4799 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10013 = _T_10012 | _T_9841; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9843 = _T_4803 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10014 = _T_10013 | _T_9843; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9845 = _T_4807 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10015 = _T_10014 | _T_9845; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9847 = _T_4811 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10016 = _T_10015 | _T_9847; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9849 = _T_4815 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10017 = _T_10016 | _T_9849; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9851 = _T_4819 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10018 = _T_10017 | _T_9851; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9853 = _T_4823 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10019 = _T_10018 | _T_9853; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9855 = _T_4827 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10020 = _T_10019 | _T_9855; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9857 = _T_4831 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10021 = _T_10020 | _T_9857; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9859 = _T_4835 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10022 = _T_10021 | _T_9859; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9861 = _T_4839 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10023 = _T_10022 | _T_9861; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9863 = _T_4843 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10024 = _T_10023 | _T_9863; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9865 = _T_4847 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10025 = _T_10024 | _T_9865; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9867 = _T_4851 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10026 = _T_10025 | _T_9867; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9869 = _T_4855 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10027 = _T_10026 | _T_9869; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9871 = _T_4859 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10028 = _T_10027 | _T_9871; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9873 = _T_4863 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10029 = _T_10028 | _T_9873; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9875 = _T_4867 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10030 = _T_10029 | _T_9875; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9877 = _T_4871 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10031 = _T_10030 | _T_9877; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9879 = _T_4875 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10032 = _T_10031 | _T_9879; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9881 = _T_4879 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10033 = _T_10032 | _T_9881; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9883 = _T_4883 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10034 = _T_10033 | _T_9883; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9885 = _T_4887 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10035 = _T_10034 | _T_9885; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9887 = _T_4891 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10036 = _T_10035 | _T_9887; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9889 = _T_4895 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10037 = _T_10036 | _T_9889; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9891 = _T_4899 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10038 = _T_10037 | _T_9891; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9893 = _T_4903 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10039 = _T_10038 | _T_9893; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9895 = _T_4907 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10040 = _T_10039 | _T_9895; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9897 = _T_4911 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10041 = _T_10040 | _T_9897; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9899 = _T_4915 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10042 = _T_10041 | _T_9899; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9901 = _T_4919 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10043 = _T_10042 | _T_9901; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9903 = _T_4923 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10044 = _T_10043 | _T_9903; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9905 = _T_4927 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10045 = _T_10044 | _T_9905; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9907 = _T_4931 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10046 = _T_10045 | _T_9907; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9909 = _T_4935 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10047 = _T_10046 | _T_9909; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9911 = _T_4939 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10048 = _T_10047 | _T_9911; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9913 = _T_4943 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10049 = _T_10048 | _T_9913; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9915 = _T_4947 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10050 = _T_10049 | _T_9915; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9917 = _T_4951 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10051 = _T_10050 | _T_9917; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9919 = _T_4955 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10052 = _T_10051 | _T_9919; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9921 = _T_4959 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10053 = _T_10052 | _T_9921; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9923 = _T_4963 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10054 = _T_10053 | _T_9923; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9925 = _T_4967 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10055 = _T_10054 | _T_9925; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9927 = _T_4971 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10056 = _T_10055 | _T_9927; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9929 = _T_4975 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10057 = _T_10056 | _T_9929; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9931 = _T_4979 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_10058 = _T_10057 | _T_9931; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9294 = _T_4471 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 745:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9296 = _T_4475 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9549 = _T_9294 | _T_9296; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9298 = _T_4479 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9550 = _T_9549 | _T_9298; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9300 = _T_4483 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9551 = _T_9550 | _T_9300; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9302 = _T_4487 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9552 = _T_9551 | _T_9302; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9304 = _T_4491 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9553 = _T_9552 | _T_9304; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9306 = _T_4495 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9554 = _T_9553 | _T_9306; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9308 = _T_4499 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9555 = _T_9554 | _T_9308; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9310 = _T_4503 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9556 = _T_9555 | _T_9310; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9312 = _T_4507 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9557 = _T_9556 | _T_9312; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9314 = _T_4511 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9558 = _T_9557 | _T_9314; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9316 = _T_4515 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9559 = _T_9558 | _T_9316; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9318 = _T_4519 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9560 = _T_9559 | _T_9318; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9320 = _T_4523 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9561 = _T_9560 | _T_9320; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9322 = _T_4527 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9562 = _T_9561 | _T_9322; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9324 = _T_4531 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9563 = _T_9562 | _T_9324; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9326 = _T_4535 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9564 = _T_9563 | _T_9326; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9328 = _T_4539 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9565 = _T_9564 | _T_9328; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9330 = _T_4543 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9566 = _T_9565 | _T_9330; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9332 = _T_4547 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9567 = _T_9566 | _T_9332; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9334 = _T_4551 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9568 = _T_9567 | _T_9334; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9336 = _T_4555 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9569 = _T_9568 | _T_9336; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9338 = _T_4559 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9570 = _T_9569 | _T_9338; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9340 = _T_4563 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9571 = _T_9570 | _T_9340; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9342 = _T_4567 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9572 = _T_9571 | _T_9342; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9344 = _T_4571 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9573 = _T_9572 | _T_9344; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9346 = _T_4575 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9574 = _T_9573 | _T_9346; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9348 = _T_4579 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9575 = _T_9574 | _T_9348; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9350 = _T_4583 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9576 = _T_9575 | _T_9350; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9352 = _T_4587 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9577 = _T_9576 | _T_9352; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9354 = _T_4591 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9578 = _T_9577 | _T_9354; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9356 = _T_4595 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9579 = _T_9578 | _T_9356; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9358 = _T_4599 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9580 = _T_9579 | _T_9358; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9360 = _T_4603 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9581 = _T_9580 | _T_9360; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9362 = _T_4607 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9582 = _T_9581 | _T_9362; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9364 = _T_4611 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9583 = _T_9582 | _T_9364; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9366 = _T_4615 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9584 = _T_9583 | _T_9366; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9368 = _T_4619 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9585 = _T_9584 | _T_9368; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9370 = _T_4623 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9586 = _T_9585 | _T_9370; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9372 = _T_4627 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9587 = _T_9586 | _T_9372; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9374 = _T_4631 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9588 = _T_9587 | _T_9374; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9376 = _T_4635 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9589 = _T_9588 | _T_9376; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9378 = _T_4639 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9590 = _T_9589 | _T_9378; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9380 = _T_4643 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9591 = _T_9590 | _T_9380; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9382 = _T_4647 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9592 = _T_9591 | _T_9382; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9384 = _T_4651 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9593 = _T_9592 | _T_9384; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9386 = _T_4655 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9594 = _T_9593 | _T_9386; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9388 = _T_4659 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9595 = _T_9594 | _T_9388; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9390 = _T_4663 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9596 = _T_9595 | _T_9390; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9392 = _T_4667 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9597 = _T_9596 | _T_9392; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9394 = _T_4671 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9598 = _T_9597 | _T_9394; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9396 = _T_4675 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9599 = _T_9598 | _T_9396; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9398 = _T_4679 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9600 = _T_9599 | _T_9398; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9400 = _T_4683 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9601 = _T_9600 | _T_9400; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9402 = _T_4687 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9602 = _T_9601 | _T_9402; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9404 = _T_4691 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9603 = _T_9602 | _T_9404; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9406 = _T_4695 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9604 = _T_9603 | _T_9406; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9408 = _T_4699 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9605 = _T_9604 | _T_9408; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9410 = _T_4703 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9606 = _T_9605 | _T_9410; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9412 = _T_4707 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9607 = _T_9606 | _T_9412; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9414 = _T_4711 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9608 = _T_9607 | _T_9414; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9416 = _T_4715 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9609 = _T_9608 | _T_9416; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9418 = _T_4719 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9610 = _T_9609 | _T_9418; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9420 = _T_4723 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9611 = _T_9610 | _T_9420; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9422 = _T_4727 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9612 = _T_9611 | _T_9422; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9424 = _T_4731 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9613 = _T_9612 | _T_9424; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9426 = _T_4735 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9614 = _T_9613 | _T_9426; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9428 = _T_4739 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9615 = _T_9614 | _T_9428; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9430 = _T_4743 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9616 = _T_9615 | _T_9430; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9432 = _T_4747 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9617 = _T_9616 | _T_9432; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9434 = _T_4751 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9618 = _T_9617 | _T_9434; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9436 = _T_4755 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9619 = _T_9618 | _T_9436; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9438 = _T_4759 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9620 = _T_9619 | _T_9438; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9440 = _T_4763 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9621 = _T_9620 | _T_9440; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9442 = _T_4767 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9622 = _T_9621 | _T_9442; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9444 = _T_4771 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9623 = _T_9622 | _T_9444; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9446 = _T_4775 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9624 = _T_9623 | _T_9446; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9448 = _T_4779 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9625 = _T_9624 | _T_9448; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9450 = _T_4783 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9626 = _T_9625 | _T_9450; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9452 = _T_4787 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9627 = _T_9626 | _T_9452; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9454 = _T_4791 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9628 = _T_9627 | _T_9454; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9456 = _T_4795 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9629 = _T_9628 | _T_9456; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9458 = _T_4799 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9630 = _T_9629 | _T_9458; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9460 = _T_4803 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9631 = _T_9630 | _T_9460; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9462 = _T_4807 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9632 = _T_9631 | _T_9462; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9464 = _T_4811 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9633 = _T_9632 | _T_9464; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9466 = _T_4815 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9634 = _T_9633 | _T_9466; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9468 = _T_4819 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9635 = _T_9634 | _T_9468; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9470 = _T_4823 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9636 = _T_9635 | _T_9470; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9472 = _T_4827 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9637 = _T_9636 | _T_9472; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9474 = _T_4831 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9638 = _T_9637 | _T_9474; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9476 = _T_4835 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9639 = _T_9638 | _T_9476; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9478 = _T_4839 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9640 = _T_9639 | _T_9478; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9480 = _T_4843 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9641 = _T_9640 | _T_9480; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9482 = _T_4847 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9642 = _T_9641 | _T_9482; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9484 = _T_4851 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9643 = _T_9642 | _T_9484; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9486 = _T_4855 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9644 = _T_9643 | _T_9486; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9488 = _T_4859 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9645 = _T_9644 | _T_9488; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9490 = _T_4863 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9646 = _T_9645 | _T_9490; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9492 = _T_4867 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9647 = _T_9646 | _T_9492; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9494 = _T_4871 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9648 = _T_9647 | _T_9494; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9496 = _T_4875 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9649 = _T_9648 | _T_9496; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9498 = _T_4879 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9650 = _T_9649 | _T_9498; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9500 = _T_4883 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9651 = _T_9650 | _T_9500; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9502 = _T_4887 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9652 = _T_9651 | _T_9502; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9504 = _T_4891 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9653 = _T_9652 | _T_9504; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9506 = _T_4895 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9654 = _T_9653 | _T_9506; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9508 = _T_4899 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9655 = _T_9654 | _T_9508; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9510 = _T_4903 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9656 = _T_9655 | _T_9510; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9512 = _T_4907 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9657 = _T_9656 | _T_9512; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9514 = _T_4911 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9658 = _T_9657 | _T_9514; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9516 = _T_4915 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9659 = _T_9658 | _T_9516; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9518 = _T_4919 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9660 = _T_9659 | _T_9518; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9520 = _T_4923 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9661 = _T_9660 | _T_9520; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9522 = _T_4927 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9662 = _T_9661 | _T_9522; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9524 = _T_4931 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9663 = _T_9662 | _T_9524; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9526 = _T_4935 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9664 = _T_9663 | _T_9526; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9528 = _T_4939 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9665 = _T_9664 | _T_9528; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9530 = _T_4943 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9666 = _T_9665 | _T_9530; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9532 = _T_4947 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9667 = _T_9666 | _T_9532; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9534 = _T_4951 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9668 = _T_9667 | _T_9534; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9536 = _T_4955 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9669 = _T_9668 | _T_9536; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9538 = _T_4959 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9670 = _T_9669 | _T_9538; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9540 = _T_4963 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9671 = _T_9670 | _T_9540; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9542 = _T_4967 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9672 = _T_9671 | _T_9542; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9544 = _T_4971 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9673 = _T_9672 | _T_9544; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9546 = _T_4975 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9674 = _T_9673 | _T_9546; // @[el2_ifu_mem_ctl.scala 745:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9548 = _T_4979 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 745:10]
  wire  _T_9675 = _T_9674 | _T_9548; // @[el2_ifu_mem_ctl.scala 745:91]
  wire [1:0] ic_tag_valid_unq = {_T_10058,_T_9675}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 818:54]
  wire [1:0] _T_10097 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10098 = ic_debug_way_ff & _T_10097; // @[el2_ifu_mem_ctl.scala 799:67]
  wire [1:0] _T_10099 = ic_tag_valid_unq & _T_10098; // @[el2_ifu_mem_ctl.scala 799:48]
  wire  ic_debug_tag_val_rd_out = |_T_10099; // @[el2_ifu_mem_ctl.scala 799:115]
  wire [65:0] _T_1210 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1211; // @[el2_ifu_mem_ctl.scala 349:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2539; // @[el2_ifu_mem_ctl.scala 359:80]
  wire  _T_1251 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 364:98]
  wire  sel_byp_data = _T_1255 & _T_1251; // @[el2_ifu_mem_ctl.scala 364:96]
  wire [63:0] _T_1262 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1263 = _T_1262 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 371:64]
  wire [63:0] _T_1265 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2101 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 440:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1615 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1663 = _T_1615 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1618 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1664 = _T_1618 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1679 = _T_1663 | _T_1664; // @[Mux.scala 27:72]
  wire  _T_1621 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1665 = _T_1621 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1680 = _T_1679 | _T_1665; // @[Mux.scala 27:72]
  wire  _T_1624 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1666 = _T_1624 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1681 = _T_1680 | _T_1666; // @[Mux.scala 27:72]
  wire  _T_1627 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1667 = _T_1627 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1682 = _T_1681 | _T_1667; // @[Mux.scala 27:72]
  wire  _T_1630 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1668 = _T_1630 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1683 = _T_1682 | _T_1668; // @[Mux.scala 27:72]
  wire  _T_1633 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1669 = _T_1633 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1684 = _T_1683 | _T_1669; // @[Mux.scala 27:72]
  wire  _T_1636 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1670 = _T_1636 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1685 = _T_1684 | _T_1670; // @[Mux.scala 27:72]
  wire  _T_1639 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1671 = _T_1639 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1686 = _T_1685 | _T_1671; // @[Mux.scala 27:72]
  wire  _T_1642 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1672 = _T_1642 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1687 = _T_1686 | _T_1672; // @[Mux.scala 27:72]
  wire  _T_1645 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1673 = _T_1645 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1688 = _T_1687 | _T_1673; // @[Mux.scala 27:72]
  wire  _T_1648 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1674 = _T_1648 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1689 = _T_1688 | _T_1674; // @[Mux.scala 27:72]
  wire  _T_1651 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1675 = _T_1651 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1690 = _T_1689 | _T_1675; // @[Mux.scala 27:72]
  wire  _T_1654 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1676 = _T_1654 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1690 | _T_1676; // @[Mux.scala 27:72]
  wire  _T_1657 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1677 = _T_1657 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1692 = _T_1691 | _T_1677; // @[Mux.scala 27:72]
  wire  _T_1660 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 437:73]
  wire [15:0] _T_1678 = _T_1660 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1692 | _T_1678; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1695 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1743 = _T_1695 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1698 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1744 = _T_1698 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1759 = _T_1743 | _T_1744; // @[Mux.scala 27:72]
  wire  _T_1701 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1745 = _T_1701 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1760 = _T_1759 | _T_1745; // @[Mux.scala 27:72]
  wire  _T_1704 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1746 = _T_1704 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1761 = _T_1760 | _T_1746; // @[Mux.scala 27:72]
  wire  _T_1707 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1747 = _T_1707 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1762 = _T_1761 | _T_1747; // @[Mux.scala 27:72]
  wire  _T_1710 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1748 = _T_1710 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1763 = _T_1762 | _T_1748; // @[Mux.scala 27:72]
  wire  _T_1713 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1749 = _T_1713 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1764 = _T_1763 | _T_1749; // @[Mux.scala 27:72]
  wire  _T_1716 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1750 = _T_1716 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1765 = _T_1764 | _T_1750; // @[Mux.scala 27:72]
  wire  _T_1719 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1751 = _T_1719 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1766 = _T_1765 | _T_1751; // @[Mux.scala 27:72]
  wire  _T_1722 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1752 = _T_1722 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1767 = _T_1766 | _T_1752; // @[Mux.scala 27:72]
  wire  _T_1725 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1753 = _T_1725 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1768 = _T_1767 | _T_1753; // @[Mux.scala 27:72]
  wire  _T_1728 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1754 = _T_1728 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1769 = _T_1768 | _T_1754; // @[Mux.scala 27:72]
  wire  _T_1731 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1755 = _T_1731 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1770 = _T_1769 | _T_1755; // @[Mux.scala 27:72]
  wire  _T_1734 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1756 = _T_1734 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1770 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1737 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1757 = _T_1737 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1772 = _T_1771 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1740 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 437:179]
  wire [31:0] _T_1758 = _T_1740 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1772 | _T_1758; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1775 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1823 = _T_1775 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1778 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1824 = _T_1778 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1839 = _T_1823 | _T_1824; // @[Mux.scala 27:72]
  wire  _T_1781 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1825 = _T_1781 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1840 = _T_1839 | _T_1825; // @[Mux.scala 27:72]
  wire  _T_1784 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1826 = _T_1784 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1841 = _T_1840 | _T_1826; // @[Mux.scala 27:72]
  wire  _T_1787 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1827 = _T_1787 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1842 = _T_1841 | _T_1827; // @[Mux.scala 27:72]
  wire  _T_1790 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1828 = _T_1790 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1843 = _T_1842 | _T_1828; // @[Mux.scala 27:72]
  wire  _T_1793 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1829 = _T_1793 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1844 = _T_1843 | _T_1829; // @[Mux.scala 27:72]
  wire  _T_1796 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1830 = _T_1796 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1845 = _T_1844 | _T_1830; // @[Mux.scala 27:72]
  wire  _T_1799 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1831 = _T_1799 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1846 = _T_1845 | _T_1831; // @[Mux.scala 27:72]
  wire  _T_1802 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1832 = _T_1802 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1847 = _T_1846 | _T_1832; // @[Mux.scala 27:72]
  wire  _T_1805 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1833 = _T_1805 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1848 = _T_1847 | _T_1833; // @[Mux.scala 27:72]
  wire  _T_1808 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1834 = _T_1808 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1849 = _T_1848 | _T_1834; // @[Mux.scala 27:72]
  wire  _T_1811 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1835 = _T_1811 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1850 = _T_1849 | _T_1835; // @[Mux.scala 27:72]
  wire  _T_1814 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1836 = _T_1814 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1850 | _T_1836; // @[Mux.scala 27:72]
  wire  _T_1817 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1837 = _T_1817 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1852 = _T_1851 | _T_1837; // @[Mux.scala 27:72]
  wire  _T_1820 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 437:285]
  wire [31:0] _T_1838 = _T_1820 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1852 | _T_1838; // @[Mux.scala 27:72]
  wire [79:0] _T_1856 = {_T_1693,_T_1773,_T_1853}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1857 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1905 = _T_1857 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1860 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1906 = _T_1860 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1921 = _T_1905 | _T_1906; // @[Mux.scala 27:72]
  wire  _T_1863 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1907 = _T_1863 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1922 = _T_1921 | _T_1907; // @[Mux.scala 27:72]
  wire  _T_1866 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1908 = _T_1866 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1923 = _T_1922 | _T_1908; // @[Mux.scala 27:72]
  wire  _T_1869 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1909 = _T_1869 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1924 = _T_1923 | _T_1909; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1910 = _T_1872 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1925 = _T_1924 | _T_1910; // @[Mux.scala 27:72]
  wire  _T_1875 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1911 = _T_1875 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1926 = _T_1925 | _T_1911; // @[Mux.scala 27:72]
  wire  _T_1878 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1912 = _T_1878 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1927 = _T_1926 | _T_1912; // @[Mux.scala 27:72]
  wire  _T_1881 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1913 = _T_1881 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1928 = _T_1927 | _T_1913; // @[Mux.scala 27:72]
  wire  _T_1884 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1914 = _T_1884 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1929 = _T_1928 | _T_1914; // @[Mux.scala 27:72]
  wire  _T_1887 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1915 = _T_1887 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1930 = _T_1929 | _T_1915; // @[Mux.scala 27:72]
  wire  _T_1890 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1916 = _T_1890 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1931 = _T_1930 | _T_1916; // @[Mux.scala 27:72]
  wire  _T_1893 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1917 = _T_1893 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1932 = _T_1931 | _T_1917; // @[Mux.scala 27:72]
  wire  _T_1896 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1918 = _T_1896 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1932 | _T_1918; // @[Mux.scala 27:72]
  wire  _T_1899 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1919 = _T_1899 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1934 = _T_1933 | _T_1919; // @[Mux.scala 27:72]
  wire  _T_1902 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 438:73]
  wire [15:0] _T_1920 = _T_1902 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1934 | _T_1920; // @[Mux.scala 27:72]
  wire [31:0] _T_1985 = _T_1615 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1986 = _T_1618 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1985 | _T_1986; // @[Mux.scala 27:72]
  wire [31:0] _T_1987 = _T_1621 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_2001 | _T_1987; // @[Mux.scala 27:72]
  wire [31:0] _T_1988 = _T_1624 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_2002 | _T_1988; // @[Mux.scala 27:72]
  wire [31:0] _T_1989 = _T_1627 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_2003 | _T_1989; // @[Mux.scala 27:72]
  wire [31:0] _T_1990 = _T_1630 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_2004 | _T_1990; // @[Mux.scala 27:72]
  wire [31:0] _T_1991 = _T_1633 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_2005 | _T_1991; // @[Mux.scala 27:72]
  wire [31:0] _T_1992 = _T_1636 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_2006 | _T_1992; // @[Mux.scala 27:72]
  wire [31:0] _T_1993 = _T_1639 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_2007 | _T_1993; // @[Mux.scala 27:72]
  wire [31:0] _T_1994 = _T_1642 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_2008 | _T_1994; // @[Mux.scala 27:72]
  wire [31:0] _T_1995 = _T_1645 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_2009 | _T_1995; // @[Mux.scala 27:72]
  wire [31:0] _T_1996 = _T_1648 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_2010 | _T_1996; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1651 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_2011 | _T_1997; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1654 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_2012 | _T_1998; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1657 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_2013 | _T_1999; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1660 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_2014 | _T_2000; // @[Mux.scala 27:72]
  wire [79:0] _T_2098 = {_T_1935,_T_2015,_T_1773}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_2101 ? _T_1856 : _T_2098; // @[el2_ifu_mem_ctl.scala 436:37]
  wire [79:0] _T_2103 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2101 ? ic_byp_data_only_pre_new : _T_2103; // @[el2_ifu_mem_ctl.scala 440:30]
  wire [79:0] _GEN_793 = {{16'd0}, _T_1265}; // @[el2_ifu_mem_ctl.scala 371:109]
  wire [79:0] _T_1266 = _GEN_793 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 371:109]
  wire [79:0] _GEN_794 = {{16'd0}, _T_1263}; // @[el2_ifu_mem_ctl.scala 371:83]
  wire [79:0] ic_premux_data = _GEN_794 | _T_1266; // @[el2_ifu_mem_ctl.scala 371:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 378:38]
  wire [1:0] _T_1275 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 382:8]
  wire [7:0] _T_1356 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1361 = ic_miss_buff_data_error[0] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  _T_2607 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 614:47]
  wire  _T_2608 = _T_2607 & _T_13; // @[el2_ifu_mem_ctl.scala 614:50]
  wire  bus_ifu_wr_data_error = _T_2608 & miss_pending; // @[el2_ifu_mem_ctl.scala 614:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1361; // @[el2_ifu_mem_ctl.scala 402:72]
  wire  _T_1365 = ic_miss_buff_data_error[1] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1365; // @[el2_ifu_mem_ctl.scala 402:72]
  wire  _T_1369 = ic_miss_buff_data_error[2] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1369; // @[el2_ifu_mem_ctl.scala 402:72]
  wire  _T_1373 = ic_miss_buff_data_error[3] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1373; // @[el2_ifu_mem_ctl.scala 402:72]
  wire  _T_1377 = ic_miss_buff_data_error[4] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1377; // @[el2_ifu_mem_ctl.scala 402:72]
  wire  _T_1381 = ic_miss_buff_data_error[5] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1381; // @[el2_ifu_mem_ctl.scala 402:72]
  wire  _T_1385 = ic_miss_buff_data_error[6] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1385; // @[el2_ifu_mem_ctl.scala 402:72]
  wire  _T_1389 = ic_miss_buff_data_error[7] & _T_1327; // @[el2_ifu_mem_ctl.scala 403:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1389; // @[el2_ifu_mem_ctl.scala 402:72]
  wire [7:0] _T_1396 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2413 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2421 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 483:65]
  wire  _T_2422 = _T_2421 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 483:88]
  wire  _T_2424 = _T_2422 & _T_2535; // @[el2_ifu_mem_ctl.scala 483:112]
  wire  _T_2425 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2426 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 488:50]
  wire  _T_2428 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2434 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2436 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2434 | _T_2436; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2428 ? _T_2426 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2425 ? _T_2426 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2413 ? _T_2424 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2413 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2427 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 489:56]
  wire  _GEN_43 = _T_2425 & _T_2427; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2413 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 474:58]
  wire  _T_2410 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 473:49]
  wire  _T_2415 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 482:87]
  wire  _T_2429 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 492:54]
  wire  _T_2430 = _T_2429 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 492:84]
  wire  _T_2439 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 513:66]
  wire  _T_2440 = io_dec_tlu_flush_err_wb & _T_2439; // @[el2_ifu_mem_ctl.scala 513:52]
  wire  _T_2442 = _T_2440 & _T_2535; // @[el2_ifu_mem_ctl.scala 513:81]
  wire  _T_2444 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 516:59]
  wire  _T_2445 = _T_2444 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 516:86]
  wire  _T_2459 = _T_2444 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 519:81]
  wire  _T_2460 = _T_2459 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 519:103]
  wire  _T_2461 = _T_2460 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 519:126]
  wire  _T_2481 = _T_2459 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 526:103]
  wire  _T_2488 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 531:62]
  wire  _T_2489 = io_dec_tlu_flush_lower_wb & _T_2488; // @[el2_ifu_mem_ctl.scala 531:60]
  wire  _T_2490 = _T_2489 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 531:88]
  wire  _T_2491 = _T_2490 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 531:115]
  wire  _GEN_50 = _T_2487 & _T_2445; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_2470 ? _T_2481 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_2470 | _T_2487; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_2443 ? _T_2461 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2443 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2438 ? _T_2442 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2503 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 548:64]
  wire  _T_2505 = _T_2503 & _T_2535; // @[el2_ifu_mem_ctl.scala 548:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2507 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 548:133]
  wire  _T_2508 = _T_2507 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 548:164]
  wire  _T_2509 = _T_2508 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 548:184]
  wire  _T_2510 = _T_2509 & miss_pending; // @[el2_ifu_mem_ctl.scala 548:204]
  wire  _T_2511 = ~_T_2510; // @[el2_ifu_mem_ctl.scala 548:112]
  wire  ifc_bus_ic_req_ff_in = _T_2505 & _T_2511; // @[el2_ifu_mem_ctl.scala 548:110]
  wire  _T_2512 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 549:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 580:45]
  wire  _T_2529 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 583:35]
  wire  _T_2530 = _T_2529 & miss_pending; // @[el2_ifu_mem_ctl.scala 583:53]
  wire  bus_cmd_sent = _T_2530 & _T_2535; // @[el2_ifu_mem_ctl.scala 583:68]
  wire [2:0] _T_2520 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2522 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2524 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 581:51]
  wire  _T_2550 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 591:73]
  wire  _T_2551 = _T_2536 & _T_2550; // @[el2_ifu_mem_ctl.scala 591:71]
  wire  _T_2553 = last_data_recieved_ff & _T_1327; // @[el2_ifu_mem_ctl.scala 591:114]
  wire  last_data_recieved_in = _T_2551 | _T_2553; // @[el2_ifu_mem_ctl.scala 591:89]
  wire [2:0] _T_2559 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 596:45]
  wire  _T_2562 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 597:81]
  wire  _T_2563 = _T_2562 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 597:97]
  wire  _T_2565 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 599:48]
  wire  _T_2566 = _T_2565 & miss_pending; // @[el2_ifu_mem_ctl.scala 599:68]
  wire  bus_inc_cmd_beat_cnt = _T_2566 & _T_2535; // @[el2_ifu_mem_ctl.scala 599:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 601:57]
  wire  _T_2570 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 602:31]
  wire  _T_2571 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 602:71]
  wire  _T_2572 = _T_2571 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 602:87]
  wire  _T_2573 = ~_T_2572; // @[el2_ifu_mem_ctl.scala 602:55]
  wire  bus_hold_cmd_beat_cnt = _T_2570 & _T_2573; // @[el2_ifu_mem_ctl.scala 602:53]
  wire  _T_2574 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 603:46]
  wire  bus_cmd_beat_en = _T_2574 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 603:62]
  wire [2:0] _T_2577 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 605:46]
  wire [2:0] _T_2579 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2580 = bus_inc_cmd_beat_cnt ? _T_2577 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2581 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2583 = _T_2579 | _T_2580; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2583 | _T_2581; // @[Mux.scala 27:72]
  wire  _T_2587 = _T_2563 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 606:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 617:62]
  wire  _T_2615 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 622:50]
  wire  _T_2616 = io_ifc_dma_access_ok & _T_2615; // @[el2_ifu_mem_ctl.scala 622:47]
  wire  _T_2617 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 622:70]
  wire  ifc_dma_access_ok_d = _T_2616 & _T_2617; // @[el2_ifu_mem_ctl.scala 622:68]
  wire  _T_2621 = _T_2616 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 623:72]
  wire  _T_2622 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 623:111]
  wire  _T_2623 = _T_2621 & _T_2622; // @[el2_ifu_mem_ctl.scala 623:97]
  wire  ifc_dma_access_q_ok = _T_2623 & _T_2617; // @[el2_ifu_mem_ctl.scala 623:127]
  wire  _T_2626 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 626:40]
  wire  _T_2627 = _T_2626 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 626:58]
  wire  _T_2630 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 627:60]
  wire  _T_2631 = _T_2626 & _T_2630; // @[el2_ifu_mem_ctl.scala 627:58]
  wire  _T_2632 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 627:104]
  wire [2:0] _T_2637 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2743 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2752 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2743}; // @[el2_lib.scala 268:22]
  wire  _T_2753 = ^_T_2752; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2761 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2770 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2761}; // @[el2_lib.scala 268:39]
  wire  _T_2771 = ^_T_2770; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2779 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2788 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2779}; // @[el2_lib.scala 268:56]
  wire  _T_2789 = ^_T_2788; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2795 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2803 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2795}; // @[el2_lib.scala 268:73]
  wire  _T_2804 = ^_T_2803; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2818 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2795}; // @[el2_lib.scala 268:90]
  wire  _T_2819 = ^_T_2818; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2824 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2825 = ^_T_2824; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2830 = {_T_2753,_T_2771,_T_2789,_T_2804,_T_2819,_T_2825}; // @[Cat.scala 29:58]
  wire  _T_2831 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2832 = ^_T_2830; // @[el2_lib.scala 269:23]
  wire  _T_2833 = _T_2831 ^ _T_2832; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2939 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2948 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2939}; // @[el2_lib.scala 268:22]
  wire  _T_2949 = ^_T_2948; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2957 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2966 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2957}; // @[el2_lib.scala 268:39]
  wire  _T_2967 = ^_T_2966; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2975 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2984 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2975}; // @[el2_lib.scala 268:56]
  wire  _T_2985 = ^_T_2984; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2991 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2999 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2991}; // @[el2_lib.scala 268:73]
  wire  _T_3000 = ^_T_2999; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3014 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2991}; // @[el2_lib.scala 268:90]
  wire  _T_3015 = ^_T_3014; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3020 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3021 = ^_T_3020; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3026 = {_T_2949,_T_2967,_T_2985,_T_3000,_T_3015,_T_3021}; // @[Cat.scala 29:58]
  wire  _T_3027 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3028 = ^_T_3026; // @[el2_lib.scala 269:23]
  wire  _T_3029 = _T_3027 ^ _T_3028; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3030 = {_T_3029,_T_2949,_T_2967,_T_2985,_T_3000,_T_3015,_T_3021}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2833,_T_2753,_T_2771,_T_2789,_T_2804,_T_2819,_T_2825,_T_3030}; // @[Cat.scala 29:58]
  wire  _T_3032 = ~_T_2626; // @[el2_ifu_mem_ctl.scala 632:45]
  wire  _T_3033 = iccm_correct_ecc & _T_3032; // @[el2_ifu_mem_ctl.scala 632:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3034 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3041 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 646:53]
  wire  _T_3373 = _T_3285[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3371 = _T_3285[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3369 = _T_3285[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3367 = _T_3285[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3365 = _T_3285[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3363 = _T_3285[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3361 = _T_3285[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3359 = _T_3285[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3357 = _T_3285[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3355 = _T_3285[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3431 = {_T_3373,_T_3371,_T_3369,_T_3367,_T_3365,_T_3363,_T_3361,_T_3359,_T_3357,_T_3355}; // @[el2_lib.scala 310:69]
  wire  _T_3353 = _T_3285[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3351 = _T_3285[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3349 = _T_3285[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3347 = _T_3285[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3345 = _T_3285[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3343 = _T_3285[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3341 = _T_3285[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3339 = _T_3285[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3337 = _T_3285[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3335 = _T_3285[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3422 = {_T_3353,_T_3351,_T_3349,_T_3347,_T_3345,_T_3343,_T_3341,_T_3339,_T_3337,_T_3335}; // @[el2_lib.scala 310:69]
  wire  _T_3333 = _T_3285[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3331 = _T_3285[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3329 = _T_3285[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3327 = _T_3285[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3325 = _T_3285[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3323 = _T_3285[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3321 = _T_3285[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3319 = _T_3285[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3317 = _T_3285[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3315 = _T_3285[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3412 = {_T_3333,_T_3331,_T_3329,_T_3327,_T_3325,_T_3323,_T_3321,_T_3319,_T_3317,_T_3315}; // @[el2_lib.scala 310:69]
  wire  _T_3313 = _T_3285[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3311 = _T_3285[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3309 = _T_3285[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3307 = _T_3285[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3305 = _T_3285[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3303 = _T_3285[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3301 = _T_3285[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3299 = _T_3285[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3297 = _T_3285[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3413 = {_T_3412,_T_3313,_T_3311,_T_3309,_T_3307,_T_3305,_T_3303,_T_3301,_T_3299,_T_3297}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3433 = {_T_3431,_T_3422,_T_3413}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3388 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3394 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3388}; // @[Cat.scala 29:58]
  wire [38:0] _T_3434 = _T_3433 ^ _T_3394; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3435 = _T_3289 ? _T_3434 : _T_3394; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3435[37:32],_T_3435[30:16],_T_3435[14:8],_T_3435[6:4],_T_3435[2]}; // @[Cat.scala 29:58]
  wire  _T_3758 = _T_3670[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3756 = _T_3670[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3754 = _T_3670[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3752 = _T_3670[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3750 = _T_3670[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3748 = _T_3670[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3746 = _T_3670[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3744 = _T_3670[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3742 = _T_3670[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3740 = _T_3670[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3816 = {_T_3758,_T_3756,_T_3754,_T_3752,_T_3750,_T_3748,_T_3746,_T_3744,_T_3742,_T_3740}; // @[el2_lib.scala 310:69]
  wire  _T_3738 = _T_3670[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3736 = _T_3670[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3734 = _T_3670[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3732 = _T_3670[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3730 = _T_3670[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3728 = _T_3670[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3726 = _T_3670[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3724 = _T_3670[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3722 = _T_3670[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3720 = _T_3670[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3807 = {_T_3738,_T_3736,_T_3734,_T_3732,_T_3730,_T_3728,_T_3726,_T_3724,_T_3722,_T_3720}; // @[el2_lib.scala 310:69]
  wire  _T_3718 = _T_3670[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3716 = _T_3670[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3714 = _T_3670[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3712 = _T_3670[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3710 = _T_3670[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3708 = _T_3670[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3706 = _T_3670[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3704 = _T_3670[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3702 = _T_3670[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3700 = _T_3670[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3797 = {_T_3718,_T_3716,_T_3714,_T_3712,_T_3710,_T_3708,_T_3706,_T_3704,_T_3702,_T_3700}; // @[el2_lib.scala 310:69]
  wire  _T_3698 = _T_3670[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3696 = _T_3670[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3694 = _T_3670[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3692 = _T_3670[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3690 = _T_3670[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3688 = _T_3670[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3686 = _T_3670[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3684 = _T_3670[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3682 = _T_3670[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3798 = {_T_3797,_T_3698,_T_3696,_T_3694,_T_3692,_T_3690,_T_3688,_T_3686,_T_3684,_T_3682}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3818 = {_T_3816,_T_3807,_T_3798}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3773 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3779 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3773}; // @[Cat.scala 29:58]
  wire [38:0] _T_3819 = _T_3818 ^ _T_3779; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3820 = _T_3674 ? _T_3819 : _T_3779; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3820[37:32],_T_3820[30:16],_T_3820[14:8],_T_3820[6:4],_T_3820[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 638:35]
  wire  _T_3293 = ~_T_3285[6]; // @[el2_lib.scala 303:55]
  wire  _T_3294 = _T_3287 & _T_3293; // @[el2_lib.scala 303:53]
  wire  _T_3678 = ~_T_3670[6]; // @[el2_lib.scala 303:55]
  wire  _T_3679 = _T_3672 & _T_3678; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3294,_T_3679}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 640:53]
  wire [63:0] _T_3045 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3046 = {iccm_dma_rdata_1_muxed,_T_3435[37:32],_T_3435[30:16],_T_3435[14:8],_T_3435[6:4],_T_3435[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 642:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 643:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 648:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 652:70]
  wire  _T_3051 = _T_2626 & _T_2615; // @[el2_ifu_mem_ctl.scala 655:65]
  wire  _T_3054 = _T_3032 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 656:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3055 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3057 = _T_3054 ? {{1'd0}, _T_3055} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 656:8]
  wire [31:0] _T_3058 = _T_3051 ? io_dma_mem_addr : {{16'd0}, _T_3057}; // @[el2_ifu_mem_ctl.scala 655:25]
  wire  _T_3447 = _T_3285 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3448 = _T_3435[38] ^ _T_3447; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3448,_T_3435[31],_T_3435[15],_T_3435[7],_T_3435[3],_T_3435[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3832 = _T_3670 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3833 = _T_3820[38] ^ _T_3832; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3833,_T_3820[31],_T_3820[15],_T_3820[7],_T_3820[3],_T_3820[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3849 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 668:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 670:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 671:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 679:62]
  wire  _T_3857 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 673:76]
  wire  _T_3858 = io_iccm_rd_ecc_single_err & _T_3857; // @[el2_ifu_mem_ctl.scala 673:74]
  wire  _T_3860 = _T_3858 & _T_317; // @[el2_ifu_mem_ctl.scala 673:104]
  wire  iccm_ecc_write_status = _T_3860 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 673:127]
  wire  _T_3861 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 674:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3861 & _T_317; // @[el2_ifu_mem_ctl.scala 674:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 678:51]
  wire [13:0] _T_3866 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 677:102]
  wire [38:0] _T_3870 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3875 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 682:41]
  wire  _T_3876 = io_ifc_fetch_req_bf & _T_3875; // @[el2_ifu_mem_ctl.scala 682:39]
  wire  _T_3877 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 682:72]
  wire  _T_3878 = _T_3876 & _T_3877; // @[el2_ifu_mem_ctl.scala 682:70]
  wire  _T_3880 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 683:34]
  wire  _T_3881 = _T_2221 & _T_3880; // @[el2_ifu_mem_ctl.scala 683:32]
  wire  _T_3884 = _T_2237 & _T_3880; // @[el2_ifu_mem_ctl.scala 684:37]
  wire  _T_3885 = _T_3881 | _T_3884; // @[el2_ifu_mem_ctl.scala 683:88]
  wire  _T_3886 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 685:19]
  wire  _T_3888 = _T_3886 & _T_3880; // @[el2_ifu_mem_ctl.scala 685:41]
  wire  _T_3889 = _T_3885 | _T_3888; // @[el2_ifu_mem_ctl.scala 684:88]
  wire  _T_3890 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 686:19]
  wire  _T_3892 = _T_3890 & _T_3880; // @[el2_ifu_mem_ctl.scala 686:35]
  wire  _T_3893 = _T_3889 | _T_3892; // @[el2_ifu_mem_ctl.scala 685:88]
  wire  _T_3896 = _T_2236 & _T_3880; // @[el2_ifu_mem_ctl.scala 687:38]
  wire  _T_3897 = _T_3893 | _T_3896; // @[el2_ifu_mem_ctl.scala 686:88]
  wire  _T_3899 = _T_2237 & miss_state_en; // @[el2_ifu_mem_ctl.scala 688:37]
  wire  _T_3900 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 688:71]
  wire  _T_3901 = _T_3899 & _T_3900; // @[el2_ifu_mem_ctl.scala 688:54]
  wire  _T_3902 = _T_3897 | _T_3901; // @[el2_ifu_mem_ctl.scala 687:57]
  wire  _T_3903 = ~_T_3902; // @[el2_ifu_mem_ctl.scala 683:5]
  wire  _T_3904 = _T_3878 & _T_3903; // @[el2_ifu_mem_ctl.scala 682:96]
  wire  _T_3905 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 689:28]
  wire  _T_3907 = _T_3905 & _T_3875; // @[el2_ifu_mem_ctl.scala 689:50]
  wire  _T_3909 = _T_3907 & _T_3877; // @[el2_ifu_mem_ctl.scala 689:81]
  wire  _T_3918 = ~_T_108; // @[el2_ifu_mem_ctl.scala 692:106]
  wire  _T_3919 = _T_2221 & _T_3918; // @[el2_ifu_mem_ctl.scala 692:104]
  wire  _T_3920 = _T_2237 | _T_3919; // @[el2_ifu_mem_ctl.scala 692:77]
  wire  _T_3924 = ~_T_51; // @[el2_ifu_mem_ctl.scala 692:172]
  wire  _T_3925 = _T_3920 & _T_3924; // @[el2_ifu_mem_ctl.scala 692:170]
  wire  _T_3926 = ~_T_3925; // @[el2_ifu_mem_ctl.scala 692:44]
  wire  _T_3930 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 695:64]
  wire  _T_3931 = ~_T_3930; // @[el2_ifu_mem_ctl.scala 695:50]
  wire  _T_3932 = _T_276 & _T_3931; // @[el2_ifu_mem_ctl.scala 695:48]
  wire  _T_3933 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 695:81]
  wire  ic_valid = _T_3932 & _T_3933; // @[el2_ifu_mem_ctl.scala 695:79]
  wire  _T_3935 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 696:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 699:14]
  wire  _T_3938 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 702:74]
  wire  _T_10080 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 776:45]
  wire  way_status_wr_en = _T_10080 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 776:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3938; // @[el2_ifu_mem_ctl.scala 702:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 704:14]
  wire [2:0] _T_3942 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 708:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 772:41]
  wire  way_status_new = _T_10080 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 775:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 710:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 712:132]
  wire  _T_3959 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3960 = _T_3959 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3961 = _T_3960 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3963 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3964 = _T_3963 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3965 = _T_3964 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3967 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3968 = _T_3967 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3969 = _T_3968 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3971 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3972 = _T_3971 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3973 = _T_3972 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3975 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3976 = _T_3975 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3977 = _T_3976 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3979 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3980 = _T_3979 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3981 = _T_3980 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3983 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3984 = _T_3983 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3985 = _T_3984 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3987 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 716:93]
  wire  _T_3988 = _T_3987 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 716:102]
  wire  _T_3989 = _T_3988 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3993 = _T_3960 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_3997 = _T_3964 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4001 = _T_3968 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4005 = _T_3972 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4009 = _T_3976 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4013 = _T_3980 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4017 = _T_3984 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4021 = _T_3988 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4025 = _T_3960 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4029 = _T_3964 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4033 = _T_3968 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4037 = _T_3972 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4041 = _T_3976 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4045 = _T_3980 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4049 = _T_3984 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4053 = _T_3988 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4057 = _T_3960 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4061 = _T_3964 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4065 = _T_3968 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4069 = _T_3972 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4073 = _T_3976 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4077 = _T_3980 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4081 = _T_3984 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4085 = _T_3988 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4089 = _T_3960 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4093 = _T_3964 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4097 = _T_3968 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4101 = _T_3972 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4105 = _T_3976 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4109 = _T_3980 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4113 = _T_3984 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4117 = _T_3988 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4121 = _T_3960 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4125 = _T_3964 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4129 = _T_3968 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4133 = _T_3972 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4137 = _T_3976 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4141 = _T_3980 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4145 = _T_3984 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4149 = _T_3988 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4153 = _T_3960 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4157 = _T_3964 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4161 = _T_3968 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4165 = _T_3972 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4169 = _T_3976 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4173 = _T_3980 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4177 = _T_3984 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4181 = _T_3988 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4185 = _T_3960 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4189 = _T_3964 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4193 = _T_3968 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4197 = _T_3972 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4201 = _T_3976 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4205 = _T_3980 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4209 = _T_3984 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4213 = _T_3988 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4217 = _T_3960 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4221 = _T_3964 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4225 = _T_3968 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4229 = _T_3972 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4233 = _T_3976 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4237 = _T_3980 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4241 = _T_3984 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4245 = _T_3988 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4249 = _T_3960 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4253 = _T_3964 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4257 = _T_3968 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4261 = _T_3972 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4265 = _T_3976 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4269 = _T_3980 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4273 = _T_3984 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4277 = _T_3988 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4281 = _T_3960 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4285 = _T_3964 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4289 = _T_3968 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4293 = _T_3972 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4297 = _T_3976 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4301 = _T_3980 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4305 = _T_3984 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4309 = _T_3988 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4313 = _T_3960 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4317 = _T_3964 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4321 = _T_3968 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4325 = _T_3972 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4329 = _T_3976 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4333 = _T_3980 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4337 = _T_3984 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4341 = _T_3988 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4345 = _T_3960 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4349 = _T_3964 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4353 = _T_3968 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4357 = _T_3972 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4361 = _T_3976 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4365 = _T_3980 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4369 = _T_3984 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4373 = _T_3988 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4377 = _T_3960 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4381 = _T_3964 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4385 = _T_3968 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4389 = _T_3972 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4393 = _T_3976 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4397 = _T_3980 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4401 = _T_3984 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4405 = _T_3988 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4409 = _T_3960 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4413 = _T_3964 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4417 = _T_3968 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4421 = _T_3972 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4425 = _T_3976 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4429 = _T_3980 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4433 = _T_3984 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4437 = _T_3988 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4441 = _T_3960 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4445 = _T_3964 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4449 = _T_3968 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4453 = _T_3972 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4457 = _T_3976 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4461 = _T_3980 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4465 = _T_3984 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_4469 = _T_3988 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 716:124]
  wire  _T_10086 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 779:84]
  wire  _T_10087 = _T_10086 & miss_pending; // @[el2_ifu_mem_ctl.scala 779:108]
  wire  bus_wren_last_1 = _T_10087 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 779:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 780:84]
  wire  _T_10089 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 781:73]
  wire  _T_10084 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 779:84]
  wire  _T_10085 = _T_10084 & miss_pending; // @[el2_ifu_mem_ctl.scala 779:108]
  wire  bus_wren_last_0 = _T_10085 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 779:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 780:84]
  wire  _T_10088 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 781:73]
  wire [1:0] ifu_tag_wren = {_T_10089,_T_10088}; // @[Cat.scala 29:58]
  wire [1:0] _T_10123 = _T_3938 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10123 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 814:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 725:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 727:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 731:14]
  wire  _T_5118 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 735:82]
  wire  _T_5120 = _T_5118 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5122 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 736:74]
  wire  _T_5124 = _T_5122 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5125 = _T_5120 | _T_5124; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5126 = _T_5125 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire  _T_5130 = _T_5118 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5134 = _T_5122 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5135 = _T_5130 | _T_5134; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5136 = _T_5135 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire [1:0] tag_valid_clken_0 = {_T_5126,_T_5136}; // @[Cat.scala 29:58]
  wire  _T_5138 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 735:82]
  wire  _T_5140 = _T_5138 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5142 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 736:74]
  wire  _T_5144 = _T_5142 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5145 = _T_5140 | _T_5144; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5146 = _T_5145 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire  _T_5150 = _T_5138 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5154 = _T_5142 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5155 = _T_5150 | _T_5154; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5156 = _T_5155 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire [1:0] tag_valid_clken_1 = {_T_5146,_T_5156}; // @[Cat.scala 29:58]
  wire  _T_5158 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 735:82]
  wire  _T_5160 = _T_5158 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5162 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 736:74]
  wire  _T_5164 = _T_5162 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5165 = _T_5160 | _T_5164; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5166 = _T_5165 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire  _T_5170 = _T_5158 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5174 = _T_5162 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5175 = _T_5170 | _T_5174; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5176 = _T_5175 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire [1:0] tag_valid_clken_2 = {_T_5166,_T_5176}; // @[Cat.scala 29:58]
  wire  _T_5178 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 735:82]
  wire  _T_5180 = _T_5178 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5182 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 736:74]
  wire  _T_5184 = _T_5182 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5185 = _T_5180 | _T_5184; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5186 = _T_5185 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire  _T_5190 = _T_5178 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5194 = _T_5182 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 736:83]
  wire  _T_5195 = _T_5190 | _T_5194; // @[el2_ifu_mem_ctl.scala 735:113]
  wire  _T_5196 = _T_5195 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 736:106]
  wire [1:0] tag_valid_clken_3 = {_T_5186,_T_5196}; // @[Cat.scala 29:58]
  wire  _T_5199 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 741:64]
  wire  _T_5200 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 741:91]
  wire  _T_5201 = _T_5199 & _T_5200; // @[el2_ifu_mem_ctl.scala 741:89]
  wire  _T_5204 = _T_4471 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5205 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5207 = _T_5205 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5209 = _T_5207 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5210 = _T_5204 | _T_5209; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5220 = _T_4475 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5221 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5223 = _T_5221 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5225 = _T_5223 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5226 = _T_5220 | _T_5225; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5236 = _T_4479 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5237 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5239 = _T_5237 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5241 = _T_5239 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5242 = _T_5236 | _T_5241; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5252 = _T_4483 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5253 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5255 = _T_5253 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5257 = _T_5255 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5258 = _T_5252 | _T_5257; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5268 = _T_4487 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5269 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5271 = _T_5269 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5273 = _T_5271 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5274 = _T_5268 | _T_5273; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5284 = _T_4491 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5285 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5287 = _T_5285 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5289 = _T_5287 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5290 = _T_5284 | _T_5289; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5300 = _T_4495 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5301 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5303 = _T_5301 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5305 = _T_5303 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5306 = _T_5300 | _T_5305; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5316 = _T_4499 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5317 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5319 = _T_5317 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5321 = _T_5319 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5322 = _T_5316 | _T_5321; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5332 = _T_4503 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5333 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5335 = _T_5333 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5337 = _T_5335 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5338 = _T_5332 | _T_5337; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5348 = _T_4507 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5349 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5351 = _T_5349 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5353 = _T_5351 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5354 = _T_5348 | _T_5353; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5364 = _T_4511 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5365 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5367 = _T_5365 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5369 = _T_5367 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5370 = _T_5364 | _T_5369; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5380 = _T_4515 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5381 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5383 = _T_5381 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5385 = _T_5383 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5386 = _T_5380 | _T_5385; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5396 = _T_4519 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5397 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5399 = _T_5397 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5401 = _T_5399 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5402 = _T_5396 | _T_5401; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5412 = _T_4523 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5413 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5415 = _T_5413 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5417 = _T_5415 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5418 = _T_5412 | _T_5417; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5428 = _T_4527 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5429 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5431 = _T_5429 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5433 = _T_5431 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5434 = _T_5428 | _T_5433; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5444 = _T_4531 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5445 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5447 = _T_5445 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5449 = _T_5447 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5450 = _T_5444 | _T_5449; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5460 = _T_4535 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5461 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5463 = _T_5461 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5465 = _T_5463 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5466 = _T_5460 | _T_5465; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5476 = _T_4539 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5477 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5479 = _T_5477 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5481 = _T_5479 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5482 = _T_5476 | _T_5481; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5492 = _T_4543 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5493 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5495 = _T_5493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5497 = _T_5495 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5498 = _T_5492 | _T_5497; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5508 = _T_4547 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5509 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5511 = _T_5509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5513 = _T_5511 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5514 = _T_5508 | _T_5513; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5524 = _T_4551 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5525 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5527 = _T_5525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5529 = _T_5527 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5530 = _T_5524 | _T_5529; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5540 = _T_4555 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5541 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5543 = _T_5541 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5545 = _T_5543 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5546 = _T_5540 | _T_5545; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5556 = _T_4559 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5557 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5559 = _T_5557 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5561 = _T_5559 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5562 = _T_5556 | _T_5561; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5572 = _T_4563 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5573 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5575 = _T_5573 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5577 = _T_5575 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5578 = _T_5572 | _T_5577; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5588 = _T_4567 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5589 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5591 = _T_5589 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5593 = _T_5591 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5594 = _T_5588 | _T_5593; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5604 = _T_4571 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5605 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5607 = _T_5605 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5609 = _T_5607 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5610 = _T_5604 | _T_5609; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5620 = _T_4575 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5621 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5623 = _T_5621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5625 = _T_5623 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5626 = _T_5620 | _T_5625; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5636 = _T_4579 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5637 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5639 = _T_5637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5641 = _T_5639 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5642 = _T_5636 | _T_5641; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5652 = _T_4583 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5653 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5655 = _T_5653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5657 = _T_5655 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5658 = _T_5652 | _T_5657; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5668 = _T_4587 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5669 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5671 = _T_5669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5673 = _T_5671 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5674 = _T_5668 | _T_5673; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5684 = _T_4591 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5685 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5687 = _T_5685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5689 = _T_5687 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5690 = _T_5684 | _T_5689; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5700 = _T_4595 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5701 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_5703 = _T_5701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5705 = _T_5703 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5706 = _T_5700 | _T_5705; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5716 = _T_4471 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5719 = _T_5205 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5721 = _T_5719 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5722 = _T_5716 | _T_5721; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5732 = _T_4475 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5735 = _T_5221 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5737 = _T_5735 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5738 = _T_5732 | _T_5737; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5748 = _T_4479 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5751 = _T_5237 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5753 = _T_5751 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5754 = _T_5748 | _T_5753; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5764 = _T_4483 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5767 = _T_5253 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5769 = _T_5767 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5770 = _T_5764 | _T_5769; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5780 = _T_4487 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5783 = _T_5269 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5785 = _T_5783 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5786 = _T_5780 | _T_5785; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5796 = _T_4491 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5799 = _T_5285 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5801 = _T_5799 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5802 = _T_5796 | _T_5801; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5812 = _T_4495 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5815 = _T_5301 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5817 = _T_5815 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5818 = _T_5812 | _T_5817; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5828 = _T_4499 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5831 = _T_5317 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5833 = _T_5831 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5834 = _T_5828 | _T_5833; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5844 = _T_4503 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5847 = _T_5333 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5849 = _T_5847 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5850 = _T_5844 | _T_5849; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5860 = _T_4507 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5863 = _T_5349 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5865 = _T_5863 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5866 = _T_5860 | _T_5865; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5876 = _T_4511 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5879 = _T_5365 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5881 = _T_5879 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5882 = _T_5876 | _T_5881; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5892 = _T_4515 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5895 = _T_5381 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5897 = _T_5895 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5898 = _T_5892 | _T_5897; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5908 = _T_4519 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5911 = _T_5397 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5913 = _T_5911 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5914 = _T_5908 | _T_5913; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5924 = _T_4523 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5927 = _T_5413 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5929 = _T_5927 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5930 = _T_5924 | _T_5929; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5940 = _T_4527 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5943 = _T_5429 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5945 = _T_5943 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5946 = _T_5940 | _T_5945; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5956 = _T_4531 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5959 = _T_5445 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5961 = _T_5959 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5962 = _T_5956 | _T_5961; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5972 = _T_4535 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5975 = _T_5461 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5977 = _T_5975 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5978 = _T_5972 | _T_5977; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_5988 = _T_4539 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_5991 = _T_5477 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_5993 = _T_5991 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_5994 = _T_5988 | _T_5993; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6004 = _T_4543 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6007 = _T_5493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6009 = _T_6007 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6010 = _T_6004 | _T_6009; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6020 = _T_4547 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6023 = _T_5509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6025 = _T_6023 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6026 = _T_6020 | _T_6025; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6036 = _T_4551 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6039 = _T_5525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6041 = _T_6039 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6042 = _T_6036 | _T_6041; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6052 = _T_4555 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6055 = _T_5541 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6057 = _T_6055 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6058 = _T_6052 | _T_6057; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6068 = _T_4559 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6071 = _T_5557 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6073 = _T_6071 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6074 = _T_6068 | _T_6073; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6084 = _T_4563 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6087 = _T_5573 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6089 = _T_6087 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6090 = _T_6084 | _T_6089; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6100 = _T_4567 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6103 = _T_5589 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6105 = _T_6103 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6106 = _T_6100 | _T_6105; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6116 = _T_4571 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6119 = _T_5605 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6121 = _T_6119 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6122 = _T_6116 | _T_6121; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6132 = _T_4575 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6135 = _T_5621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6137 = _T_6135 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6138 = _T_6132 | _T_6137; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6148 = _T_4579 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6151 = _T_5637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6153 = _T_6151 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6154 = _T_6148 | _T_6153; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6164 = _T_4583 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6167 = _T_5653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6169 = _T_6167 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6170 = _T_6164 | _T_6169; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6180 = _T_4587 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6183 = _T_5669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6185 = _T_6183 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6186 = _T_6180 | _T_6185; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6196 = _T_4591 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6199 = _T_5685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6201 = _T_6199 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6202 = _T_6196 | _T_6201; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6212 = _T_4595 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6215 = _T_5701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6217 = _T_6215 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6218 = _T_6212 | _T_6217; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6228 = _T_4599 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6229 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6231 = _T_6229 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6233 = _T_6231 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6234 = _T_6228 | _T_6233; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6244 = _T_4603 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6245 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6247 = _T_6245 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6249 = _T_6247 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6250 = _T_6244 | _T_6249; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6260 = _T_4607 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6261 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6263 = _T_6261 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6265 = _T_6263 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6266 = _T_6260 | _T_6265; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6276 = _T_4611 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6277 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6279 = _T_6277 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6281 = _T_6279 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6282 = _T_6276 | _T_6281; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6292 = _T_4615 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6293 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6295 = _T_6293 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6297 = _T_6295 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6298 = _T_6292 | _T_6297; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6308 = _T_4619 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6309 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6311 = _T_6309 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6313 = _T_6311 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6314 = _T_6308 | _T_6313; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6324 = _T_4623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6325 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6327 = _T_6325 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6329 = _T_6327 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6330 = _T_6324 | _T_6329; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6340 = _T_4627 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6341 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6343 = _T_6341 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6345 = _T_6343 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6346 = _T_6340 | _T_6345; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6356 = _T_4631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6357 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6359 = _T_6357 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6361 = _T_6359 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6362 = _T_6356 | _T_6361; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6372 = _T_4635 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6373 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6375 = _T_6373 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6377 = _T_6375 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6378 = _T_6372 | _T_6377; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6388 = _T_4639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6389 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6391 = _T_6389 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6393 = _T_6391 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6394 = _T_6388 | _T_6393; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6404 = _T_4643 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6405 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6407 = _T_6405 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6409 = _T_6407 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6410 = _T_6404 | _T_6409; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6420 = _T_4647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6421 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6423 = _T_6421 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6425 = _T_6423 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6426 = _T_6420 | _T_6425; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6436 = _T_4651 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6437 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6439 = _T_6437 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6441 = _T_6439 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6442 = _T_6436 | _T_6441; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6452 = _T_4655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6453 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6455 = _T_6453 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6457 = _T_6455 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6458 = _T_6452 | _T_6457; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6468 = _T_4659 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6469 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6471 = _T_6469 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6473 = _T_6471 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6474 = _T_6468 | _T_6473; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6484 = _T_4663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6485 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6487 = _T_6485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6489 = _T_6487 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6490 = _T_6484 | _T_6489; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6500 = _T_4667 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6501 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6503 = _T_6501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6505 = _T_6503 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6506 = _T_6500 | _T_6505; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6516 = _T_4671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6517 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6519 = _T_6517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6521 = _T_6519 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6522 = _T_6516 | _T_6521; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6532 = _T_4675 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6533 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6535 = _T_6533 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6537 = _T_6535 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6538 = _T_6532 | _T_6537; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6548 = _T_4679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6549 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6551 = _T_6549 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6553 = _T_6551 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6554 = _T_6548 | _T_6553; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6564 = _T_4683 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6565 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6567 = _T_6565 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6569 = _T_6567 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6570 = _T_6564 | _T_6569; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6580 = _T_4687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6581 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6583 = _T_6581 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6585 = _T_6583 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6586 = _T_6580 | _T_6585; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6596 = _T_4691 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6597 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6599 = _T_6597 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6601 = _T_6599 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6602 = _T_6596 | _T_6601; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6612 = _T_4695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6613 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6615 = _T_6613 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6617 = _T_6615 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6618 = _T_6612 | _T_6617; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6628 = _T_4699 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6629 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6631 = _T_6629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6633 = _T_6631 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6634 = _T_6628 | _T_6633; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6644 = _T_4703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6645 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6647 = _T_6645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6649 = _T_6647 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6650 = _T_6644 | _T_6649; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6660 = _T_4707 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6661 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6663 = _T_6661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6665 = _T_6663 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6666 = _T_6660 | _T_6665; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6676 = _T_4711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6677 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6679 = _T_6677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6681 = _T_6679 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6682 = _T_6676 | _T_6681; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6692 = _T_4715 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6693 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6695 = _T_6693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6697 = _T_6695 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6698 = _T_6692 | _T_6697; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6708 = _T_4719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6709 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6711 = _T_6709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6713 = _T_6711 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6714 = _T_6708 | _T_6713; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6724 = _T_4723 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6725 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_6727 = _T_6725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6729 = _T_6727 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6730 = _T_6724 | _T_6729; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6740 = _T_4599 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6743 = _T_6229 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6745 = _T_6743 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6746 = _T_6740 | _T_6745; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6756 = _T_4603 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6759 = _T_6245 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6761 = _T_6759 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6762 = _T_6756 | _T_6761; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6772 = _T_4607 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6775 = _T_6261 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6777 = _T_6775 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6778 = _T_6772 | _T_6777; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6788 = _T_4611 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6791 = _T_6277 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6793 = _T_6791 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6794 = _T_6788 | _T_6793; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6804 = _T_4615 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6807 = _T_6293 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6809 = _T_6807 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6810 = _T_6804 | _T_6809; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6820 = _T_4619 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6823 = _T_6309 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6825 = _T_6823 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6826 = _T_6820 | _T_6825; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6836 = _T_4623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6839 = _T_6325 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6841 = _T_6839 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6842 = _T_6836 | _T_6841; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6852 = _T_4627 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6855 = _T_6341 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6857 = _T_6855 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6858 = _T_6852 | _T_6857; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6868 = _T_4631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6871 = _T_6357 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6873 = _T_6871 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6874 = _T_6868 | _T_6873; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6884 = _T_4635 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6887 = _T_6373 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6889 = _T_6887 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6890 = _T_6884 | _T_6889; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6900 = _T_4639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6903 = _T_6389 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6905 = _T_6903 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6906 = _T_6900 | _T_6905; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6916 = _T_4643 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6919 = _T_6405 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6921 = _T_6919 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6922 = _T_6916 | _T_6921; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6932 = _T_4647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6935 = _T_6421 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6937 = _T_6935 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6938 = _T_6932 | _T_6937; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6948 = _T_4651 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6951 = _T_6437 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6953 = _T_6951 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6954 = _T_6948 | _T_6953; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6964 = _T_4655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6967 = _T_6453 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6969 = _T_6967 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6970 = _T_6964 | _T_6969; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6980 = _T_4659 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6983 = _T_6469 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_6985 = _T_6983 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_6986 = _T_6980 | _T_6985; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_6996 = _T_4663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_6999 = _T_6485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7001 = _T_6999 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7002 = _T_6996 | _T_7001; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7012 = _T_4667 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7015 = _T_6501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7017 = _T_7015 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7018 = _T_7012 | _T_7017; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7028 = _T_4671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7031 = _T_6517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7033 = _T_7031 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7034 = _T_7028 | _T_7033; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7044 = _T_4675 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7047 = _T_6533 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7049 = _T_7047 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7050 = _T_7044 | _T_7049; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7060 = _T_4679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7063 = _T_6549 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7065 = _T_7063 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7066 = _T_7060 | _T_7065; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7076 = _T_4683 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7079 = _T_6565 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7081 = _T_7079 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7082 = _T_7076 | _T_7081; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7092 = _T_4687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7095 = _T_6581 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7097 = _T_7095 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7098 = _T_7092 | _T_7097; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7108 = _T_4691 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7111 = _T_6597 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7113 = _T_7111 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7114 = _T_7108 | _T_7113; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7124 = _T_4695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7127 = _T_6613 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7129 = _T_7127 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7130 = _T_7124 | _T_7129; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7140 = _T_4699 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7143 = _T_6629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7145 = _T_7143 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7146 = _T_7140 | _T_7145; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7156 = _T_4703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7159 = _T_6645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7161 = _T_7159 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7162 = _T_7156 | _T_7161; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7172 = _T_4707 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7175 = _T_6661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7177 = _T_7175 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7178 = _T_7172 | _T_7177; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7188 = _T_4711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7191 = _T_6677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7193 = _T_7191 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7194 = _T_7188 | _T_7193; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7204 = _T_4715 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7207 = _T_6693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7209 = _T_7207 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7210 = _T_7204 | _T_7209; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7220 = _T_4719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7223 = _T_6709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7225 = _T_7223 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7226 = _T_7220 | _T_7225; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7236 = _T_4723 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7239 = _T_6725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7241 = _T_7239 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7242 = _T_7236 | _T_7241; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7252 = _T_4727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7253 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7255 = _T_7253 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7257 = _T_7255 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7258 = _T_7252 | _T_7257; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7268 = _T_4731 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7269 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7271 = _T_7269 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7273 = _T_7271 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7274 = _T_7268 | _T_7273; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7284 = _T_4735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7285 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7287 = _T_7285 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7289 = _T_7287 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7290 = _T_7284 | _T_7289; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7300 = _T_4739 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7301 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7303 = _T_7301 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7305 = _T_7303 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7306 = _T_7300 | _T_7305; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7316 = _T_4743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7317 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7319 = _T_7317 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7321 = _T_7319 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7322 = _T_7316 | _T_7321; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7332 = _T_4747 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7333 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7335 = _T_7333 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7337 = _T_7335 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7338 = _T_7332 | _T_7337; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7348 = _T_4751 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7349 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7351 = _T_7349 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7353 = _T_7351 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7354 = _T_7348 | _T_7353; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7364 = _T_4755 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7365 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7367 = _T_7365 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7369 = _T_7367 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7370 = _T_7364 | _T_7369; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7380 = _T_4759 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7381 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7383 = _T_7381 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7385 = _T_7383 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7386 = _T_7380 | _T_7385; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7396 = _T_4763 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7397 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7399 = _T_7397 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7401 = _T_7399 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7402 = _T_7396 | _T_7401; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7412 = _T_4767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7413 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7415 = _T_7413 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7417 = _T_7415 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7418 = _T_7412 | _T_7417; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7428 = _T_4771 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7429 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7431 = _T_7429 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7433 = _T_7431 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7434 = _T_7428 | _T_7433; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7444 = _T_4775 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7445 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7447 = _T_7445 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7449 = _T_7447 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7450 = _T_7444 | _T_7449; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7460 = _T_4779 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7461 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7463 = _T_7461 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7465 = _T_7463 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7466 = _T_7460 | _T_7465; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7476 = _T_4783 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7477 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7479 = _T_7477 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7481 = _T_7479 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7482 = _T_7476 | _T_7481; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7492 = _T_4787 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7493 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7495 = _T_7493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7497 = _T_7495 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7498 = _T_7492 | _T_7497; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7508 = _T_4791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7509 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7511 = _T_7509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7513 = _T_7511 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7514 = _T_7508 | _T_7513; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7524 = _T_4795 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7525 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7527 = _T_7525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7529 = _T_7527 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7530 = _T_7524 | _T_7529; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7540 = _T_4799 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7541 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7543 = _T_7541 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7545 = _T_7543 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7546 = _T_7540 | _T_7545; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7556 = _T_4803 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7557 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7559 = _T_7557 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7561 = _T_7559 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7562 = _T_7556 | _T_7561; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7572 = _T_4807 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7573 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7575 = _T_7573 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7577 = _T_7575 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7578 = _T_7572 | _T_7577; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7588 = _T_4811 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7589 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7591 = _T_7589 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7593 = _T_7591 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7594 = _T_7588 | _T_7593; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7604 = _T_4815 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7605 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7607 = _T_7605 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7609 = _T_7607 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7610 = _T_7604 | _T_7609; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7620 = _T_4819 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7621 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7623 = _T_7621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7625 = _T_7623 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7626 = _T_7620 | _T_7625; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7636 = _T_4823 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7637 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7639 = _T_7637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7641 = _T_7639 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7642 = _T_7636 | _T_7641; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7652 = _T_4827 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7653 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7655 = _T_7653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7657 = _T_7655 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7658 = _T_7652 | _T_7657; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7668 = _T_4831 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7669 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7671 = _T_7669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7673 = _T_7671 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7674 = _T_7668 | _T_7673; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7684 = _T_4835 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7685 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7687 = _T_7685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7689 = _T_7687 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7690 = _T_7684 | _T_7689; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7700 = _T_4839 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7701 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7703 = _T_7701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7705 = _T_7703 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7706 = _T_7700 | _T_7705; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7716 = _T_4843 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7717 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7719 = _T_7717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7721 = _T_7719 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7722 = _T_7716 | _T_7721; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7732 = _T_4847 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7733 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7735 = _T_7733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7737 = _T_7735 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7738 = _T_7732 | _T_7737; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7748 = _T_4851 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7749 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_7751 = _T_7749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7753 = _T_7751 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7754 = _T_7748 | _T_7753; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7764 = _T_4727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7767 = _T_7253 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7769 = _T_7767 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7770 = _T_7764 | _T_7769; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7780 = _T_4731 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7783 = _T_7269 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7785 = _T_7783 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7786 = _T_7780 | _T_7785; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7796 = _T_4735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7799 = _T_7285 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7801 = _T_7799 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7802 = _T_7796 | _T_7801; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7812 = _T_4739 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7815 = _T_7301 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7817 = _T_7815 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7818 = _T_7812 | _T_7817; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7828 = _T_4743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7831 = _T_7317 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7833 = _T_7831 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7834 = _T_7828 | _T_7833; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7844 = _T_4747 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7847 = _T_7333 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7849 = _T_7847 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7850 = _T_7844 | _T_7849; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7860 = _T_4751 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7863 = _T_7349 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7865 = _T_7863 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7866 = _T_7860 | _T_7865; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7876 = _T_4755 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7879 = _T_7365 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7881 = _T_7879 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7882 = _T_7876 | _T_7881; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7892 = _T_4759 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7895 = _T_7381 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7897 = _T_7895 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7898 = _T_7892 | _T_7897; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7908 = _T_4763 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7911 = _T_7397 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7913 = _T_7911 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7914 = _T_7908 | _T_7913; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7924 = _T_4767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7927 = _T_7413 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7929 = _T_7927 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7930 = _T_7924 | _T_7929; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7940 = _T_4771 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7943 = _T_7429 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7945 = _T_7943 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7946 = _T_7940 | _T_7945; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7956 = _T_4775 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7959 = _T_7445 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7961 = _T_7959 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7962 = _T_7956 | _T_7961; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7972 = _T_4779 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7975 = _T_7461 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7977 = _T_7975 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7978 = _T_7972 | _T_7977; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_7988 = _T_4783 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_7991 = _T_7477 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_7993 = _T_7991 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_7994 = _T_7988 | _T_7993; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8004 = _T_4787 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8007 = _T_7493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8009 = _T_8007 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8010 = _T_8004 | _T_8009; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8020 = _T_4791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8023 = _T_7509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8025 = _T_8023 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8026 = _T_8020 | _T_8025; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8036 = _T_4795 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8039 = _T_7525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8041 = _T_8039 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8042 = _T_8036 | _T_8041; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8052 = _T_4799 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8055 = _T_7541 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8057 = _T_8055 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8058 = _T_8052 | _T_8057; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8068 = _T_4803 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8071 = _T_7557 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8073 = _T_8071 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8074 = _T_8068 | _T_8073; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8084 = _T_4807 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8087 = _T_7573 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8089 = _T_8087 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8090 = _T_8084 | _T_8089; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8100 = _T_4811 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8103 = _T_7589 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8105 = _T_8103 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8106 = _T_8100 | _T_8105; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8116 = _T_4815 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8119 = _T_7605 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8121 = _T_8119 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8122 = _T_8116 | _T_8121; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8132 = _T_4819 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8135 = _T_7621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8137 = _T_8135 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8138 = _T_8132 | _T_8137; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8148 = _T_4823 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8151 = _T_7637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8153 = _T_8151 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8154 = _T_8148 | _T_8153; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8164 = _T_4827 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8167 = _T_7653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8169 = _T_8167 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8170 = _T_8164 | _T_8169; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8180 = _T_4831 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8183 = _T_7669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8185 = _T_8183 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8186 = _T_8180 | _T_8185; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8196 = _T_4835 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8199 = _T_7685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8201 = _T_8199 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8202 = _T_8196 | _T_8201; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8212 = _T_4839 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8215 = _T_7701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8217 = _T_8215 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8218 = _T_8212 | _T_8217; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8228 = _T_4843 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8231 = _T_7717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8233 = _T_8231 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8234 = _T_8228 | _T_8233; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8244 = _T_4847 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8247 = _T_7733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8249 = _T_8247 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8250 = _T_8244 | _T_8249; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8260 = _T_4851 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8263 = _T_7749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8265 = _T_8263 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8266 = _T_8260 | _T_8265; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8276 = _T_4855 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8277 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8279 = _T_8277 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8281 = _T_8279 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8282 = _T_8276 | _T_8281; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8292 = _T_4859 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8293 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8295 = _T_8293 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8297 = _T_8295 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8298 = _T_8292 | _T_8297; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8308 = _T_4863 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8309 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8311 = _T_8309 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8313 = _T_8311 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8314 = _T_8308 | _T_8313; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8324 = _T_4867 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8325 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8327 = _T_8325 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8329 = _T_8327 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8330 = _T_8324 | _T_8329; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8340 = _T_4871 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8341 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8343 = _T_8341 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8345 = _T_8343 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8346 = _T_8340 | _T_8345; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8356 = _T_4875 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8357 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8359 = _T_8357 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8361 = _T_8359 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8362 = _T_8356 | _T_8361; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8372 = _T_4879 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8373 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8375 = _T_8373 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8377 = _T_8375 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8378 = _T_8372 | _T_8377; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8388 = _T_4883 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8389 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8391 = _T_8389 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8393 = _T_8391 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8394 = _T_8388 | _T_8393; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8404 = _T_4887 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8405 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8407 = _T_8405 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8409 = _T_8407 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8410 = _T_8404 | _T_8409; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8420 = _T_4891 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8421 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8423 = _T_8421 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8425 = _T_8423 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8426 = _T_8420 | _T_8425; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8436 = _T_4895 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8437 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8439 = _T_8437 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8441 = _T_8439 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8442 = _T_8436 | _T_8441; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8452 = _T_4899 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8453 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8455 = _T_8453 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8457 = _T_8455 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8458 = _T_8452 | _T_8457; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8468 = _T_4903 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8469 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8471 = _T_8469 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8473 = _T_8471 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8474 = _T_8468 | _T_8473; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8484 = _T_4907 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8485 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8487 = _T_8485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8489 = _T_8487 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8490 = _T_8484 | _T_8489; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8500 = _T_4911 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8501 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8503 = _T_8501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8505 = _T_8503 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8506 = _T_8500 | _T_8505; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8516 = _T_4915 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8517 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8519 = _T_8517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8521 = _T_8519 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8522 = _T_8516 | _T_8521; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8532 = _T_4919 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8533 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8535 = _T_8533 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8537 = _T_8535 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8538 = _T_8532 | _T_8537; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8548 = _T_4923 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8549 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8551 = _T_8549 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8553 = _T_8551 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8554 = _T_8548 | _T_8553; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8564 = _T_4927 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8565 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8567 = _T_8565 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8569 = _T_8567 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8570 = _T_8564 | _T_8569; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8580 = _T_4931 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8581 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8583 = _T_8581 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8585 = _T_8583 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8586 = _T_8580 | _T_8585; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8596 = _T_4935 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8597 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8599 = _T_8597 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8601 = _T_8599 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8602 = _T_8596 | _T_8601; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8612 = _T_4939 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8613 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8615 = _T_8613 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8617 = _T_8615 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8618 = _T_8612 | _T_8617; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8628 = _T_4943 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8629 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8631 = _T_8629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8633 = _T_8631 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8634 = _T_8628 | _T_8633; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8644 = _T_4947 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8645 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8647 = _T_8645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8649 = _T_8647 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8650 = _T_8644 | _T_8649; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8660 = _T_4951 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8661 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8663 = _T_8661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8665 = _T_8663 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8666 = _T_8660 | _T_8665; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8676 = _T_4955 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8677 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8679 = _T_8677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8681 = _T_8679 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8682 = _T_8676 | _T_8681; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8692 = _T_4959 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8693 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8695 = _T_8693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8697 = _T_8695 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8698 = _T_8692 | _T_8697; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8708 = _T_4963 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8709 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8711 = _T_8709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8713 = _T_8711 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8714 = _T_8708 | _T_8713; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8724 = _T_4967 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8725 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8727 = _T_8725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8729 = _T_8727 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8730 = _T_8724 | _T_8729; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8740 = _T_4971 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8741 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8743 = _T_8741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8745 = _T_8743 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8746 = _T_8740 | _T_8745; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8756 = _T_4975 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8757 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8759 = _T_8757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8761 = _T_8759 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8762 = _T_8756 | _T_8761; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8772 = _T_4979 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8773 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 742:101]
  wire  _T_8775 = _T_8773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8777 = _T_8775 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8778 = _T_8772 | _T_8777; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8788 = _T_4855 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8791 = _T_8277 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8793 = _T_8791 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8794 = _T_8788 | _T_8793; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8804 = _T_4859 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8807 = _T_8293 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8809 = _T_8807 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8810 = _T_8804 | _T_8809; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8820 = _T_4863 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8823 = _T_8309 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8825 = _T_8823 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8826 = _T_8820 | _T_8825; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8836 = _T_4867 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8839 = _T_8325 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8841 = _T_8839 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8842 = _T_8836 | _T_8841; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8852 = _T_4871 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8855 = _T_8341 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8857 = _T_8855 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8858 = _T_8852 | _T_8857; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8868 = _T_4875 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8871 = _T_8357 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8873 = _T_8871 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8874 = _T_8868 | _T_8873; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8884 = _T_4879 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8887 = _T_8373 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8889 = _T_8887 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8890 = _T_8884 | _T_8889; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8900 = _T_4883 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8903 = _T_8389 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8905 = _T_8903 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8906 = _T_8900 | _T_8905; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8916 = _T_4887 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8919 = _T_8405 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8921 = _T_8919 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8922 = _T_8916 | _T_8921; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8932 = _T_4891 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8935 = _T_8421 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8937 = _T_8935 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8938 = _T_8932 | _T_8937; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8948 = _T_4895 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8951 = _T_8437 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8953 = _T_8951 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8954 = _T_8948 | _T_8953; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8964 = _T_4899 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8967 = _T_8453 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8969 = _T_8967 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8970 = _T_8964 | _T_8969; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8980 = _T_4903 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8983 = _T_8469 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_8985 = _T_8983 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_8986 = _T_8980 | _T_8985; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_8996 = _T_4907 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_8999 = _T_8485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9001 = _T_8999 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9002 = _T_8996 | _T_9001; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9012 = _T_4911 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9015 = _T_8501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9017 = _T_9015 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9018 = _T_9012 | _T_9017; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9028 = _T_4915 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9031 = _T_8517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9033 = _T_9031 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9034 = _T_9028 | _T_9033; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9044 = _T_4919 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9047 = _T_8533 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9049 = _T_9047 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9050 = _T_9044 | _T_9049; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9060 = _T_4923 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9063 = _T_8549 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9065 = _T_9063 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9066 = _T_9060 | _T_9065; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9076 = _T_4927 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9079 = _T_8565 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9081 = _T_9079 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9082 = _T_9076 | _T_9081; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9092 = _T_4931 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9095 = _T_8581 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9097 = _T_9095 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9098 = _T_9092 | _T_9097; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9108 = _T_4935 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9111 = _T_8597 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9113 = _T_9111 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9114 = _T_9108 | _T_9113; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9124 = _T_4939 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9127 = _T_8613 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9129 = _T_9127 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9130 = _T_9124 | _T_9129; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9140 = _T_4943 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9143 = _T_8629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9145 = _T_9143 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9146 = _T_9140 | _T_9145; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9156 = _T_4947 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9159 = _T_8645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9161 = _T_9159 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9162 = _T_9156 | _T_9161; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9172 = _T_4951 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9175 = _T_8661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9177 = _T_9175 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9178 = _T_9172 | _T_9177; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9188 = _T_4955 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9191 = _T_8677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9193 = _T_9191 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9194 = _T_9188 | _T_9193; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9204 = _T_4959 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9207 = _T_8693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9209 = _T_9207 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9210 = _T_9204 | _T_9209; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9220 = _T_4963 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9223 = _T_8709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9225 = _T_9223 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9226 = _T_9220 | _T_9225; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9236 = _T_4967 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9239 = _T_8725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9241 = _T_9239 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9242 = _T_9236 | _T_9241; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9252 = _T_4971 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9255 = _T_8741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9257 = _T_9255 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9258 = _T_9252 | _T_9257; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9268 = _T_4975 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9271 = _T_8757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9273 = _T_9271 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9274 = _T_9268 | _T_9273; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_9284 = _T_4979 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:58]
  wire  _T_9287 = _T_8773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 742:123]
  wire  _T_9289 = _T_9287 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 742:144]
  wire  _T_9290 = _T_9284 | _T_9289; // @[el2_ifu_mem_ctl.scala 742:80]
  wire  _T_10091 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 796:63]
  wire  _T_10092 = _T_10091 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 796:85]
  wire [1:0] _T_10094 = _T_10092 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10101; // @[el2_ifu_mem_ctl.scala 801:57]
  reg  _T_10102; // @[el2_ifu_mem_ctl.scala 802:56]
  reg  _T_10103; // @[el2_ifu_mem_ctl.scala 803:59]
  wire  _T_10104 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 804:80]
  wire  _T_10105 = ifu_bus_arvalid_ff & _T_10104; // @[el2_ifu_mem_ctl.scala 804:78]
  wire  _T_10106 = _T_10105 & miss_pending; // @[el2_ifu_mem_ctl.scala 804:100]
  reg  _T_10107; // @[el2_ifu_mem_ctl.scala 804:58]
  reg  _T_10108; // @[el2_ifu_mem_ctl.scala 805:58]
  wire  _T_10111 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 812:71]
  wire  _T_10113 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 812:124]
  wire  _T_10115 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 813:50]
  wire  _T_10117 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 813:103]
  wire [3:0] _T_10120 = {_T_10111,_T_10113,_T_10115,_T_10117}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 815:53]
  reg  _T_10131; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 324:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 323:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 187:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3926; // @[el2_ifu_mem_ctl.scala 692:21]
  assign io_ifu_pmu_ic_miss = _T_10101; // @[el2_ifu_mem_ctl.scala 801:22]
  assign io_ifu_pmu_ic_hit = _T_10102; // @[el2_ifu_mem_ctl.scala 802:21]
  assign io_ifu_pmu_bus_error = _T_10103; // @[el2_ifu_mem_ctl.scala 803:24]
  assign io_ifu_pmu_bus_busy = _T_10107; // @[el2_ifu_mem_ctl.scala 804:23]
  assign io_ifu_pmu_bus_trxn = _T_10108; // @[el2_ifu_mem_ctl.scala 805:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 138:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 137:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 132:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 136:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 145:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 147:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 142:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 140:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 131:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 129:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 130:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 143:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 554:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2520; // @[el2_ifu_mem_ctl.scala 555:19]
  assign io_ifu_axi_araddr = _T_2522 & _T_2524; // @[el2_ifu_mem_ctl.scala 556:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 559:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 557:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 560:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 135:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 558:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 141:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 561:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 651:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 649:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 653:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 644:20]
  assign io_iccm_ready = _T_2623 & _T_2617; // @[el2_ifu_mem_ctl.scala 624:17]
  assign io_ic_rw_addr = _T_340 | _T_341; // @[el2_ifu_mem_ctl.scala 333:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 691:15]
  assign io_ic_rd_en = _T_3904 | _T_3909; // @[el2_ifu_mem_ctl.scala 682:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 340:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 340:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 341:23]
  assign io_ifu_ic_debug_rd_data = _T_1211; // @[el2_ifu_mem_ctl.scala 349:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 808:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 810:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 811:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 809:25]
  assign io_ic_debug_way = _T_10120[1:0]; // @[el2_ifu_mem_ctl.scala 812:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10094; // @[el2_ifu_mem_ctl.scala 796:19]
  assign io_iccm_rw_addr = _T_3058[14:0]; // @[el2_ifu_mem_ctl.scala 655:19]
  assign io_iccm_wren = _T_2627 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 626:16]
  assign io_iccm_rden = _T_2631 | _T_2632; // @[el2_ifu_mem_ctl.scala 627:16]
  assign io_iccm_wr_data = _T_3033 ? _T_3034 : _T_3041; // @[el2_ifu_mem_ctl.scala 632:19]
  assign io_iccm_wr_size = _T_2637 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 629:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 285:15]
  assign io_ic_access_fault_f = _T_2405 & _T_317; // @[el2_ifu_mem_ctl.scala 380:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1275; // @[el2_ifu_mem_ctl.scala 381:29]
  assign io_iccm_rd_ecc_single_err = _T_3849 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 668:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 669:29]
  assign io_ic_error_start = _T_1199 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 343:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 186:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 185:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 385:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 377:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 374:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 375:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10131; // @[el2_ifu_mem_ctl.scala 819:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2410; // @[el2_ifu_mem_ctl.scala 473:27]
  assign io_iccm_correction_state = _T_2438 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 508:28 el2_ifu_mem_ctl.scala 521:32 el2_ifu_mem_ctl.scala 528:32 el2_ifu_mem_ctl.scala 535:32]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_5114 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4470 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4466 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4462 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4458 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4454 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4450 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4446 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4442 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4438 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4434 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4430 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4426 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4422 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4418 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4414 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4410 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4406 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4402 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4398 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4394 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4390 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4386 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4382 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4378 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4374 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4370 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4366 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4362 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4358 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4354 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4350 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4346 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4342 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4338 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4334 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4330 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4326 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4322 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4318 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4314 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4310 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4306 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4302 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4298 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4294 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4290 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4286 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4282 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_4278 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_4274 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_4270 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_4266 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_4262 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_4258 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_4254 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_4250 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_4246 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_4242 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4238 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4234 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4230 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4226 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_4222 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_4218 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_4214 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_4210 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4206 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4202 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4198 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4194 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4190 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4186 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4182 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4178 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_4174 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4170 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_4166 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_4162 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_4158 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_4154 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_4150 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_4146 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_4142 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_4138 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_4134 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_4130 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_4126 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_4122 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_4118 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_4114 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_4110 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_4106 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_4102 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_4098 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_4094 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_4090 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_4086 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_4082 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_4078 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_4074 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_4070 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_4066 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_4062 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_4058 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_4054 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_4050 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_4046 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4042 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4038 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4034 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4030 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_4026 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_4022 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_4018 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_4014 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_4010 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_4006 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_4002 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3998 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3994 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3990 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3986 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3982 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3978 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3974 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3970 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3966 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3962 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  _T_1295 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  _T_1297 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  _T_1299 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  _T_1301 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  _T_1303 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  _T_1305 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  _T_1307 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  _T_1309 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  _T_1311 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  _T_1313 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  _T_1315 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  _T_1317 = _RAND_175[63:0];
  _RAND_176 = {2{`RANDOM}};
  _T_1319 = _RAND_176[63:0];
  _RAND_177 = {2{`RANDOM}};
  _T_1321 = _RAND_177[63:0];
  _RAND_178 = {2{`RANDOM}};
  _T_1323 = _RAND_178[63:0];
  _RAND_179 = {2{`RANDOM}};
  _T_1325 = _RAND_179[63:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_1211 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_10101 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10102 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10103 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10107 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10108 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10131 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_4470 <= 3'h0;
    end else if (_T_4469) begin
      _T_4470 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4466 <= 3'h0;
    end else if (_T_4465) begin
      _T_4466 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4462 <= 3'h0;
    end else if (_T_4461) begin
      _T_4462 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4458 <= 3'h0;
    end else if (_T_4457) begin
      _T_4458 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4454 <= 3'h0;
    end else if (_T_4453) begin
      _T_4454 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4450 <= 3'h0;
    end else if (_T_4449) begin
      _T_4450 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4446 <= 3'h0;
    end else if (_T_4445) begin
      _T_4446 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4442 <= 3'h0;
    end else if (_T_4441) begin
      _T_4442 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4438 <= 3'h0;
    end else if (_T_4437) begin
      _T_4438 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4434 <= 3'h0;
    end else if (_T_4433) begin
      _T_4434 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4430 <= 3'h0;
    end else if (_T_4429) begin
      _T_4430 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4426 <= 3'h0;
    end else if (_T_4425) begin
      _T_4426 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4422 <= 3'h0;
    end else if (_T_4421) begin
      _T_4422 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4418 <= 3'h0;
    end else if (_T_4417) begin
      _T_4418 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4414 <= 3'h0;
    end else if (_T_4413) begin
      _T_4414 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4410 <= 3'h0;
    end else if (_T_4409) begin
      _T_4410 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4406 <= 3'h0;
    end else if (_T_4405) begin
      _T_4406 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4402 <= 3'h0;
    end else if (_T_4401) begin
      _T_4402 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4398 <= 3'h0;
    end else if (_T_4397) begin
      _T_4398 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4394 <= 3'h0;
    end else if (_T_4393) begin
      _T_4394 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4390 <= 3'h0;
    end else if (_T_4389) begin
      _T_4390 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4386 <= 3'h0;
    end else if (_T_4385) begin
      _T_4386 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4382 <= 3'h0;
    end else if (_T_4381) begin
      _T_4382 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4378 <= 3'h0;
    end else if (_T_4377) begin
      _T_4378 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4374 <= 3'h0;
    end else if (_T_4373) begin
      _T_4374 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4370 <= 3'h0;
    end else if (_T_4369) begin
      _T_4370 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4366 <= 3'h0;
    end else if (_T_4365) begin
      _T_4366 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4362 <= 3'h0;
    end else if (_T_4361) begin
      _T_4362 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4358 <= 3'h0;
    end else if (_T_4357) begin
      _T_4358 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4354 <= 3'h0;
    end else if (_T_4353) begin
      _T_4354 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4350 <= 3'h0;
    end else if (_T_4349) begin
      _T_4350 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4346 <= 3'h0;
    end else if (_T_4345) begin
      _T_4346 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4342 <= 3'h0;
    end else if (_T_4341) begin
      _T_4342 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4338 <= 3'h0;
    end else if (_T_4337) begin
      _T_4338 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4334 <= 3'h0;
    end else if (_T_4333) begin
      _T_4334 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4330 <= 3'h0;
    end else if (_T_4329) begin
      _T_4330 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4326 <= 3'h0;
    end else if (_T_4325) begin
      _T_4326 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4322 <= 3'h0;
    end else if (_T_4321) begin
      _T_4322 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4318 <= 3'h0;
    end else if (_T_4317) begin
      _T_4318 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4314 <= 3'h0;
    end else if (_T_4313) begin
      _T_4314 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4310 <= 3'h0;
    end else if (_T_4309) begin
      _T_4310 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4306 <= 3'h0;
    end else if (_T_4305) begin
      _T_4306 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4302 <= 3'h0;
    end else if (_T_4301) begin
      _T_4302 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4298 <= 3'h0;
    end else if (_T_4297) begin
      _T_4298 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4294 <= 3'h0;
    end else if (_T_4293) begin
      _T_4294 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4290 <= 3'h0;
    end else if (_T_4289) begin
      _T_4290 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4286 <= 3'h0;
    end else if (_T_4285) begin
      _T_4286 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4282 <= 3'h0;
    end else if (_T_4281) begin
      _T_4282 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4278 <= 3'h0;
    end else if (_T_4277) begin
      _T_4278 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4274 <= 3'h0;
    end else if (_T_4273) begin
      _T_4274 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4270 <= 3'h0;
    end else if (_T_4269) begin
      _T_4270 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4266 <= 3'h0;
    end else if (_T_4265) begin
      _T_4266 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4262 <= 3'h0;
    end else if (_T_4261) begin
      _T_4262 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4258 <= 3'h0;
    end else if (_T_4257) begin
      _T_4258 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4254 <= 3'h0;
    end else if (_T_4253) begin
      _T_4254 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4250 <= 3'h0;
    end else if (_T_4249) begin
      _T_4250 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4246 <= 3'h0;
    end else if (_T_4245) begin
      _T_4246 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4242 <= 3'h0;
    end else if (_T_4241) begin
      _T_4242 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4238 <= 3'h0;
    end else if (_T_4237) begin
      _T_4238 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4234 <= 3'h0;
    end else if (_T_4233) begin
      _T_4234 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4230 <= 3'h0;
    end else if (_T_4229) begin
      _T_4230 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4226 <= 3'h0;
    end else if (_T_4225) begin
      _T_4226 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4222 <= 3'h0;
    end else if (_T_4221) begin
      _T_4222 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4218 <= 3'h0;
    end else if (_T_4217) begin
      _T_4218 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4214 <= 3'h0;
    end else if (_T_4213) begin
      _T_4214 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4210 <= 3'h0;
    end else if (_T_4209) begin
      _T_4210 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4206 <= 3'h0;
    end else if (_T_4205) begin
      _T_4206 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4202 <= 3'h0;
    end else if (_T_4201) begin
      _T_4202 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4198 <= 3'h0;
    end else if (_T_4197) begin
      _T_4198 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4194 <= 3'h0;
    end else if (_T_4193) begin
      _T_4194 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4190 <= 3'h0;
    end else if (_T_4189) begin
      _T_4190 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4186 <= 3'h0;
    end else if (_T_4185) begin
      _T_4186 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4182 <= 3'h0;
    end else if (_T_4181) begin
      _T_4182 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4178 <= 3'h0;
    end else if (_T_4177) begin
      _T_4178 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4174 <= 3'h0;
    end else if (_T_4173) begin
      _T_4174 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4170 <= 3'h0;
    end else if (_T_4169) begin
      _T_4170 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4166 <= 3'h0;
    end else if (_T_4165) begin
      _T_4166 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4162 <= 3'h0;
    end else if (_T_4161) begin
      _T_4162 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4158 <= 3'h0;
    end else if (_T_4157) begin
      _T_4158 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4154 <= 3'h0;
    end else if (_T_4153) begin
      _T_4154 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4150 <= 3'h0;
    end else if (_T_4149) begin
      _T_4150 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4146 <= 3'h0;
    end else if (_T_4145) begin
      _T_4146 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4142 <= 3'h0;
    end else if (_T_4141) begin
      _T_4142 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4138 <= 3'h0;
    end else if (_T_4137) begin
      _T_4138 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4134 <= 3'h0;
    end else if (_T_4133) begin
      _T_4134 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4130 <= 3'h0;
    end else if (_T_4129) begin
      _T_4130 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4126 <= 3'h0;
    end else if (_T_4125) begin
      _T_4126 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4122 <= 3'h0;
    end else if (_T_4121) begin
      _T_4122 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4118 <= 3'h0;
    end else if (_T_4117) begin
      _T_4118 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4114 <= 3'h0;
    end else if (_T_4113) begin
      _T_4114 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4110 <= 3'h0;
    end else if (_T_4109) begin
      _T_4110 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4106 <= 3'h0;
    end else if (_T_4105) begin
      _T_4106 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4102 <= 3'h0;
    end else if (_T_4101) begin
      _T_4102 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4098 <= 3'h0;
    end else if (_T_4097) begin
      _T_4098 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4094 <= 3'h0;
    end else if (_T_4093) begin
      _T_4094 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4090 <= 3'h0;
    end else if (_T_4089) begin
      _T_4090 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4086 <= 3'h0;
    end else if (_T_4085) begin
      _T_4086 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4082 <= 3'h0;
    end else if (_T_4081) begin
      _T_4082 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4078 <= 3'h0;
    end else if (_T_4077) begin
      _T_4078 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4074 <= 3'h0;
    end else if (_T_4073) begin
      _T_4074 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4070 <= 3'h0;
    end else if (_T_4069) begin
      _T_4070 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4066 <= 3'h0;
    end else if (_T_4065) begin
      _T_4066 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4062 <= 3'h0;
    end else if (_T_4061) begin
      _T_4062 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4058 <= 3'h0;
    end else if (_T_4057) begin
      _T_4058 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4054 <= 3'h0;
    end else if (_T_4053) begin
      _T_4054 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4050 <= 3'h0;
    end else if (_T_4049) begin
      _T_4050 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4046 <= 3'h0;
    end else if (_T_4045) begin
      _T_4046 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4042 <= 3'h0;
    end else if (_T_4041) begin
      _T_4042 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4038 <= 3'h0;
    end else if (_T_4037) begin
      _T_4038 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4034 <= 3'h0;
    end else if (_T_4033) begin
      _T_4034 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4030 <= 3'h0;
    end else if (_T_4029) begin
      _T_4030 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4026 <= 3'h0;
    end else if (_T_4025) begin
      _T_4026 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4022 <= 3'h0;
    end else if (_T_4021) begin
      _T_4022 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4018 <= 3'h0;
    end else if (_T_4017) begin
      _T_4018 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4014 <= 3'h0;
    end else if (_T_4013) begin
      _T_4014 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4010 <= 3'h0;
    end else if (_T_4009) begin
      _T_4010 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4006 <= 3'h0;
    end else if (_T_4005) begin
      _T_4006 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4002 <= 3'h0;
    end else if (_T_4001) begin
      _T_4002 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3998 <= 3'h0;
    end else if (_T_3997) begin
      _T_3998 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3994 <= 3'h0;
    end else if (_T_3993) begin
      _T_3994 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3990 <= 3'h0;
    end else if (_T_3989) begin
      _T_3990 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3986 <= 3'h0;
    end else if (_T_3985) begin
      _T_3986 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3982 <= 3'h0;
    end else if (_T_3981) begin
      _T_3982 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3978 <= 3'h0;
    end else if (_T_3977) begin
      _T_3978 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3974 <= 3'h0;
    end else if (_T_3973) begin
      _T_3974 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3970 <= 3'h0;
    end else if (_T_3969) begin
      _T_3970 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3966 <= 3'h0;
    end else if (_T_3965) begin
      _T_3966 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3962 <= 3'h0;
    end else if (_T_3961) begin
      _T_3962 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_289;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2563) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2559;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1295 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1295 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1297 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1297 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1299 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1299 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1301 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1301 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1303 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1303 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1305 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1305 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1307 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1307 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1309 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1309 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1311 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1311 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1313 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1313 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1315 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1315 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1317 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1317 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1319 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1319 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1321 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1321 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1323 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1323 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1325 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1325 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5722) begin
      ic_tag_valid_out_1_0 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5738) begin
      ic_tag_valid_out_1_1 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5754) begin
      ic_tag_valid_out_1_2 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5770) begin
      ic_tag_valid_out_1_3 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5786) begin
      ic_tag_valid_out_1_4 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5802) begin
      ic_tag_valid_out_1_5 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5818) begin
      ic_tag_valid_out_1_6 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5834) begin
      ic_tag_valid_out_1_7 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5850) begin
      ic_tag_valid_out_1_8 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5866) begin
      ic_tag_valid_out_1_9 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5882) begin
      ic_tag_valid_out_1_10 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5898) begin
      ic_tag_valid_out_1_11 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5914) begin
      ic_tag_valid_out_1_12 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5930) begin
      ic_tag_valid_out_1_13 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5946) begin
      ic_tag_valid_out_1_14 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5962) begin
      ic_tag_valid_out_1_15 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5978) begin
      ic_tag_valid_out_1_16 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5994) begin
      ic_tag_valid_out_1_17 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6010) begin
      ic_tag_valid_out_1_18 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6026) begin
      ic_tag_valid_out_1_19 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6042) begin
      ic_tag_valid_out_1_20 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6058) begin
      ic_tag_valid_out_1_21 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6074) begin
      ic_tag_valid_out_1_22 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6090) begin
      ic_tag_valid_out_1_23 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6106) begin
      ic_tag_valid_out_1_24 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6122) begin
      ic_tag_valid_out_1_25 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6138) begin
      ic_tag_valid_out_1_26 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6154) begin
      ic_tag_valid_out_1_27 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6170) begin
      ic_tag_valid_out_1_28 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6186) begin
      ic_tag_valid_out_1_29 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6202) begin
      ic_tag_valid_out_1_30 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6218) begin
      ic_tag_valid_out_1_31 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6746) begin
      ic_tag_valid_out_1_32 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6762) begin
      ic_tag_valid_out_1_33 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6778) begin
      ic_tag_valid_out_1_34 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6794) begin
      ic_tag_valid_out_1_35 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6810) begin
      ic_tag_valid_out_1_36 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6826) begin
      ic_tag_valid_out_1_37 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6842) begin
      ic_tag_valid_out_1_38 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6858) begin
      ic_tag_valid_out_1_39 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6874) begin
      ic_tag_valid_out_1_40 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6890) begin
      ic_tag_valid_out_1_41 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6906) begin
      ic_tag_valid_out_1_42 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6922) begin
      ic_tag_valid_out_1_43 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6938) begin
      ic_tag_valid_out_1_44 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6954) begin
      ic_tag_valid_out_1_45 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6970) begin
      ic_tag_valid_out_1_46 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6986) begin
      ic_tag_valid_out_1_47 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7002) begin
      ic_tag_valid_out_1_48 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7018) begin
      ic_tag_valid_out_1_49 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7034) begin
      ic_tag_valid_out_1_50 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7050) begin
      ic_tag_valid_out_1_51 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7066) begin
      ic_tag_valid_out_1_52 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7082) begin
      ic_tag_valid_out_1_53 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7098) begin
      ic_tag_valid_out_1_54 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7114) begin
      ic_tag_valid_out_1_55 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7130) begin
      ic_tag_valid_out_1_56 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7146) begin
      ic_tag_valid_out_1_57 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7162) begin
      ic_tag_valid_out_1_58 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7178) begin
      ic_tag_valid_out_1_59 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7194) begin
      ic_tag_valid_out_1_60 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7210) begin
      ic_tag_valid_out_1_61 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7226) begin
      ic_tag_valid_out_1_62 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7242) begin
      ic_tag_valid_out_1_63 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7770) begin
      ic_tag_valid_out_1_64 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7786) begin
      ic_tag_valid_out_1_65 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7802) begin
      ic_tag_valid_out_1_66 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7818) begin
      ic_tag_valid_out_1_67 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7834) begin
      ic_tag_valid_out_1_68 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7850) begin
      ic_tag_valid_out_1_69 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7866) begin
      ic_tag_valid_out_1_70 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7882) begin
      ic_tag_valid_out_1_71 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7898) begin
      ic_tag_valid_out_1_72 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7914) begin
      ic_tag_valid_out_1_73 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7930) begin
      ic_tag_valid_out_1_74 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7946) begin
      ic_tag_valid_out_1_75 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7962) begin
      ic_tag_valid_out_1_76 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7978) begin
      ic_tag_valid_out_1_77 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7994) begin
      ic_tag_valid_out_1_78 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8010) begin
      ic_tag_valid_out_1_79 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8026) begin
      ic_tag_valid_out_1_80 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8042) begin
      ic_tag_valid_out_1_81 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8058) begin
      ic_tag_valid_out_1_82 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8074) begin
      ic_tag_valid_out_1_83 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8090) begin
      ic_tag_valid_out_1_84 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8106) begin
      ic_tag_valid_out_1_85 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8122) begin
      ic_tag_valid_out_1_86 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8138) begin
      ic_tag_valid_out_1_87 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8154) begin
      ic_tag_valid_out_1_88 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8170) begin
      ic_tag_valid_out_1_89 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8186) begin
      ic_tag_valid_out_1_90 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8202) begin
      ic_tag_valid_out_1_91 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8218) begin
      ic_tag_valid_out_1_92 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8234) begin
      ic_tag_valid_out_1_93 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8250) begin
      ic_tag_valid_out_1_94 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8266) begin
      ic_tag_valid_out_1_95 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8794) begin
      ic_tag_valid_out_1_96 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8810) begin
      ic_tag_valid_out_1_97 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8826) begin
      ic_tag_valid_out_1_98 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8842) begin
      ic_tag_valid_out_1_99 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8858) begin
      ic_tag_valid_out_1_100 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8874) begin
      ic_tag_valid_out_1_101 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8890) begin
      ic_tag_valid_out_1_102 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8906) begin
      ic_tag_valid_out_1_103 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8922) begin
      ic_tag_valid_out_1_104 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8938) begin
      ic_tag_valid_out_1_105 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8954) begin
      ic_tag_valid_out_1_106 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8970) begin
      ic_tag_valid_out_1_107 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8986) begin
      ic_tag_valid_out_1_108 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9002) begin
      ic_tag_valid_out_1_109 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9018) begin
      ic_tag_valid_out_1_110 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9034) begin
      ic_tag_valid_out_1_111 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9050) begin
      ic_tag_valid_out_1_112 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9066) begin
      ic_tag_valid_out_1_113 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9082) begin
      ic_tag_valid_out_1_114 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9098) begin
      ic_tag_valid_out_1_115 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9114) begin
      ic_tag_valid_out_1_116 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9130) begin
      ic_tag_valid_out_1_117 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9146) begin
      ic_tag_valid_out_1_118 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9162) begin
      ic_tag_valid_out_1_119 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9178) begin
      ic_tag_valid_out_1_120 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9194) begin
      ic_tag_valid_out_1_121 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9210) begin
      ic_tag_valid_out_1_122 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9226) begin
      ic_tag_valid_out_1_123 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9242) begin
      ic_tag_valid_out_1_124 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9258) begin
      ic_tag_valid_out_1_125 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9274) begin
      ic_tag_valid_out_1_126 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9290) begin
      ic_tag_valid_out_1_127 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5210) begin
      ic_tag_valid_out_0_0 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5226) begin
      ic_tag_valid_out_0_1 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5242) begin
      ic_tag_valid_out_0_2 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5258) begin
      ic_tag_valid_out_0_3 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5274) begin
      ic_tag_valid_out_0_4 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5290) begin
      ic_tag_valid_out_0_5 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5306) begin
      ic_tag_valid_out_0_6 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5322) begin
      ic_tag_valid_out_0_7 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5338) begin
      ic_tag_valid_out_0_8 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5354) begin
      ic_tag_valid_out_0_9 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5370) begin
      ic_tag_valid_out_0_10 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5386) begin
      ic_tag_valid_out_0_11 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5402) begin
      ic_tag_valid_out_0_12 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5418) begin
      ic_tag_valid_out_0_13 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5434) begin
      ic_tag_valid_out_0_14 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5450) begin
      ic_tag_valid_out_0_15 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5466) begin
      ic_tag_valid_out_0_16 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5482) begin
      ic_tag_valid_out_0_17 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5498) begin
      ic_tag_valid_out_0_18 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5514) begin
      ic_tag_valid_out_0_19 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5530) begin
      ic_tag_valid_out_0_20 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5546) begin
      ic_tag_valid_out_0_21 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5562) begin
      ic_tag_valid_out_0_22 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5578) begin
      ic_tag_valid_out_0_23 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5594) begin
      ic_tag_valid_out_0_24 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5610) begin
      ic_tag_valid_out_0_25 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5626) begin
      ic_tag_valid_out_0_26 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5642) begin
      ic_tag_valid_out_0_27 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5658) begin
      ic_tag_valid_out_0_28 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5674) begin
      ic_tag_valid_out_0_29 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5690) begin
      ic_tag_valid_out_0_30 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5706) begin
      ic_tag_valid_out_0_31 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6234) begin
      ic_tag_valid_out_0_32 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6250) begin
      ic_tag_valid_out_0_33 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6266) begin
      ic_tag_valid_out_0_34 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6282) begin
      ic_tag_valid_out_0_35 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6298) begin
      ic_tag_valid_out_0_36 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6314) begin
      ic_tag_valid_out_0_37 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6330) begin
      ic_tag_valid_out_0_38 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6346) begin
      ic_tag_valid_out_0_39 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6362) begin
      ic_tag_valid_out_0_40 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6378) begin
      ic_tag_valid_out_0_41 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6394) begin
      ic_tag_valid_out_0_42 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6410) begin
      ic_tag_valid_out_0_43 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6426) begin
      ic_tag_valid_out_0_44 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6442) begin
      ic_tag_valid_out_0_45 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6458) begin
      ic_tag_valid_out_0_46 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6474) begin
      ic_tag_valid_out_0_47 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6490) begin
      ic_tag_valid_out_0_48 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6506) begin
      ic_tag_valid_out_0_49 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6522) begin
      ic_tag_valid_out_0_50 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6538) begin
      ic_tag_valid_out_0_51 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6554) begin
      ic_tag_valid_out_0_52 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6570) begin
      ic_tag_valid_out_0_53 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6586) begin
      ic_tag_valid_out_0_54 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6602) begin
      ic_tag_valid_out_0_55 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6618) begin
      ic_tag_valid_out_0_56 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6634) begin
      ic_tag_valid_out_0_57 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6650) begin
      ic_tag_valid_out_0_58 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6666) begin
      ic_tag_valid_out_0_59 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6682) begin
      ic_tag_valid_out_0_60 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6698) begin
      ic_tag_valid_out_0_61 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6714) begin
      ic_tag_valid_out_0_62 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6730) begin
      ic_tag_valid_out_0_63 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7258) begin
      ic_tag_valid_out_0_64 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7274) begin
      ic_tag_valid_out_0_65 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7290) begin
      ic_tag_valid_out_0_66 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7306) begin
      ic_tag_valid_out_0_67 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7322) begin
      ic_tag_valid_out_0_68 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7338) begin
      ic_tag_valid_out_0_69 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7354) begin
      ic_tag_valid_out_0_70 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7370) begin
      ic_tag_valid_out_0_71 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7386) begin
      ic_tag_valid_out_0_72 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7402) begin
      ic_tag_valid_out_0_73 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7418) begin
      ic_tag_valid_out_0_74 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7434) begin
      ic_tag_valid_out_0_75 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7450) begin
      ic_tag_valid_out_0_76 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7466) begin
      ic_tag_valid_out_0_77 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7482) begin
      ic_tag_valid_out_0_78 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7498) begin
      ic_tag_valid_out_0_79 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7514) begin
      ic_tag_valid_out_0_80 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7530) begin
      ic_tag_valid_out_0_81 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7546) begin
      ic_tag_valid_out_0_82 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7562) begin
      ic_tag_valid_out_0_83 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7578) begin
      ic_tag_valid_out_0_84 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7594) begin
      ic_tag_valid_out_0_85 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7610) begin
      ic_tag_valid_out_0_86 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7626) begin
      ic_tag_valid_out_0_87 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7642) begin
      ic_tag_valid_out_0_88 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7658) begin
      ic_tag_valid_out_0_89 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7674) begin
      ic_tag_valid_out_0_90 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7690) begin
      ic_tag_valid_out_0_91 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7706) begin
      ic_tag_valid_out_0_92 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7722) begin
      ic_tag_valid_out_0_93 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7738) begin
      ic_tag_valid_out_0_94 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7754) begin
      ic_tag_valid_out_0_95 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8282) begin
      ic_tag_valid_out_0_96 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8298) begin
      ic_tag_valid_out_0_97 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8314) begin
      ic_tag_valid_out_0_98 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8330) begin
      ic_tag_valid_out_0_99 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8346) begin
      ic_tag_valid_out_0_100 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8362) begin
      ic_tag_valid_out_0_101 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8378) begin
      ic_tag_valid_out_0_102 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8394) begin
      ic_tag_valid_out_0_103 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8410) begin
      ic_tag_valid_out_0_104 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8426) begin
      ic_tag_valid_out_0_105 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8442) begin
      ic_tag_valid_out_0_106 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8458) begin
      ic_tag_valid_out_0_107 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8474) begin
      ic_tag_valid_out_0_108 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8490) begin
      ic_tag_valid_out_0_109 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8506) begin
      ic_tag_valid_out_0_110 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8522) begin
      ic_tag_valid_out_0_111 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8538) begin
      ic_tag_valid_out_0_112 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8554) begin
      ic_tag_valid_out_0_113 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8570) begin
      ic_tag_valid_out_0_114 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8586) begin
      ic_tag_valid_out_0_115 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8602) begin
      ic_tag_valid_out_0_116 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8618) begin
      ic_tag_valid_out_0_117 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8634) begin
      ic_tag_valid_out_0_118 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8650) begin
      ic_tag_valid_out_0_119 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8666) begin
      ic_tag_valid_out_0_120 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8682) begin
      ic_tag_valid_out_0_121 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8698) begin
      ic_tag_valid_out_0_122 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8714) begin
      ic_tag_valid_out_0_123 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8730) begin
      ic_tag_valid_out_0_124 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8746) begin
      ic_tag_valid_out_0_125 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8762) begin
      ic_tag_valid_out_0_126 <= _T_5201;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8778) begin
      ic_tag_valid_out_0_127 <= _T_5201;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1211 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1211 <= {{5'd0}, _T_1210};
    end else begin
      _T_1211 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2512) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2587) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2631;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2413) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2415) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2425) begin
        perr_state <= 3'h0;
      end else if (_T_2428) begin
        if (_T_2430) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2434) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2438) begin
        err_stop_state <= 2'h1;
      end else if (_T_2443) begin
        if (_T_2445) begin
          err_stop_state <= 2'h0;
        end else if (_T_2466) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2470) begin
        if (_T_2445) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2487) begin
        if (_T_2491) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1356;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_5114 <= 7'h0;
    end else if (_T_3935) begin
      _T_5114 <= io_ic_debug_addr[9:3];
    end else begin
      _T_5114 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1396;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3870;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3045;
    end else begin
      iccm_dma_rdata <= _T_3046;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3866;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3935) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3938) begin
      way_status_new_ff <= _T_3942;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3938) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10131 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10131 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10101 <= 1'h0;
    end else begin
      _T_10101 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10102 <= 1'h0;
    end else begin
      _T_10102 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10103 <= 1'h0;
    end else begin
      _T_10103 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10107 <= 1'h0;
    end else begin
      _T_10107 <= _T_10106;
    end
    if (reset) begin
      _T_10108 <= 1'h0;
    end else begin
      _T_10108 <= bus_cmd_sent;
    end
  end
endmodule
