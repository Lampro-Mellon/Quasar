module el2_ifu_mem_ctl(
  input          clock,
  input          reset,
  input          io_free_clk,
  input          io_active_clk,
  input          io_exu_flush_final,
  input          io_dec_tlu_flush_lower_wb,
  input          io_dec_tlu_flush_err_wb,
  input          io_dec_tlu_i0_commit_cmt,
  input          io_dec_tlu_force_halt,
  input  [30:0]  io_ifc_fetch_addr_bf,
  input          io_ifc_fetch_uncacheable_bf,
  input          io_ifc_fetch_req_bf,
  input          io_ifc_fetch_req_bf_raw,
  input          io_ifc_iccm_access_bf,
  input          io_ifc_region_acc_fault_bf,
  input          io_ifc_dma_access_ok,
  input          io_dec_tlu_fence_i_wb,
  input          io_ifu_bp_hit_taken_f,
  input          io_ifu_bp_inst_mask_f,
  input          io_ifu_axi_arready,
  input          io_ifu_axi_rvalid,
  input  [2:0]   io_ifu_axi_rid,
  input  [63:0]  io_ifu_axi_rdata,
  input  [1:0]   io_ifu_axi_rresp,
  input          io_ifu_bus_clk_en,
  input          io_dma_iccm_req,
  input  [31:0]  io_dma_mem_addr,
  input  [2:0]   io_dma_mem_sz,
  input          io_dma_mem_write,
  input  [63:0]  io_dma_mem_wdata,
  input  [2:0]   io_dma_mem_tag,
  input  [63:0]  io_ic_rd_data,
  input  [70:0]  io_ic_debug_rd_data,
  input  [25:0]  io_ictag_debug_rd_data,
  input  [1:0]   io_ic_eccerr,
  input  [1:0]   io_ic_parerr,
  input  [1:0]   io_ic_rd_hit,
  input          io_ic_tag_perr,
  input  [63:0]  io_iccm_rd_data,
  input  [77:0]  io_iccm_rd_data_ecc,
  input  [1:0]   io_ifu_fetch_val,
  input  [70:0]  io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0]  io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input          io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input          io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output         io_ifu_miss_state_idle,
  output         io_ifu_ic_mb_empty,
  output         io_ic_dma_active,
  output         io_ic_write_stall,
  output         io_ifu_pmu_ic_miss,
  output         io_ifu_pmu_ic_hit,
  output         io_ifu_pmu_bus_error,
  output         io_ifu_pmu_bus_busy,
  output         io_ifu_pmu_bus_trxn,
  output         io_ifu_axi_awvalid,
  output [2:0]   io_ifu_axi_awid,
  output [31:0]  io_ifu_axi_awaddr,
  output [3:0]   io_ifu_axi_awregion,
  output [7:0]   io_ifu_axi_awlen,
  output [2:0]   io_ifu_axi_awsize,
  output [1:0]   io_ifu_axi_awburst,
  output         io_ifu_axi_awlock,
  output [3:0]   io_ifu_axi_awcache,
  output [2:0]   io_ifu_axi_awprot,
  output [3:0]   io_ifu_axi_awqos,
  output         io_ifu_axi_wvalid,
  output [63:0]  io_ifu_axi_wdata,
  output [7:0]   io_ifu_axi_wstrb,
  output         io_ifu_axi_wlast,
  output         io_ifu_axi_bready,
  output         io_ifu_axi_arvalid,
  output [2:0]   io_ifu_axi_arid,
  output [31:0]  io_ifu_axi_araddr,
  output [3:0]   io_ifu_axi_arregion,
  output [7:0]   io_ifu_axi_arlen,
  output [2:0]   io_ifu_axi_arsize,
  output [1:0]   io_ifu_axi_arburst,
  output         io_ifu_axi_arlock,
  output [3:0]   io_ifu_axi_arcache,
  output [2:0]   io_ifu_axi_arprot,
  output [3:0]   io_ifu_axi_arqos,
  output         io_ifu_axi_rready,
  output         io_iccm_dma_ecc_error,
  output         io_iccm_dma_rvalid,
  output [63:0]  io_iccm_dma_rdata,
  output [2:0]   io_iccm_dma_rtag,
  output         io_iccm_ready,
  output [30:0]  io_ic_rw_addr,
  output [1:0]   io_ic_wr_en,
  output         io_ic_rd_en,
  output [70:0]  io_ic_wr_data_0,
  output [70:0]  io_ic_wr_data_1,
  output [70:0]  io_ic_debug_wr_data,
  output [70:0]  io_ifu_ic_debug_rd_data,
  output [9:0]   io_ic_debug_addr,
  output         io_ic_debug_rd_en,
  output         io_ic_debug_wr_en,
  output         io_ic_debug_tag_array,
  output [1:0]   io_ic_debug_way,
  output [1:0]   io_ic_tag_valid,
  output [14:0]  io_iccm_rw_addr,
  output         io_iccm_wren,
  output         io_iccm_rden,
  output [77:0]  io_iccm_wr_data,
  output [2:0]   io_iccm_wr_size,
  output         io_ic_hit_f,
  output         io_ic_access_fault_f,
  output [1:0]   io_ic_access_fault_type_f,
  output         io_iccm_rd_ecc_single_err,
  output         io_iccm_rd_ecc_double_err,
  output         io_ic_error_start,
  output         io_ifu_async_error_start,
  output         io_iccm_dma_sb_error,
  output [1:0]   io_ic_fetch_val_f,
  output [31:0]  io_ic_data_f,
  output [63:0]  io_ic_premux_data,
  output         io_ic_sel_premux_data,
  input          io_dec_tlu_core_ecc_disable,
  output         io_ifu_ic_debug_rd_data_valid,
  output         io_iccm_buf_correct_ecc,
  output         io_iccm_correction_state,
  input          io_scan_mode,
  output [255:0] io_valids,
  output [1:0]   io_tagv_mb_in,
  output         io_test,
  output [127:0] io_test_way_status_out,
  output [15:0]  io_test_way_status_clken
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [63:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 189:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 324:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 325:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 325:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 257:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 551:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 553:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 191:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 312:34]
  wire [4:0] _GEN_464 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 668:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_464 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 668:53]
  wire [1:0] _GEN_465 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 671:91]
  wire [1:0] _T_3121 = ic_fetch_val_shift_right[3:2] & _GEN_465; // @[el2_ifu_mem_ctl.scala 671:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 326:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 279:46]
  wire [1:0] _GEN_466 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 671:113]
  wire [1:0] _T_3122 = _T_3121 & _GEN_466; // @[el2_ifu_mem_ctl.scala 671:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 657:59]
  wire [1:0] _GEN_467 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 671:130]
  wire [1:0] _T_3123 = _T_3122 | _GEN_467; // @[el2_ifu_mem_ctl.scala 671:130]
  wire  _T_3124 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 671:154]
  wire [1:0] _GEN_468 = {{1'd0}, _T_3124}; // @[el2_ifu_mem_ctl.scala 671:152]
  wire [1:0] _T_3125 = _T_3123 & _GEN_468; // @[el2_ifu_mem_ctl.scala 671:152]
  wire [1:0] _T_3114 = ic_fetch_val_shift_right[1:0] & _GEN_465; // @[el2_ifu_mem_ctl.scala 671:91]
  wire [1:0] _T_3115 = _T_3114 & _GEN_466; // @[el2_ifu_mem_ctl.scala 671:113]
  wire [1:0] _T_3116 = _T_3115 | _GEN_467; // @[el2_ifu_mem_ctl.scala 671:130]
  wire [1:0] _T_3118 = _T_3116 & _GEN_468; // @[el2_ifu_mem_ctl.scala 671:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3125,_T_3118}; // @[Cat.scala 29:58]
  wire  _T_3225 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3226 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3227 = _T_3225 ^ _T_3226; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3235 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3236 = ^_T_3235; // @[el2_lib.scala 301:83]
  wire  _T_3237 = io_iccm_rd_data_ecc[37] ^ _T_3236; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3244 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3252 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3244}; // @[el2_lib.scala 301:103]
  wire  _T_3253 = ^_T_3252; // @[el2_lib.scala 301:110]
  wire  _T_3254 = io_iccm_rd_data_ecc[36] ^ _T_3253; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3261 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3269 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3261}; // @[el2_lib.scala 301:130]
  wire  _T_3270 = ^_T_3269; // @[el2_lib.scala 301:137]
  wire  _T_3271 = io_iccm_rd_data_ecc[35] ^ _T_3270; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3280 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3289 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3280}; // @[el2_lib.scala 301:157]
  wire  _T_3290 = ^_T_3289; // @[el2_lib.scala 301:164]
  wire  _T_3291 = io_iccm_rd_data_ecc[34] ^ _T_3290; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3300 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3309 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3300}; // @[el2_lib.scala 301:184]
  wire  _T_3310 = ^_T_3309; // @[el2_lib.scala 301:191]
  wire  _T_3311 = io_iccm_rd_data_ecc[33] ^ _T_3310; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3320 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3329 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3320}; // @[el2_lib.scala 301:211]
  wire  _T_3330 = ^_T_3329; // @[el2_lib.scala 301:218]
  wire  _T_3331 = io_iccm_rd_data_ecc[32] ^ _T_3330; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3337 = {_T_3227,_T_3237,_T_3254,_T_3271,_T_3291,_T_3311,_T_3331}; // @[Cat.scala 29:58]
  wire  _T_3338 = _T_3337 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3339 = iccm_ecc_word_enable[0] & _T_3338; // @[el2_lib.scala 302:32]
  wire  _T_3341 = _T_3339 & _T_3337[6]; // @[el2_lib.scala 302:53]
  wire  _T_3610 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3611 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3612 = _T_3610 ^ _T_3611; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3620 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3621 = ^_T_3620; // @[el2_lib.scala 301:83]
  wire  _T_3622 = io_iccm_rd_data_ecc[76] ^ _T_3621; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3629 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3637 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3629}; // @[el2_lib.scala 301:103]
  wire  _T_3638 = ^_T_3637; // @[el2_lib.scala 301:110]
  wire  _T_3639 = io_iccm_rd_data_ecc[75] ^ _T_3638; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3646 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3654 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3646}; // @[el2_lib.scala 301:130]
  wire  _T_3655 = ^_T_3654; // @[el2_lib.scala 301:137]
  wire  _T_3656 = io_iccm_rd_data_ecc[74] ^ _T_3655; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3665 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3674 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3665}; // @[el2_lib.scala 301:157]
  wire  _T_3675 = ^_T_3674; // @[el2_lib.scala 301:164]
  wire  _T_3676 = io_iccm_rd_data_ecc[73] ^ _T_3675; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3685 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3694 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3685}; // @[el2_lib.scala 301:184]
  wire  _T_3695 = ^_T_3694; // @[el2_lib.scala 301:191]
  wire  _T_3696 = io_iccm_rd_data_ecc[72] ^ _T_3695; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3705 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3714 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3705}; // @[el2_lib.scala 301:211]
  wire  _T_3715 = ^_T_3714; // @[el2_lib.scala 301:218]
  wire  _T_3716 = io_iccm_rd_data_ecc[71] ^ _T_3715; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3722 = {_T_3612,_T_3622,_T_3639,_T_3656,_T_3676,_T_3696,_T_3716}; // @[Cat.scala 29:58]
  wire  _T_3723 = _T_3722 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3724 = iccm_ecc_word_enable[1] & _T_3723; // @[el2_lib.scala 302:32]
  wire  _T_3726 = _T_3724 & _T_3722[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3341,_T_3726}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 194:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 635:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 195:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 196:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 480:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 196:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 196:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 196:72]
  wire  _T_2490 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2495 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2515 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 530:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 394:42]
  wire  _T_2517 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 530:79]
  wire  _T_2518 = _T_2515 | _T_2517; // @[el2_ifu_mem_ctl.scala 530:56]
  wire  _T_2519 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 530:122]
  wire  _T_2520 = ~_T_2519; // @[el2_ifu_mem_ctl.scala 530:101]
  wire  _T_2521 = _T_2518 & _T_2520; // @[el2_ifu_mem_ctl.scala 530:99]
  wire  _T_2522 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2536 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 537:45]
  wire  _T_2537 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 537:69]
  wire  _T_2538 = _T_2536 & _T_2537; // @[el2_ifu_mem_ctl.scala 537:67]
  wire  _T_2539 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_2522 ? _T_2538 : _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2495 ? _T_2521 : _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2490 ? 1'h0 : _GEN_59; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 196:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 198:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 198:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 287:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 287:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 703:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 287:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 278:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 278:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 328:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 278:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 278:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 287:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 287:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 287:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 287:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 287:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 550:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 592:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 619:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 314:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 600:56]
  wire  _T_2641 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 617:69]
  wire  _T_2642 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 617:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2641 : _T_2642; // @[el2_ifu_mem_ctl.scala 617:28]
  wire  _T_2588 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 596:68]
  wire  _T_2589 = ic_act_miss_f | _T_2588; // @[el2_ifu_mem_ctl.scala 596:48]
  wire  bus_reset_data_beat_cnt = _T_2589 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 596:91]
  wire  _T_2585 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 595:50]
  wire  _T_2586 = bus_ifu_wr_en_ff & _T_2585; // @[el2_ifu_mem_ctl.scala 595:48]
  wire  _T_2587 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 595:72]
  wire  bus_inc_data_beat_cnt = _T_2586 & _T_2587; // @[el2_ifu_mem_ctl.scala 595:70]
  wire [2:0] _T_2593 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 599:115]
  wire [2:0] _T_2595 = bus_inc_data_beat_cnt ? _T_2593 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2590 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 597:32]
  wire  _T_2591 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 597:57]
  wire  bus_hold_data_beat_cnt = _T_2590 & _T_2591; // @[el2_ifu_mem_ctl.scala 597:55]
  wire [2:0] _T_2596 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2595 | _T_2596; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 198:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 198:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 199:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 198:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 199:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 205:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 430:45]
  wire  _T_2120 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 451:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 407:60]
  wire  _T_2151 = _T_2120 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2124 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2152 = _T_2124 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2159 = _T_2151 | _T_2152; // @[Mux.scala 27:72]
  wire  _T_2128 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2153 = _T_2128 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2160 = _T_2159 | _T_2153; // @[Mux.scala 27:72]
  wire  _T_2132 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2154 = _T_2132 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2161 = _T_2160 | _T_2154; // @[Mux.scala 27:72]
  wire  _T_2136 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2155 = _T_2136 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2162 = _T_2161 | _T_2155; // @[Mux.scala 27:72]
  wire  _T_2140 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2156 = _T_2140 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2163 = _T_2162 | _T_2156; // @[Mux.scala 27:72]
  wire  _T_2144 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2157 = _T_2144 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2164 = _T_2163 | _T_2157; // @[Mux.scala 27:72]
  wire  _T_2148 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 451:127]
  wire  _T_2158 = _T_2148 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2164 | _T_2158; // @[Mux.scala 27:72]
  wire  _T_2206 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 453:69]
  wire  _T_2207 = ic_miss_buff_data_valid_bypass_index & _T_2206; // @[el2_ifu_mem_ctl.scala 453:67]
  wire  _T_2209 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 453:91]
  wire  _T_2210 = _T_2207 & _T_2209; // @[el2_ifu_mem_ctl.scala 453:89]
  wire  _T_2215 = _T_2207 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 454:65]
  wire  _T_2216 = _T_2210 | _T_2215; // @[el2_ifu_mem_ctl.scala 453:112]
  wire  _T_2218 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 455:43]
  wire  _T_2221 = _T_2218 & _T_2209; // @[el2_ifu_mem_ctl.scala 455:65]
  wire  _T_2222 = _T_2216 | _T_2221; // @[el2_ifu_mem_ctl.scala 454:88]
  wire  _T_2226 = _T_2218 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 456:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 433:75]
  wire  _T_2166 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2190 = _T_2166 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2169 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2191 = _T_2169 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2190 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2172 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2192 = _T_2172 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2199 = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2193 = _T_2175 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2199 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2178 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2194 = _T_2178 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2181 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2195 = _T_2181 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2184 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2196 = _T_2184 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2187 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 452:110]
  wire  _T_2197 = _T_2187 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2227 = _T_2226 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 456:87]
  wire  _T_2228 = _T_2222 | _T_2227; // @[el2_ifu_mem_ctl.scala 455:88]
  wire  _T_2232 = ic_miss_buff_data_valid_bypass_index & _T_2148; // @[el2_ifu_mem_ctl.scala 457:43]
  wire  miss_buff_hit_unq_f = _T_2228 | _T_2232; // @[el2_ifu_mem_ctl.scala 456:131]
  wire  _T_2248 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 462:55]
  wire  _T_2249 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 462:87]
  wire  _T_2250 = _T_2248 | _T_2249; // @[el2_ifu_mem_ctl.scala 462:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2250; // @[el2_ifu_mem_ctl.scala 462:41]
  wire  _T_2233 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 459:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 315:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 450:51]
  wire  _T_2234 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 459:68]
  wire  _T_2235 = miss_buff_hit_unq_f & _T_2234; // @[el2_ifu_mem_ctl.scala 459:66]
  wire  stream_hit_f = _T_2233 & _T_2235; // @[el2_ifu_mem_ctl.scala 459:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 282:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 282:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 282:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 602:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 629:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 209:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 209:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 209:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 209:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 210:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 210:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 210:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 211:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 211:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 211:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 211:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 212:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 213:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 213:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 213:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 201:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 213:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 213:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 214:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 214:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 214:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 214:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 215:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 216:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 216:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 216:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 215:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 214:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 213:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 212:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 211:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 210:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 209:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2245 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 461:60]
  wire  _T_2246 = _T_2245 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 461:94]
  wire  stream_eol_f = _T_2246 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 461:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 224:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 224:87]
  wire  _T_113 = _T_111 & _T_2587; // @[el2_ifu_mem_ctl.scala 224:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 228:48]
  wire  _T_126 = _T_124 & _T_2587; // @[el2_ifu_mem_ctl.scala 228:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 288:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 288:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 288:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 288:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 288:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 289:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 288:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 289:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 342:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 289:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 289:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 289:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 232:50]
  wire  _T_137 = _T_135 & _T_2587; // @[el2_ifu_mem_ctl.scala 232:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 290:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 291:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 291:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 290:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 233:35]
  wire  _T_143 = _T_141 & _T_2587; // @[el2_ifu_mem_ctl.scala 233:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 233:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 232:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 238:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 237:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 237:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 242:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 242:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 199:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 199:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 199:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 199:91]
  wire  _T_30 = ic_act_miss_f & _T_2587; // @[el2_ifu_mem_ctl.scala 206:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 217:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 217:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 217:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 217:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 217:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 221:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 221:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 225:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 229:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 229:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 234:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 234:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 234:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 239:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 239:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 258:95]
  wire  _T_175 = _T_2248 & _T_174; // @[el2_ifu_mem_ctl.scala 258:93]
  wire  crit_wd_byp_ok_ff = _T_2249 | _T_175; // @[el2_ifu_mem_ctl.scala 258:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 259:36]
  wire  _T_180 = _T_2248 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 259:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 259:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 259:70]
  wire  _T_184 = _T_2248 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 260:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 259:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 260:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 261:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 261:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 260:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 263:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 263:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 271:35]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 737:14]
  wire  _T_5297 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5299 = _T_5297 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5300 = _T_5299 & _GEN_473; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5293 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5295 = _T_5293 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire [5:0] _GEN_474 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5296 = _T_5295 & _GEN_474; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5289 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5291 = _T_5289 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5292 = _T_5291 & _GEN_475; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5285 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5287 = _T_5285 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire [5:0] _GEN_476 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5288 = _T_5287 & _GEN_476; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5281 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5283 = _T_5281 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5284 = _T_5283 & _GEN_477; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5277 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5279 = _T_5277 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire [5:0] _GEN_478 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5280 = _T_5279 & _GEN_478; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5273 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5275 = _T_5273 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5276 = _T_5275 & _GEN_479; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5269 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5271 = _T_5269 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire [5:0] _GEN_480 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5272 = _T_5271 & _GEN_480; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5265 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5267 = _T_5265 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5268 = _T_5267 & _GEN_481; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5261 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5263 = _T_5261 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire [5:0] _GEN_482 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5264 = _T_5263 & _GEN_482; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [59:0] _T_5309 = {_T_5300,_T_5296,_T_5292,_T_5288,_T_5284,_T_5280,_T_5276,_T_5272,_T_5268,_T_5264}; // @[Cat.scala 29:58]
  wire  _T_5257 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5259 = _T_5257 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5260 = _T_5259 & _GEN_483; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5253 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5255 = _T_5253 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire [5:0] _GEN_484 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5256 = _T_5255 & _GEN_484; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5249 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5251 = _T_5249 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5252 = _T_5251 & _GEN_485; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5245 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5247 = _T_5245 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire [5:0] _GEN_486 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5248 = _T_5247 & _GEN_486; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5241 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5243 = _T_5241 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5244 = _T_5243 & _GEN_487; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5237 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5239 = _T_5237 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire [5:0] _GEN_488 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5240 = _T_5239 & _GEN_488; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5233 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5235 = _T_5233 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5236 = _T_5235 & _GEN_489; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5229 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5231 = _T_5229 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire [5:0] _GEN_490 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5232 = _T_5231 & _GEN_490; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5225 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5227 = _T_5225 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5228 = _T_5227 & _GEN_491; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [113:0] _T_5318 = {_T_5309,_T_5260,_T_5256,_T_5252,_T_5248,_T_5244,_T_5240,_T_5236,_T_5232,_T_5228}; // @[Cat.scala 29:58]
  wire  _T_5221 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5223 = _T_5221 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire [5:0] _GEN_492 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5224 = _T_5223 & _GEN_492; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5217 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5219 = _T_5217 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5220 = _T_5219 & _GEN_493; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5213 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5215 = _T_5213 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire [5:0] _GEN_494 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5216 = _T_5215 & _GEN_494; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5209 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5211 = _T_5209 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5212 = _T_5211 & _GEN_495; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5205 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5207 = _T_5205 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire [5:0] _GEN_496 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5208 = _T_5207 & _GEN_496; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5201 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5203 = _T_5201 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5204 = _T_5203 & _GEN_497; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5197 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5199 = _T_5197 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire [5:0] _GEN_498 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5200 = _T_5199 & _GEN_498; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5193 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5195 = _T_5193 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5196 = _T_5195 & _GEN_499; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5189 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5191 = _T_5189 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire [5:0] _GEN_500 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5192 = _T_5191 & _GEN_500; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [167:0] _T_5327 = {_T_5318,_T_5224,_T_5220,_T_5216,_T_5212,_T_5208,_T_5204,_T_5200,_T_5196,_T_5192}; // @[Cat.scala 29:58]
  wire  _T_5185 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5187 = _T_5185 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5188 = _T_5187 & _GEN_501; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5181 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5183 = _T_5181 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire [5:0] _GEN_502 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5184 = _T_5183 & _GEN_502; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5177 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5179 = _T_5177 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5180 = _T_5179 & _GEN_503; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5173 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5175 = _T_5173 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire [5:0] _GEN_504 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5176 = _T_5175 & _GEN_504; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5169 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5171 = _T_5169 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5172 = _T_5171 & _GEN_505; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5165 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5167 = _T_5165 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire [5:0] _GEN_506 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5168 = _T_5167 & _GEN_506; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5161 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5163 = _T_5161 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5164 = _T_5163 & _GEN_507; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5157 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5159 = _T_5157 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire [5:0] _GEN_508 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5160 = _T_5159 & _GEN_508; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5153 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5155 = _T_5153 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5156 = _T_5155 & _GEN_509; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [221:0] _T_5336 = {_T_5327,_T_5188,_T_5184,_T_5180,_T_5176,_T_5172,_T_5168,_T_5164,_T_5160,_T_5156}; // @[Cat.scala 29:58]
  wire  _T_5149 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5151 = _T_5149 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire [5:0] _GEN_510 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5152 = _T_5151 & _GEN_510; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5145 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5147 = _T_5145 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5148 = _T_5147 & _GEN_511; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5141 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5143 = _T_5141 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire [5:0] _GEN_512 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5144 = _T_5143 & _GEN_512; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5137 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5139 = _T_5137 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5140 = _T_5139 & _GEN_513; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5133 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5135 = _T_5133 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire [5:0] _GEN_514 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5136 = _T_5135 & _GEN_514; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5129 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5131 = _T_5129 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5132 = _T_5131 & _GEN_515; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5125 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5127 = _T_5125 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire [5:0] _GEN_516 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5128 = _T_5127 & _GEN_516; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5121 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5123 = _T_5121 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5124 = _T_5123 & _GEN_517; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5117 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5119 = _T_5117 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire [5:0] _GEN_518 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5120 = _T_5119 & _GEN_518; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [275:0] _T_5345 = {_T_5336,_T_5152,_T_5148,_T_5144,_T_5140,_T_5136,_T_5132,_T_5128,_T_5124,_T_5120}; // @[Cat.scala 29:58]
  wire  _T_5113 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5115 = _T_5113 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5116 = _T_5115 & _GEN_519; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5109 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5111 = _T_5109 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire [5:0] _GEN_520 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5112 = _T_5111 & _GEN_520; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5105 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5107 = _T_5105 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5108 = _T_5107 & _GEN_521; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5101 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5103 = _T_5101 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire [5:0] _GEN_522 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5104 = _T_5103 & _GEN_522; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5097 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5099 = _T_5097 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5100 = _T_5099 & _GEN_523; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5093 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5095 = _T_5093 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire [5:0] _GEN_524 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5096 = _T_5095 & _GEN_524; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5089 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5091 = _T_5089 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5092 = _T_5091 & _GEN_525; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5085 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5087 = _T_5085 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire [5:0] _GEN_526 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5088 = _T_5087 & _GEN_526; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5081 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5083 = _T_5081 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5084 = _T_5083 & _GEN_527; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [329:0] _T_5354 = {_T_5345,_T_5116,_T_5112,_T_5108,_T_5104,_T_5100,_T_5096,_T_5092,_T_5088,_T_5084}; // @[Cat.scala 29:58]
  wire  _T_5077 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5079 = _T_5077 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire [5:0] _GEN_528 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5080 = _T_5079 & _GEN_528; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5073 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5075 = _T_5073 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5076 = _T_5075 & _GEN_529; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5069 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5071 = _T_5069 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire [5:0] _GEN_530 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5072 = _T_5071 & _GEN_530; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5065 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5067 = _T_5065 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5068 = _T_5067 & _GEN_531; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5061 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5063 = _T_5061 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire [5:0] _GEN_532 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5064 = _T_5063 & _GEN_532; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5057 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5059 = _T_5057 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5060 = _T_5059 & _GEN_533; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5053 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5055 = _T_5053 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire [5:0] _GEN_534 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5056 = _T_5055 & _GEN_534; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5049 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5051 = _T_5049 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5052 = _T_5051 & _GEN_535; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5045 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5047 = _T_5045 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire [5:0] _GEN_536 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5048 = _T_5047 & _GEN_536; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [383:0] _T_5363 = {_T_5354,_T_5080,_T_5076,_T_5072,_T_5068,_T_5064,_T_5060,_T_5056,_T_5052,_T_5048}; // @[Cat.scala 29:58]
  wire  _T_5041 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5043 = _T_5041 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5044 = _T_5043 & _GEN_537; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5037 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5039 = _T_5037 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire [5:0] _GEN_538 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5040 = _T_5039 & _GEN_538; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5033 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5035 = _T_5033 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5036 = _T_5035 & _GEN_539; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5029 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5031 = _T_5029 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire [5:0] _GEN_540 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5032 = _T_5031 & _GEN_540; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5025 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5027 = _T_5025 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5028 = _T_5027 & _GEN_541; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5021 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5023 = _T_5021 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire [5:0] _GEN_542 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5024 = _T_5023 & _GEN_542; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5017 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5019 = _T_5017 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5020 = _T_5019 & _GEN_543; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5013 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5015 = _T_5013 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire [5:0] _GEN_544 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5016 = _T_5015 & _GEN_544; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5009 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5011 = _T_5009 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5012 = _T_5011 & _GEN_545; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [437:0] _T_5372 = {_T_5363,_T_5044,_T_5040,_T_5036,_T_5032,_T_5028,_T_5024,_T_5020,_T_5016,_T_5012}; // @[Cat.scala 29:58]
  wire  _T_5005 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5007 = _T_5005 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire [5:0] _GEN_546 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5008 = _T_5007 & _GEN_546; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_5001 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_5003 = _T_5001 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5004 = _T_5003 & _GEN_547; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4997 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4999 = _T_4997 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire [5:0] _GEN_548 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_5000 = _T_4999 & _GEN_548; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4993 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4995 = _T_4993 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4996 = _T_4995 & _GEN_549; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4989 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4991 = _T_4989 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire [5:0] _GEN_550 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4992 = _T_4991 & _GEN_550; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4985 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4987 = _T_4985 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4988 = _T_4987 & _GEN_551; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4981 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4983 = _T_4981 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire [5:0] _GEN_552 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4984 = _T_4983 & _GEN_552; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4977 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4979 = _T_4977 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4980 = _T_4979 & _GEN_553; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4973 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4975 = _T_4973 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire [5:0] _GEN_554 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4976 = _T_4975 & _GEN_554; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [491:0] _T_5381 = {_T_5372,_T_5008,_T_5004,_T_5000,_T_4996,_T_4992,_T_4988,_T_4984,_T_4980,_T_4976}; // @[Cat.scala 29:58]
  wire  _T_4969 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4971 = _T_4969 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4972 = _T_4971 & _GEN_555; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4965 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4967 = _T_4965 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire [5:0] _GEN_556 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4968 = _T_4967 & _GEN_556; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4961 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4963 = _T_4961 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4964 = _T_4963 & _GEN_557; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4957 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4959 = _T_4957 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire [5:0] _GEN_558 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4960 = _T_4959 & _GEN_558; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4953 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4955 = _T_4953 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4956 = _T_4955 & _GEN_559; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4949 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4951 = _T_4949 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire [5:0] _GEN_560 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4952 = _T_4951 & _GEN_560; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4945 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4947 = _T_4945 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4948 = _T_4947 & _GEN_561; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4941 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4943 = _T_4941 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire [5:0] _GEN_562 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4944 = _T_4943 & _GEN_562; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4937 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4939 = _T_4937 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4940 = _T_4939 & _GEN_563; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [545:0] _T_5390 = {_T_5381,_T_4972,_T_4968,_T_4964,_T_4960,_T_4956,_T_4952,_T_4948,_T_4944,_T_4940}; // @[Cat.scala 29:58]
  wire  _T_4933 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4935 = _T_4933 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire [5:0] _GEN_564 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4936 = _T_4935 & _GEN_564; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4929 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4931 = _T_4929 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4932 = _T_4931 & _GEN_565; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4925 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4927 = _T_4925 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire [5:0] _GEN_566 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4928 = _T_4927 & _GEN_566; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4921 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4923 = _T_4921 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4924 = _T_4923 & _GEN_567; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4917 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4919 = _T_4917 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire [5:0] _GEN_568 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4920 = _T_4919 & _GEN_568; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4913 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4915 = _T_4913 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4916 = _T_4915 & _GEN_569; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4909 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4911 = _T_4909 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire [5:0] _GEN_570 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4912 = _T_4911 & _GEN_570; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4905 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4907 = _T_4905 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4908 = _T_4907 & _GEN_571; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4901 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4903 = _T_4901 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire [5:0] _GEN_572 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4904 = _T_4903 & _GEN_572; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [599:0] _T_5399 = {_T_5390,_T_4936,_T_4932,_T_4928,_T_4924,_T_4920,_T_4916,_T_4912,_T_4908,_T_4904}; // @[Cat.scala 29:58]
  wire  _T_4897 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4899 = _T_4897 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4900 = _T_4899 & _GEN_573; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4893 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4895 = _T_4893 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire [5:0] _GEN_574 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4896 = _T_4895 & _GEN_574; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4889 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4891 = _T_4889 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4892 = _T_4891 & _GEN_575; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4885 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4887 = _T_4885 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire [5:0] _GEN_576 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4888 = _T_4887 & _GEN_576; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4881 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4883 = _T_4881 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4884 = _T_4883 & _GEN_577; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4877 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4879 = _T_4877 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire [5:0] _GEN_578 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4880 = _T_4879 & _GEN_578; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4873 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4875 = _T_4873 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4876 = _T_4875 & _GEN_579; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4869 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4871 = _T_4869 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire [5:0] _GEN_580 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4872 = _T_4871 & _GEN_580; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4865 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4867 = _T_4865 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4868 = _T_4867 & _GEN_581; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [653:0] _T_5408 = {_T_5399,_T_4900,_T_4896,_T_4892,_T_4888,_T_4884,_T_4880,_T_4876,_T_4872,_T_4868}; // @[Cat.scala 29:58]
  wire  _T_4861 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4863 = _T_4861 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire [5:0] _GEN_582 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4864 = _T_4863 & _GEN_582; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4857 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4859 = _T_4857 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4860 = _T_4859 & _GEN_583; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4853 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4855 = _T_4853 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire [5:0] _GEN_584 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4856 = _T_4855 & _GEN_584; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4849 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4851 = _T_4849 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4852 = _T_4851 & _GEN_585; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4845 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4847 = _T_4845 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire [5:0] _GEN_586 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4848 = _T_4847 & _GEN_586; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4841 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4843 = _T_4841 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4844 = _T_4843 & _GEN_587; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4837 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4839 = _T_4837 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire [5:0] _GEN_588 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4840 = _T_4839 & _GEN_588; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4833 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4835 = _T_4833 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4836 = _T_4835 & _GEN_589; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4829 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4831 = _T_4829 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire [5:0] _GEN_590 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4832 = _T_4831 & _GEN_590; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [707:0] _T_5417 = {_T_5408,_T_4864,_T_4860,_T_4856,_T_4852,_T_4848,_T_4844,_T_4840,_T_4836,_T_4832}; // @[Cat.scala 29:58]
  wire  _T_4825 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4827 = _T_4825 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4828 = _T_4827 & _GEN_591; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4821 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4823 = _T_4821 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire [5:0] _GEN_592 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4824 = _T_4823 & _GEN_592; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4817 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4819 = _T_4817 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4820 = _T_4819 & _GEN_593; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4813 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4815 = _T_4813 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire [5:0] _GEN_594 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4816 = _T_4815 & _GEN_594; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4809 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4811 = _T_4809 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4812 = _T_4811 & _GEN_595; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4805 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4807 = _T_4805 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire [5:0] _GEN_596 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4808 = _T_4807 & _GEN_596; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4801 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4803 = _T_4801 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4804 = _T_4803 & _GEN_597; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4797 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4799 = _T_4797 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire [5:0] _GEN_598 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4800 = _T_4799 & _GEN_598; // @[el2_ifu_mem_ctl.scala 733:128]
  wire  _T_4793 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4795 = _T_4793 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4796 = _T_4795 & _GEN_599; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [761:0] _T_5426 = {_T_5417,_T_4828,_T_4824,_T_4820,_T_4816,_T_4812,_T_4808,_T_4804,_T_4800,_T_4796}; // @[Cat.scala 29:58]
  wire  _T_4789 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 733:119]
  wire [5:0] _T_4791 = _T_4789 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [5:0] _T_4792 = _T_4791 & _GEN_600; // @[el2_ifu_mem_ctl.scala 733:128]
  wire [767:0] _T_5427 = {_T_5426,_T_4792}; // @[Cat.scala 29:58]
  wire  way_status = _T_5427[0]; // @[el2_ifu_mem_ctl.scala 733:14]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 266:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 266:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 272:29]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 270:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 275:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 280:59]
  wire  _T_214 = _T_212 | _T_2233; // @[el2_ifu_mem_ctl.scala 280:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 280:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 286:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 286:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 286:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 293:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 293:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 293:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 294:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 294:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 297:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 297:135]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2662 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 625:48]
  wire  _T_2663 = _T_2662 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 625:52]
  wire  bus_ifu_wr_data_error_ff = _T_2663 & miss_pending; // @[el2_ifu_mem_ctl.scala 625:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 370:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 369:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 297:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 297:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 300:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 300:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 301:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 320:30]
  wire  _T_10888 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 789:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 321:24]
  wire  _T_10890 = _T_10888 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 789:51]
  wire  _T_10892 = _T_10890 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 789:67]
  wire  _T_10894 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 789:86]
  wire  replace_way_mb_any_0 = _T_10892 | _T_10894; // @[el2_ifu_mem_ctl.scala 789:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10897 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:50]
  wire  _T_10899 = _T_10897 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 790:66]
  wire  _T_10901 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 790:85]
  wire  _T_10903 = _T_10901 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:100]
  wire  replace_way_mb_any_1 = _T_10899 | _T_10903; // @[el2_ifu_mem_ctl.scala 790:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 305:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 305:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 306:56]
  wire [1:0] _T_296 = miss_pending ? tagv_mb_ff : _T_295; // @[el2_ifu_mem_ctl.scala 306:6]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 309:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 309:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 310:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 309:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 309:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 311:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 319:23]
  wire  _T_313 = _T_2248 & flush_final_f; // @[el2_ifu_mem_ctl.scala 323:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 323:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 323:53]
  wire  _T_2240 = ~_T_2235; // @[el2_ifu_mem_ctl.scala 460:46]
  wire  _T_2241 = _T_2233 & _T_2240; // @[el2_ifu_mem_ctl.scala 460:44]
  wire  stream_miss_f = _T_2241 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 460:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 323:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 323:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 329:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_2233; // @[el2_ifu_mem_ctl.scala 331:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 331:82]
  wire  _T_2254 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 465:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2254}; // @[Cat.scala 29:58]
  wire  _T_2255 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2279 = _T_2255 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2258 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2280 = _T_2258 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2287 = _T_2279 | _T_2280; // @[Mux.scala 27:72]
  wire  _T_2261 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2281 = _T_2261 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2287 | _T_2281; // @[Mux.scala 27:72]
  wire  _T_2264 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2282 = _T_2264 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2288 | _T_2282; // @[Mux.scala 27:72]
  wire  _T_2267 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2283 = _T_2267 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2289 | _T_2283; // @[Mux.scala 27:72]
  wire  _T_2270 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2284 = _T_2270 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2290 | _T_2284; // @[Mux.scala 27:72]
  wire  _T_2273 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2285 = _T_2273 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2291 | _T_2285; // @[Mux.scala 27:72]
  wire  _T_2276 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 466:81]
  wire  _T_2286 = _T_2276 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2292 | _T_2286; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 467:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 335:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 335:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 622:61]
  wire  _T_2656 = ic_act_miss_f_delayed & _T_2249; // @[el2_ifu_mem_ctl.scala 623:53]
  wire  reset_tag_valid_for_miss = _T_2656 & _T_17; // @[el2_ifu_mem_ctl.scala 623:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 335:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 337:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 339:84]
  wire  _T_2650 = ~_T_2662; // @[el2_ifu_mem_ctl.scala 620:84]
  wire  _T_2651 = _T_100 & _T_2650; // @[el2_ifu_mem_ctl.scala 620:82]
  wire  bus_ifu_wr_en_ff_q = _T_2651 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 620:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 339:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 340:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_567 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 384:13]
  wire  _T_568 = ^_T_567; // @[el2_lib.scala 384:20]
  wire [6:0] _T_574 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_581 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 384:30]
  wire [14:0] _T_582 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_574}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_589 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 384:30]
  wire [30:0] _T_598 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_582}; // @[el2_lib.scala 384:30]
  wire  _T_599 = ^_T_598; // @[el2_lib.scala 384:37]
  wire [6:0] _T_605 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 384:47]
  wire [14:0] _T_613 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_605}; // @[el2_lib.scala 384:47]
  wire [30:0] _T_629 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_613}; // @[el2_lib.scala 384:47]
  wire  _T_630 = ^_T_629; // @[el2_lib.scala 384:54]
  wire [6:0] _T_636 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 384:64]
  wire [14:0] _T_644 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_636}; // @[el2_lib.scala 384:64]
  wire [30:0] _T_660 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_581,_T_644}; // @[el2_lib.scala 384:64]
  wire  _T_661 = ^_T_660; // @[el2_lib.scala 384:71]
  wire [7:0] _T_668 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 384:81]
  wire [16:0] _T_677 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_668}; // @[el2_lib.scala 384:81]
  wire [8:0] _T_685 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 384:81]
  wire [17:0] _T_694 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_685}; // @[el2_lib.scala 384:81]
  wire [34:0] _T_695 = {_T_694,_T_677}; // @[el2_lib.scala 384:81]
  wire  _T_696 = ^_T_695; // @[el2_lib.scala 384:88]
  wire [7:0] _T_703 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 384:98]
  wire [16:0] _T_712 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_703}; // @[el2_lib.scala 384:98]
  wire [8:0] _T_720 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 384:98]
  wire [17:0] _T_729 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_720}; // @[el2_lib.scala 384:98]
  wire [34:0] _T_730 = {_T_729,_T_712}; // @[el2_lib.scala 384:98]
  wire  _T_731 = ^_T_730; // @[el2_lib.scala 384:105]
  wire [7:0] _T_738 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 384:115]
  wire [16:0] _T_747 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_738}; // @[el2_lib.scala 384:115]
  wire [8:0] _T_755 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 384:115]
  wire [17:0] _T_764 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_755}; // @[el2_lib.scala 384:115]
  wire [34:0] _T_765 = {_T_764,_T_747}; // @[el2_lib.scala 384:115]
  wire  _T_766 = ^_T_765; // @[el2_lib.scala 384:122]
  wire [3:0] _T_2295 = {ifu_bus_rid_ff[2:1],_T_2254,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2296 = _T_2295 == 4'h0; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2343 = _T_2296 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2299 = _T_2295 == 4'h1; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2344 = _T_2299 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2343 | _T_2344; // @[Mux.scala 27:72]
  wire  _T_2302 = _T_2295 == 4'h2; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2345 = _T_2302 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2360 = _T_2359 | _T_2345; // @[Mux.scala 27:72]
  wire  _T_2305 = _T_2295 == 4'h3; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2346 = _T_2305 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2360 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2308 = _T_2295 == 4'h4; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2347 = _T_2308 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire  _T_2311 = _T_2295 == 4'h5; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2348 = _T_2311 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2363 = _T_2362 | _T_2348; // @[Mux.scala 27:72]
  wire  _T_2314 = _T_2295 == 4'h6; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2349 = _T_2314 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2364 = _T_2363 | _T_2349; // @[Mux.scala 27:72]
  wire  _T_2317 = _T_2295 == 4'h7; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2350 = _T_2317 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2365 = _T_2364 | _T_2350; // @[Mux.scala 27:72]
  wire  _T_2320 = _T_2295 == 4'h8; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2351 = _T_2320 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2366 = _T_2365 | _T_2351; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2295 == 4'h9; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2352 = _T_2323 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2367 = _T_2366 | _T_2352; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2295 == 4'ha; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2353 = _T_2326 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2368 = _T_2367 | _T_2353; // @[Mux.scala 27:72]
  wire  _T_2329 = _T_2295 == 4'hb; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2354 = _T_2329 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2369 = _T_2368 | _T_2354; // @[Mux.scala 27:72]
  wire  _T_2332 = _T_2295 == 4'hc; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2355 = _T_2332 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 27:72]
  wire  _T_2335 = _T_2295 == 4'hd; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2356 = _T_2335 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2371 = _T_2370 | _T_2356; // @[Mux.scala 27:72]
  wire  _T_2338 = _T_2295 == 4'he; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2357 = _T_2338 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2372 = _T_2371 | _T_2357; // @[Mux.scala 27:72]
  wire  _T_2341 = _T_2295 == 4'hf; // @[el2_ifu_mem_ctl.scala 468:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2358 = _T_2341 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2373 = _T_2372 | _T_2358; // @[Mux.scala 27:72]
  wire [3:0] _T_2375 = {ifu_bus_rid_ff[2:1],_T_2254,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2376 = _T_2375 == 4'h0; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2423 = _T_2376 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2375 == 4'h1; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2424 = _T_2379 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2439 = _T_2423 | _T_2424; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2375 == 4'h2; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2425 = _T_2382 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2440 = _T_2439 | _T_2425; // @[Mux.scala 27:72]
  wire  _T_2385 = _T_2375 == 4'h3; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2426 = _T_2385 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2441 = _T_2440 | _T_2426; // @[Mux.scala 27:72]
  wire  _T_2388 = _T_2375 == 4'h4; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2427 = _T_2388 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2442 = _T_2441 | _T_2427; // @[Mux.scala 27:72]
  wire  _T_2391 = _T_2375 == 4'h5; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2428 = _T_2391 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2443 = _T_2442 | _T_2428; // @[Mux.scala 27:72]
  wire  _T_2394 = _T_2375 == 4'h6; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2429 = _T_2394 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2444 = _T_2443 | _T_2429; // @[Mux.scala 27:72]
  wire  _T_2397 = _T_2375 == 4'h7; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2430 = _T_2397 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2445 = _T_2444 | _T_2430; // @[Mux.scala 27:72]
  wire  _T_2400 = _T_2375 == 4'h8; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2431 = _T_2400 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2446 = _T_2445 | _T_2431; // @[Mux.scala 27:72]
  wire  _T_2403 = _T_2375 == 4'h9; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2432 = _T_2403 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2447 = _T_2446 | _T_2432; // @[Mux.scala 27:72]
  wire  _T_2406 = _T_2375 == 4'ha; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2433 = _T_2406 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2448 = _T_2447 | _T_2433; // @[Mux.scala 27:72]
  wire  _T_2409 = _T_2375 == 4'hb; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2434 = _T_2409 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2449 = _T_2448 | _T_2434; // @[Mux.scala 27:72]
  wire  _T_2412 = _T_2375 == 4'hc; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2435 = _T_2412 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2450 = _T_2449 | _T_2435; // @[Mux.scala 27:72]
  wire  _T_2415 = _T_2375 == 4'hd; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2436 = _T_2415 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2451 = _T_2450 | _T_2436; // @[Mux.scala 27:72]
  wire  _T_2418 = _T_2375 == 4'he; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2437 = _T_2418 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2452 = _T_2451 | _T_2437; // @[Mux.scala 27:72]
  wire  _T_2421 = _T_2375 == 4'hf; // @[el2_ifu_mem_ctl.scala 469:66]
  wire [31:0] _T_2438 = _T_2421 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2453 = _T_2452 | _T_2438; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [6:0] _T_989 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 384:13]
  wire  _T_990 = ^_T_989; // @[el2_lib.scala 384:20]
  wire [6:0] _T_996 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_1003 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 384:30]
  wire [14:0] _T_1004 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_996}; // @[el2_lib.scala 384:30]
  wire [7:0] _T_1011 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 384:30]
  wire [30:0] _T_1020 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1004}; // @[el2_lib.scala 384:30]
  wire  _T_1021 = ^_T_1020; // @[el2_lib.scala 384:37]
  wire [6:0] _T_1027 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 384:47]
  wire [14:0] _T_1035 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1027}; // @[el2_lib.scala 384:47]
  wire [30:0] _T_1051 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1035}; // @[el2_lib.scala 384:47]
  wire  _T_1052 = ^_T_1051; // @[el2_lib.scala 384:54]
  wire [6:0] _T_1058 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 384:64]
  wire [14:0] _T_1066 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1058}; // @[el2_lib.scala 384:64]
  wire [30:0] _T_1082 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1003,_T_1066}; // @[el2_lib.scala 384:64]
  wire  _T_1083 = ^_T_1082; // @[el2_lib.scala 384:71]
  wire [7:0] _T_1090 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 384:81]
  wire [16:0] _T_1099 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1090}; // @[el2_lib.scala 384:81]
  wire [8:0] _T_1107 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 384:81]
  wire [17:0] _T_1116 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1107}; // @[el2_lib.scala 384:81]
  wire [34:0] _T_1117 = {_T_1116,_T_1099}; // @[el2_lib.scala 384:81]
  wire  _T_1118 = ^_T_1117; // @[el2_lib.scala 384:88]
  wire [7:0] _T_1125 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 384:98]
  wire [16:0] _T_1134 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1125}; // @[el2_lib.scala 384:98]
  wire [8:0] _T_1142 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 384:98]
  wire [17:0] _T_1151 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1142}; // @[el2_lib.scala 384:98]
  wire [34:0] _T_1152 = {_T_1151,_T_1134}; // @[el2_lib.scala 384:98]
  wire  _T_1153 = ^_T_1152; // @[el2_lib.scala 384:105]
  wire [7:0] _T_1160 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 384:115]
  wire [16:0] _T_1169 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1160}; // @[el2_lib.scala 384:115]
  wire [8:0] _T_1177 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 384:115]
  wire [17:0] _T_1186 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1177}; // @[el2_lib.scala 384:115]
  wire [34:0] _T_1187 = {_T_1186,_T_1169}; // @[el2_lib.scala 384:115]
  wire  _T_1188 = ^_T_1187; // @[el2_lib.scala 384:122]
  wire [70:0] _T_1233 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1232 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [141:0] _T_1234 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff,_T_1232}; // @[Cat.scala 29:58]
  wire [141:0] _T_1237 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453,_T_1233}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1234 : _T_1237; // @[el2_ifu_mem_ctl.scala 361:28]
  wire  _T_1196 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 351:56]
  wire  _T_1197 = _T_1196 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 351:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 415:28]
  wire  _T_1413 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 618:35]
  wire  _T_1282 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1339 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 406:118]
  wire  _T_1340 = ic_miss_buff_data_valid[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1340; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1436 = _T_1413 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1343 = ic_miss_buff_data_valid[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1343; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1437 = _T_1416 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1444 = _T_1436 | _T_1437; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1284 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1346 = ic_miss_buff_data_valid[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1346; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1438 = _T_1419 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1444 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1349 = ic_miss_buff_data_valid[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1349; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1439 = _T_1422 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1425 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1352 = ic_miss_buff_data_valid[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1352; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1440 = _T_1425 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1428 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1355 = ic_miss_buff_data_valid[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1355; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1441 = _T_1428 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1431 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1358 = ic_miss_buff_data_valid[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1358; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1442 = _T_1431 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1434 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 417:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 400:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 400:73]
  wire  _T_1361 = ic_miss_buff_data_valid[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 406:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1361; // @[el2_ifu_mem_ctl.scala 406:88]
  wire  _T_1443 = _T_1434 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1452 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 418:58]
  wire  _T_1453 = bypass_valid_value_check & _T_1452; // @[el2_ifu_mem_ctl.scala 418:56]
  wire  _T_1455 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 418:77]
  wire  _T_1456 = _T_1453 & _T_1455; // @[el2_ifu_mem_ctl.scala 418:75]
  wire  _T_1461 = _T_1453 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 419:75]
  wire  _T_1462 = _T_1456 | _T_1461; // @[el2_ifu_mem_ctl.scala 418:95]
  wire  _T_1464 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 420:56]
  wire  _T_1467 = _T_1464 & _T_1455; // @[el2_ifu_mem_ctl.scala 420:74]
  wire  _T_1468 = _T_1462 | _T_1467; // @[el2_ifu_mem_ctl.scala 419:94]
  wire  _T_1472 = _T_1464 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 421:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 416:70]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1489 = _T_1473 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1490 = _T_1475 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1497 = _T_1489 | _T_1490; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1491 = _T_1477 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1498 = _T_1497 | _T_1491; // @[Mux.scala 27:72]
  wire  _T_1479 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1492 = _T_1479 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1498 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1481 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1493 = _T_1481 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1499 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1483 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1494 = _T_1483 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1500 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1485 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1495 = _T_1485 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1501 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1487 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 421:132]
  wire  _T_1496 = _T_1487 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1502 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1472 & _T_1503; // @[el2_ifu_mem_ctl.scala 421:69]
  wire  _T_1506 = _T_1468 | _T_1505; // @[el2_ifu_mem_ctl.scala 420:94]
  wire [4:0] _GEN_601 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 422:95]
  wire  _T_1509 = _GEN_601 == 5'h1f; // @[el2_ifu_mem_ctl.scala 422:95]
  wire  _T_1510 = bypass_valid_value_check & _T_1509; // @[el2_ifu_mem_ctl.scala 422:56]
  wire  bypass_data_ready_in = _T_1506 | _T_1510; // @[el2_ifu_mem_ctl.scala 421:181]
  wire  _T_1511 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 426:53]
  wire  _T_1512 = _T_1511 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 426:73]
  wire  _T_1514 = _T_1512 & _T_317; // @[el2_ifu_mem_ctl.scala 426:96]
  wire  _T_1516 = _T_1514 & _T_58; // @[el2_ifu_mem_ctl.scala 426:118]
  wire  _T_1518 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 427:73]
  wire  _T_1520 = _T_1518 & _T_317; // @[el2_ifu_mem_ctl.scala 427:96]
  wire  _T_1522 = _T_1520 & _T_58; // @[el2_ifu_mem_ctl.scala 427:118]
  wire  _T_1523 = _T_1516 | _T_1522; // @[el2_ifu_mem_ctl.scala 426:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 429:58]
  wire  _T_1524 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 428:54]
  wire  _T_1525 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 428:76]
  wire  _T_1526 = _T_1524 & _T_1525; // @[el2_ifu_mem_ctl.scala 428:74]
  wire  _T_1528 = _T_1526 & _T_317; // @[el2_ifu_mem_ctl.scala 428:96]
  wire  ic_crit_wd_rdy_new_in = _T_1523 | _T_1528; // @[el2_ifu_mem_ctl.scala 427:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 628:43]
  wire  _T_1249 = ic_crit_wd_rdy | _T_2233; // @[el2_ifu_mem_ctl.scala 374:38]
  wire  _T_1251 = _T_1249 | _T_2249; // @[el2_ifu_mem_ctl.scala 374:64]
  wire  _T_1252 = ~_T_1251; // @[el2_ifu_mem_ctl.scala 374:21]
  wire  _T_1253 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 374:98]
  wire  sel_ic_data = _T_1252 & _T_1253; // @[el2_ifu_mem_ctl.scala 374:96]
  wire  _T_2456 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 473:44]
  wire  _T_1622 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 440:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 412:60]
  wire  _T_1566 = _T_1413 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1416 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1566 | _T_1567; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1419 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1574 | _T_1568; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1422 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1575 | _T_1569; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1425 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1570; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1428 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1571; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1431 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1572; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1434 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1579 | _T_1573; // @[Mux.scala 27:72]
  wire  _T_1605 = _T_2166 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1606 = _T_2169 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1613 = _T_1605 | _T_1606; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_2172 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1614 = _T_1613 | _T_1607; // @[Mux.scala 27:72]
  wire  _T_1608 = _T_2175 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1615 = _T_1614 | _T_1608; // @[Mux.scala 27:72]
  wire  _T_1609 = _T_2178 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1616 = _T_1615 | _T_1609; // @[Mux.scala 27:72]
  wire  _T_1610 = _T_2181 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1617 = _T_1616 | _T_1610; // @[Mux.scala 27:72]
  wire  _T_1611 = _T_2184 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1618 = _T_1617 | _T_1611; // @[Mux.scala 27:72]
  wire  _T_1612 = _T_2187 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1618 | _T_1612; // @[Mux.scala 27:72]
  wire  _T_1623 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 442:70]
  wire  ifu_byp_data_err_new = _T_1622 ? ic_miss_buff_data_error_bypass : _T_1623; // @[el2_ifu_mem_ctl.scala 440:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 385:42]
  wire  _T_2457 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 473:91]
  wire  _T_2458 = ~_T_2457; // @[el2_ifu_mem_ctl.scala 473:60]
  wire  ic_rd_parity_final_err = _T_2456 & _T_2458; // @[el2_ifu_mem_ctl.scala 473:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_10506 = _T_4789 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 764:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_10508 = _T_4793 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10761 = _T_10506 | _T_10508; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_10510 = _T_4797 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10762 = _T_10761 | _T_10510; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_10512 = _T_4801 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10763 = _T_10762 | _T_10512; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_10514 = _T_4805 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10764 = _T_10763 | _T_10514; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_10516 = _T_4809 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10765 = _T_10764 | _T_10516; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_10518 = _T_4813 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10766 = _T_10765 | _T_10518; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_10520 = _T_4817 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10767 = _T_10766 | _T_10520; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_10522 = _T_4821 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10768 = _T_10767 | _T_10522; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_10524 = _T_4825 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10769 = _T_10768 | _T_10524; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_10526 = _T_4829 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10770 = _T_10769 | _T_10526; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_10528 = _T_4833 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10771 = _T_10770 | _T_10528; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_10530 = _T_4837 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10772 = _T_10771 | _T_10530; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_10532 = _T_4841 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10773 = _T_10772 | _T_10532; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_10534 = _T_4845 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10774 = _T_10773 | _T_10534; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_10536 = _T_4849 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10775 = _T_10774 | _T_10536; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_10538 = _T_4853 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10776 = _T_10775 | _T_10538; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_10540 = _T_4857 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10777 = _T_10776 | _T_10540; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_10542 = _T_4861 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10778 = _T_10777 | _T_10542; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_10544 = _T_4865 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10779 = _T_10778 | _T_10544; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_10546 = _T_4869 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10780 = _T_10779 | _T_10546; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_10548 = _T_4873 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10781 = _T_10780 | _T_10548; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_10550 = _T_4877 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10782 = _T_10781 | _T_10550; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_10552 = _T_4881 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10783 = _T_10782 | _T_10552; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_10554 = _T_4885 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10784 = _T_10783 | _T_10554; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_10556 = _T_4889 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10785 = _T_10784 | _T_10556; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_10558 = _T_4893 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10786 = _T_10785 | _T_10558; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_10560 = _T_4897 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10787 = _T_10786 | _T_10560; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_10562 = _T_4901 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10788 = _T_10787 | _T_10562; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_10564 = _T_4905 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10789 = _T_10788 | _T_10564; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_10566 = _T_4909 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10790 = _T_10789 | _T_10566; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_10568 = _T_4913 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10791 = _T_10790 | _T_10568; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_10570 = _T_4917 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10792 = _T_10791 | _T_10570; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_10572 = _T_4921 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10793 = _T_10792 | _T_10572; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_10574 = _T_4925 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10794 = _T_10793 | _T_10574; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_10576 = _T_4929 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10795 = _T_10794 | _T_10576; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_10578 = _T_4933 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10796 = _T_10795 | _T_10578; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_10580 = _T_4937 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10797 = _T_10796 | _T_10580; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_10582 = _T_4941 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10798 = _T_10797 | _T_10582; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_10584 = _T_4945 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10799 = _T_10798 | _T_10584; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_10586 = _T_4949 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10800 = _T_10799 | _T_10586; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_10588 = _T_4953 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10801 = _T_10800 | _T_10588; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_10590 = _T_4957 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10802 = _T_10801 | _T_10590; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_10592 = _T_4961 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10803 = _T_10802 | _T_10592; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_10594 = _T_4965 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10804 = _T_10803 | _T_10594; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_10596 = _T_4969 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10805 = _T_10804 | _T_10596; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_10598 = _T_4973 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10806 = _T_10805 | _T_10598; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_10600 = _T_4977 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10807 = _T_10806 | _T_10600; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_10602 = _T_4981 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10808 = _T_10807 | _T_10602; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_10604 = _T_4985 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10809 = _T_10808 | _T_10604; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_10606 = _T_4989 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10810 = _T_10809 | _T_10606; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_10608 = _T_4993 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10811 = _T_10810 | _T_10608; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_10610 = _T_4997 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10812 = _T_10811 | _T_10610; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_10612 = _T_5001 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10813 = _T_10812 | _T_10612; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_10614 = _T_5005 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10814 = _T_10813 | _T_10614; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_10616 = _T_5009 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10815 = _T_10814 | _T_10616; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_10618 = _T_5013 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10816 = _T_10815 | _T_10618; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_10620 = _T_5017 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10817 = _T_10816 | _T_10620; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_10622 = _T_5021 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10818 = _T_10817 | _T_10622; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_10624 = _T_5025 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10819 = _T_10818 | _T_10624; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_10626 = _T_5029 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10820 = _T_10819 | _T_10626; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_10628 = _T_5033 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10821 = _T_10820 | _T_10628; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_10630 = _T_5037 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10822 = _T_10821 | _T_10630; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_10632 = _T_5041 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10823 = _T_10822 | _T_10632; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_10634 = _T_5045 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10824 = _T_10823 | _T_10634; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_10636 = _T_5049 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10825 = _T_10824 | _T_10636; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_10638 = _T_5053 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10826 = _T_10825 | _T_10638; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_10640 = _T_5057 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10827 = _T_10826 | _T_10640; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_10642 = _T_5061 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10828 = _T_10827 | _T_10642; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_10644 = _T_5065 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10829 = _T_10828 | _T_10644; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_10646 = _T_5069 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10830 = _T_10829 | _T_10646; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_10648 = _T_5073 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10831 = _T_10830 | _T_10648; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_10650 = _T_5077 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10832 = _T_10831 | _T_10650; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_10652 = _T_5081 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10833 = _T_10832 | _T_10652; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_10654 = _T_5085 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10834 = _T_10833 | _T_10654; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_10656 = _T_5089 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10835 = _T_10834 | _T_10656; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_10658 = _T_5093 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10836 = _T_10835 | _T_10658; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_10660 = _T_5097 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10837 = _T_10836 | _T_10660; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_10662 = _T_5101 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10838 = _T_10837 | _T_10662; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_10664 = _T_5105 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10839 = _T_10838 | _T_10664; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_10666 = _T_5109 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10840 = _T_10839 | _T_10666; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_10668 = _T_5113 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10841 = _T_10840 | _T_10668; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_10670 = _T_5117 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10842 = _T_10841 | _T_10670; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_10672 = _T_5121 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10843 = _T_10842 | _T_10672; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_10674 = _T_5125 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10844 = _T_10843 | _T_10674; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_10676 = _T_5129 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10845 = _T_10844 | _T_10676; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_10678 = _T_5133 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10846 = _T_10845 | _T_10678; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_10680 = _T_5137 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10847 = _T_10846 | _T_10680; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_10682 = _T_5141 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10848 = _T_10847 | _T_10682; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_10684 = _T_5145 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10849 = _T_10848 | _T_10684; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_10686 = _T_5149 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10850 = _T_10849 | _T_10686; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_10688 = _T_5153 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10851 = _T_10850 | _T_10688; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_10690 = _T_5157 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10852 = _T_10851 | _T_10690; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_10692 = _T_5161 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10853 = _T_10852 | _T_10692; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_10694 = _T_5165 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10854 = _T_10853 | _T_10694; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_10696 = _T_5169 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10855 = _T_10854 | _T_10696; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_10698 = _T_5173 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10856 = _T_10855 | _T_10698; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_10700 = _T_5177 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10857 = _T_10856 | _T_10700; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_10702 = _T_5181 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10858 = _T_10857 | _T_10702; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_10704 = _T_5185 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10859 = _T_10858 | _T_10704; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_10706 = _T_5189 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10860 = _T_10859 | _T_10706; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_10708 = _T_5193 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10861 = _T_10860 | _T_10708; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_10710 = _T_5197 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10862 = _T_10861 | _T_10710; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_10712 = _T_5201 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10863 = _T_10862 | _T_10712; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_10714 = _T_5205 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10864 = _T_10863 | _T_10714; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_10716 = _T_5209 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10865 = _T_10864 | _T_10716; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_10718 = _T_5213 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10866 = _T_10865 | _T_10718; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_10720 = _T_5217 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10867 = _T_10866 | _T_10720; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_10722 = _T_5221 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10868 = _T_10867 | _T_10722; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_10724 = _T_5225 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10869 = _T_10868 | _T_10724; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_10726 = _T_5229 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10870 = _T_10869 | _T_10726; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_10728 = _T_5233 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10871 = _T_10870 | _T_10728; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_10730 = _T_5237 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10872 = _T_10871 | _T_10730; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_10732 = _T_5241 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10873 = _T_10872 | _T_10732; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_10734 = _T_5245 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10874 = _T_10873 | _T_10734; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_10736 = _T_5249 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10875 = _T_10874 | _T_10736; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_10738 = _T_5253 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10876 = _T_10875 | _T_10738; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_10740 = _T_5257 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10877 = _T_10876 | _T_10740; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_10742 = _T_5261 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10878 = _T_10877 | _T_10742; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_10744 = _T_5265 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10879 = _T_10878 | _T_10744; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_10746 = _T_5269 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10880 = _T_10879 | _T_10746; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_10748 = _T_5273 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10881 = _T_10880 | _T_10748; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_10750 = _T_5277 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10882 = _T_10881 | _T_10750; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_10752 = _T_5281 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10883 = _T_10882 | _T_10752; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_10754 = _T_5285 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10884 = _T_10883 | _T_10754; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_10756 = _T_5289 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10885 = _T_10884 | _T_10756; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_10758 = _T_5293 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10886 = _T_10885 | _T_10758; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_10760 = _T_5297 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10887 = _T_10886 | _T_10760; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_10123 = _T_4789 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 764:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_10125 = _T_4793 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10378 = _T_10123 | _T_10125; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_10127 = _T_4797 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10379 = _T_10378 | _T_10127; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_10129 = _T_4801 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10380 = _T_10379 | _T_10129; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_10131 = _T_4805 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10381 = _T_10380 | _T_10131; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_10133 = _T_4809 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10382 = _T_10381 | _T_10133; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_10135 = _T_4813 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10383 = _T_10382 | _T_10135; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_10137 = _T_4817 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10384 = _T_10383 | _T_10137; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_10139 = _T_4821 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10385 = _T_10384 | _T_10139; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_10141 = _T_4825 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10386 = _T_10385 | _T_10141; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_10143 = _T_4829 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10387 = _T_10386 | _T_10143; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_10145 = _T_4833 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10388 = _T_10387 | _T_10145; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_10147 = _T_4837 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10389 = _T_10388 | _T_10147; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_10149 = _T_4841 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10390 = _T_10389 | _T_10149; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_10151 = _T_4845 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10391 = _T_10390 | _T_10151; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_10153 = _T_4849 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10392 = _T_10391 | _T_10153; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_10155 = _T_4853 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10393 = _T_10392 | _T_10155; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_10157 = _T_4857 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10394 = _T_10393 | _T_10157; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_10159 = _T_4861 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10395 = _T_10394 | _T_10159; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_10161 = _T_4865 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10396 = _T_10395 | _T_10161; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_10163 = _T_4869 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10397 = _T_10396 | _T_10163; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_10165 = _T_4873 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10398 = _T_10397 | _T_10165; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_10167 = _T_4877 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10399 = _T_10398 | _T_10167; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_10169 = _T_4881 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10400 = _T_10399 | _T_10169; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_10171 = _T_4885 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10401 = _T_10400 | _T_10171; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_10173 = _T_4889 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10402 = _T_10401 | _T_10173; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_10175 = _T_4893 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10403 = _T_10402 | _T_10175; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_10177 = _T_4897 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10404 = _T_10403 | _T_10177; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_10179 = _T_4901 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10405 = _T_10404 | _T_10179; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_10181 = _T_4905 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10406 = _T_10405 | _T_10181; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_10183 = _T_4909 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10407 = _T_10406 | _T_10183; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_10185 = _T_4913 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10408 = _T_10407 | _T_10185; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_10187 = _T_4917 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10409 = _T_10408 | _T_10187; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_10189 = _T_4921 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10410 = _T_10409 | _T_10189; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_10191 = _T_4925 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10411 = _T_10410 | _T_10191; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_10193 = _T_4929 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10412 = _T_10411 | _T_10193; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_10195 = _T_4933 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10413 = _T_10412 | _T_10195; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_10197 = _T_4937 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10414 = _T_10413 | _T_10197; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_10199 = _T_4941 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10415 = _T_10414 | _T_10199; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_10201 = _T_4945 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10416 = _T_10415 | _T_10201; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_10203 = _T_4949 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10417 = _T_10416 | _T_10203; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_10205 = _T_4953 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10418 = _T_10417 | _T_10205; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_10207 = _T_4957 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10419 = _T_10418 | _T_10207; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_10209 = _T_4961 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10420 = _T_10419 | _T_10209; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_10211 = _T_4965 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10421 = _T_10420 | _T_10211; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_10213 = _T_4969 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10422 = _T_10421 | _T_10213; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_10215 = _T_4973 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10423 = _T_10422 | _T_10215; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_10217 = _T_4977 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10424 = _T_10423 | _T_10217; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_10219 = _T_4981 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10425 = _T_10424 | _T_10219; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_10221 = _T_4985 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10426 = _T_10425 | _T_10221; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_10223 = _T_4989 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10427 = _T_10426 | _T_10223; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_10225 = _T_4993 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10428 = _T_10427 | _T_10225; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_10227 = _T_4997 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10429 = _T_10428 | _T_10227; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_10229 = _T_5001 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10430 = _T_10429 | _T_10229; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_10231 = _T_5005 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10431 = _T_10430 | _T_10231; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_10233 = _T_5009 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10432 = _T_10431 | _T_10233; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_10235 = _T_5013 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10433 = _T_10432 | _T_10235; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_10237 = _T_5017 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10434 = _T_10433 | _T_10237; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_10239 = _T_5021 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10435 = _T_10434 | _T_10239; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_10241 = _T_5025 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10436 = _T_10435 | _T_10241; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_10243 = _T_5029 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10437 = _T_10436 | _T_10243; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_10245 = _T_5033 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10438 = _T_10437 | _T_10245; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_10247 = _T_5037 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10439 = _T_10438 | _T_10247; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_10249 = _T_5041 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10440 = _T_10439 | _T_10249; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_10251 = _T_5045 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10441 = _T_10440 | _T_10251; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_10253 = _T_5049 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10442 = _T_10441 | _T_10253; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_10255 = _T_5053 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10443 = _T_10442 | _T_10255; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_10257 = _T_5057 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10444 = _T_10443 | _T_10257; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_10259 = _T_5061 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10445 = _T_10444 | _T_10259; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_10261 = _T_5065 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10446 = _T_10445 | _T_10261; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_10263 = _T_5069 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10447 = _T_10446 | _T_10263; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_10265 = _T_5073 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10448 = _T_10447 | _T_10265; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_10267 = _T_5077 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10449 = _T_10448 | _T_10267; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_10269 = _T_5081 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10450 = _T_10449 | _T_10269; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_10271 = _T_5085 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10451 = _T_10450 | _T_10271; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_10273 = _T_5089 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10452 = _T_10451 | _T_10273; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_10275 = _T_5093 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10453 = _T_10452 | _T_10275; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_10277 = _T_5097 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10454 = _T_10453 | _T_10277; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_10279 = _T_5101 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10455 = _T_10454 | _T_10279; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_10281 = _T_5105 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10456 = _T_10455 | _T_10281; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_10283 = _T_5109 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10457 = _T_10456 | _T_10283; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_10285 = _T_5113 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10458 = _T_10457 | _T_10285; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_10287 = _T_5117 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10459 = _T_10458 | _T_10287; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_10289 = _T_5121 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10460 = _T_10459 | _T_10289; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_10291 = _T_5125 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10461 = _T_10460 | _T_10291; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_10293 = _T_5129 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10462 = _T_10461 | _T_10293; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_10295 = _T_5133 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10463 = _T_10462 | _T_10295; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_10297 = _T_5137 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10464 = _T_10463 | _T_10297; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_10299 = _T_5141 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10465 = _T_10464 | _T_10299; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_10301 = _T_5145 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10466 = _T_10465 | _T_10301; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_10303 = _T_5149 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10467 = _T_10466 | _T_10303; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_10305 = _T_5153 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10468 = _T_10467 | _T_10305; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_10307 = _T_5157 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10469 = _T_10468 | _T_10307; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_10309 = _T_5161 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10470 = _T_10469 | _T_10309; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_10311 = _T_5165 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10471 = _T_10470 | _T_10311; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_10313 = _T_5169 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10472 = _T_10471 | _T_10313; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_10315 = _T_5173 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10473 = _T_10472 | _T_10315; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_10317 = _T_5177 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10474 = _T_10473 | _T_10317; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_10319 = _T_5181 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10475 = _T_10474 | _T_10319; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_10321 = _T_5185 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10476 = _T_10475 | _T_10321; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_10323 = _T_5189 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10477 = _T_10476 | _T_10323; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_10325 = _T_5193 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10478 = _T_10477 | _T_10325; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_10327 = _T_5197 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10479 = _T_10478 | _T_10327; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_10329 = _T_5201 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10480 = _T_10479 | _T_10329; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_10331 = _T_5205 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10481 = _T_10480 | _T_10331; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_10333 = _T_5209 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10482 = _T_10481 | _T_10333; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_10335 = _T_5213 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10483 = _T_10482 | _T_10335; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_10337 = _T_5217 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10484 = _T_10483 | _T_10337; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_10339 = _T_5221 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10485 = _T_10484 | _T_10339; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_10341 = _T_5225 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10486 = _T_10485 | _T_10341; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_10343 = _T_5229 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10487 = _T_10486 | _T_10343; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_10345 = _T_5233 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10488 = _T_10487 | _T_10345; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_10347 = _T_5237 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10489 = _T_10488 | _T_10347; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_10349 = _T_5241 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10490 = _T_10489 | _T_10349; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_10351 = _T_5245 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10491 = _T_10490 | _T_10351; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_10353 = _T_5249 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10492 = _T_10491 | _T_10353; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_10355 = _T_5253 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10493 = _T_10492 | _T_10355; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_10357 = _T_5257 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10494 = _T_10493 | _T_10357; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_10359 = _T_5261 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10495 = _T_10494 | _T_10359; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_10361 = _T_5265 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10496 = _T_10495 | _T_10361; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_10363 = _T_5269 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10497 = _T_10496 | _T_10363; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_10365 = _T_5273 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10498 = _T_10497 | _T_10365; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_10367 = _T_5277 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10499 = _T_10498 | _T_10367; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_10369 = _T_5281 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10500 = _T_10499 | _T_10369; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_10371 = _T_5285 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10501 = _T_10500 | _T_10371; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_10373 = _T_5289 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10502 = _T_10501 | _T_10373; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_10375 = _T_5293 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10503 = _T_10502 | _T_10375; // @[el2_ifu_mem_ctl.scala 764:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_10377 = _T_5297 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 764:10]
  wire  _T_10504 = _T_10503 | _T_10377; // @[el2_ifu_mem_ctl.scala 764:91]
  wire [1:0] ic_tag_valid_unq = {_T_10887,_T_10504}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 838:54]
  wire [1:0] _T_10927 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10928 = ic_debug_way_ff & _T_10927; // @[el2_ifu_mem_ctl.scala 819:67]
  wire [1:0] _T_10929 = ic_tag_valid_unq & _T_10928; // @[el2_ifu_mem_ctl.scala 819:48]
  wire  ic_debug_tag_val_rd_out = |_T_10929; // @[el2_ifu_mem_ctl.scala 819:115]
  wire [65:0] _T_1208 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1209; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2591; // @[el2_ifu_mem_ctl.scala 368:80]
  wire  _T_1247 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 373:98]
  wire  sel_byp_data = _T_1251 & _T_1247; // @[el2_ifu_mem_ctl.scala 373:96]
  wire [63:0] _T_1258 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1259 = _T_1258 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 380:64]
  wire [63:0] _T_1261 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2113 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 448:31]
  wire  _T_1626 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 444:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1627 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1675 = _T_1627 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1630 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1676 = _T_1630 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1675 | _T_1676; // @[Mux.scala 27:72]
  wire  _T_1633 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1677 = _T_1633 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1692 = _T_1691 | _T_1677; // @[Mux.scala 27:72]
  wire  _T_1636 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1678 = _T_1636 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1692 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1639 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1679 = _T_1639 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire  _T_1642 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1680 = _T_1642 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1695 = _T_1694 | _T_1680; // @[Mux.scala 27:72]
  wire  _T_1645 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1681 = _T_1645 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1696 = _T_1695 | _T_1681; // @[Mux.scala 27:72]
  wire  _T_1648 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1682 = _T_1648 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1697 = _T_1696 | _T_1682; // @[Mux.scala 27:72]
  wire  _T_1651 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1683 = _T_1651 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1698 = _T_1697 | _T_1683; // @[Mux.scala 27:72]
  wire  _T_1654 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1684 = _T_1654 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1699 = _T_1698 | _T_1684; // @[Mux.scala 27:72]
  wire  _T_1657 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1685 = _T_1657 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1700 = _T_1699 | _T_1685; // @[Mux.scala 27:72]
  wire  _T_1660 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1686 = _T_1660 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1701 = _T_1700 | _T_1686; // @[Mux.scala 27:72]
  wire  _T_1663 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1687 = _T_1663 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1702 = _T_1701 | _T_1687; // @[Mux.scala 27:72]
  wire  _T_1666 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1688 = _T_1666 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1703 = _T_1702 | _T_1688; // @[Mux.scala 27:72]
  wire  _T_1669 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1689 = _T_1669 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1704 = _T_1703 | _T_1689; // @[Mux.scala 27:72]
  wire  _T_1672 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 445:73]
  wire [15:0] _T_1690 = _T_1672 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1705 = _T_1704 | _T_1690; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1707 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1755 = _T_1707 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1710 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1756 = _T_1710 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1755 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1713 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1757 = _T_1713 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1772 = _T_1771 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1716 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1758 = _T_1716 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1772 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1719 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1759 = _T_1719 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1722 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1760 = _T_1722 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1775 = _T_1774 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1725 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1761 = _T_1725 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1776 = _T_1775 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1728 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1762 = _T_1728 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1777 = _T_1776 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1731 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1763 = _T_1731 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1778 = _T_1777 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1734 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1764 = _T_1734 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1779 = _T_1778 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1737 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1765 = _T_1737 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1780 = _T_1779 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1740 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1766 = _T_1740 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1781 = _T_1780 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1743 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1767 = _T_1743 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1782 = _T_1781 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1746 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1768 = _T_1746 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1783 = _T_1782 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1749 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1769 = _T_1749 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1784 = _T_1783 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1752 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 445:179]
  wire [31:0] _T_1770 = _T_1752 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1785 = _T_1784 | _T_1770; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1787 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1835 = _T_1787 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1790 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1836 = _T_1790 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1835 | _T_1836; // @[Mux.scala 27:72]
  wire  _T_1793 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1837 = _T_1793 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1852 = _T_1851 | _T_1837; // @[Mux.scala 27:72]
  wire  _T_1796 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1838 = _T_1796 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1852 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1799 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1839 = _T_1799 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire  _T_1802 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1840 = _T_1802 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1855 = _T_1854 | _T_1840; // @[Mux.scala 27:72]
  wire  _T_1805 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1841 = _T_1805 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1856 = _T_1855 | _T_1841; // @[Mux.scala 27:72]
  wire  _T_1808 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1842 = _T_1808 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1857 = _T_1856 | _T_1842; // @[Mux.scala 27:72]
  wire  _T_1811 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1843 = _T_1811 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1858 = _T_1857 | _T_1843; // @[Mux.scala 27:72]
  wire  _T_1814 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1844 = _T_1814 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1859 = _T_1858 | _T_1844; // @[Mux.scala 27:72]
  wire  _T_1817 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1845 = _T_1817 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1860 = _T_1859 | _T_1845; // @[Mux.scala 27:72]
  wire  _T_1820 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1846 = _T_1820 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1861 = _T_1860 | _T_1846; // @[Mux.scala 27:72]
  wire  _T_1823 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1847 = _T_1823 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1862 = _T_1861 | _T_1847; // @[Mux.scala 27:72]
  wire  _T_1826 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1848 = _T_1826 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1863 = _T_1862 | _T_1848; // @[Mux.scala 27:72]
  wire  _T_1829 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1849 = _T_1829 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1864 = _T_1863 | _T_1849; // @[Mux.scala 27:72]
  wire  _T_1832 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 445:285]
  wire [31:0] _T_1850 = _T_1832 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1865 = _T_1864 | _T_1850; // @[Mux.scala 27:72]
  wire [79:0] _T_1868 = {_T_1705,_T_1785,_T_1865}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1869 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1917 = _T_1869 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1918 = _T_1872 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1917 | _T_1918; // @[Mux.scala 27:72]
  wire  _T_1875 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1919 = _T_1875 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1934 = _T_1933 | _T_1919; // @[Mux.scala 27:72]
  wire  _T_1878 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1920 = _T_1878 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1934 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1881 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1921 = _T_1881 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire  _T_1884 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1922 = _T_1884 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1937 = _T_1936 | _T_1922; // @[Mux.scala 27:72]
  wire  _T_1887 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1923 = _T_1887 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1938 = _T_1937 | _T_1923; // @[Mux.scala 27:72]
  wire  _T_1890 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1924 = _T_1890 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1939 = _T_1938 | _T_1924; // @[Mux.scala 27:72]
  wire  _T_1893 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1925 = _T_1893 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1940 = _T_1939 | _T_1925; // @[Mux.scala 27:72]
  wire  _T_1896 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1926 = _T_1896 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1941 = _T_1940 | _T_1926; // @[Mux.scala 27:72]
  wire  _T_1899 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1927 = _T_1899 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1942 = _T_1941 | _T_1927; // @[Mux.scala 27:72]
  wire  _T_1902 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1928 = _T_1902 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1943 = _T_1942 | _T_1928; // @[Mux.scala 27:72]
  wire  _T_1905 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1929 = _T_1905 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1944 = _T_1943 | _T_1929; // @[Mux.scala 27:72]
  wire  _T_1908 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1930 = _T_1908 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1945 = _T_1944 | _T_1930; // @[Mux.scala 27:72]
  wire  _T_1911 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1931 = _T_1911 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1946 = _T_1945 | _T_1931; // @[Mux.scala 27:72]
  wire  _T_1914 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 446:73]
  wire [15:0] _T_1932 = _T_1914 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1947 = _T_1946 | _T_1932; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1627 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1630 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_1997 | _T_1998; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1633 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_2013 | _T_1999; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1636 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_2014 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1639 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1642 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2017 = _T_2016 | _T_2002; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_1645 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2018 = _T_2017 | _T_2003; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_1648 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2019 = _T_2018 | _T_2004; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_1651 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2020 = _T_2019 | _T_2005; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_1654 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2021 = _T_2020 | _T_2006; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_1657 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2022 = _T_2021 | _T_2007; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_1660 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2023 = _T_2022 | _T_2008; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_1663 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2024 = _T_2023 | _T_2009; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_1666 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2025 = _T_2024 | _T_2010; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_1669 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2026 = _T_2025 | _T_2011; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_1672 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2027 = _T_2026 | _T_2012; // @[Mux.scala 27:72]
  wire [79:0] _T_2110 = {_T_1947,_T_2027,_T_1785}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1626 ? _T_1868 : _T_2110; // @[el2_ifu_mem_ctl.scala 444:37]
  wire [79:0] _T_2115 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2113 ? ic_byp_data_only_pre_new : _T_2115; // @[el2_ifu_mem_ctl.scala 448:30]
  wire [79:0] _GEN_602 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 380:109]
  wire [79:0] _T_1262 = _GEN_602 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 380:109]
  wire [79:0] _GEN_603 = {{16'd0}, _T_1259}; // @[el2_ifu_mem_ctl.scala 380:83]
  wire [79:0] ic_premux_data = _GEN_603 | _T_1262; // @[el2_ifu_mem_ctl.scala 380:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 387:38]
  wire [1:0] _T_1271 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 391:8]
  wire  _T_1273 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 393:45]
  wire  _T_1275 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 393:80]
  wire  _T_1276 = ~_T_1275; // @[el2_ifu_mem_ctl.scala 393:71]
  wire  _T_1277 = _T_1273 & _T_1276; // @[el2_ifu_mem_ctl.scala 393:69]
  wire  _T_1278 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 393:131]
  wire  _T_1279 = _T_1277 & _T_1278; // @[el2_ifu_mem_ctl.scala 393:114]
  wire [7:0] _T_1368 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1373 = ic_miss_buff_data_error[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  _T_2659 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 624:47]
  wire  _T_2660 = _T_2659 & _T_13; // @[el2_ifu_mem_ctl.scala 624:50]
  wire  bus_ifu_wr_data_error = _T_2660 & miss_pending; // @[el2_ifu_mem_ctl.scala 624:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1373; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1377 = ic_miss_buff_data_error[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1377; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1381 = ic_miss_buff_data_error[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1381; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1385 = ic_miss_buff_data_error[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1385; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1389 = ic_miss_buff_data_error[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1389; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1393 = ic_miss_buff_data_error[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1393; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1397 = ic_miss_buff_data_error[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1397; // @[el2_ifu_mem_ctl.scala 410:72]
  wire  _T_1401 = ic_miss_buff_data_error[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 411:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1401; // @[el2_ifu_mem_ctl.scala 410:72]
  wire [7:0] _T_1408 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2465 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2473 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 493:65]
  wire  _T_2474 = _T_2473 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 493:88]
  wire  _T_2476 = _T_2474 & _T_2587; // @[el2_ifu_mem_ctl.scala 493:112]
  wire  _T_2477 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2478 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 498:50]
  wire  _T_2480 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2486 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2488 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_2486 | _T_2488; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2480 ? _T_2478 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_2477 ? _T_2478 : _GEN_41; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2465 ? _T_2476 : _GEN_43; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2465 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2479 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 499:56]
  wire  _GEN_44 = _T_2477 & _T_2479; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2465 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 484:58]
  wire  _T_2462 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 483:49]
  wire  _T_2467 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 492:87]
  wire  _T_2481 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 502:54]
  wire  _T_2482 = _T_2481 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 502:84]
  wire  _T_2491 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 523:66]
  wire  _T_2492 = io_dec_tlu_flush_err_wb & _T_2491; // @[el2_ifu_mem_ctl.scala 523:52]
  wire  _T_2494 = _T_2492 & _T_2587; // @[el2_ifu_mem_ctl.scala 523:81]
  wire  _T_2496 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 526:59]
  wire  _T_2497 = _T_2496 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 526:86]
  wire  _T_2511 = _T_2496 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 529:81]
  wire  _T_2512 = _T_2511 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 529:103]
  wire  _T_2513 = _T_2512 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 529:126]
  wire  _T_2533 = _T_2511 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 536:103]
  wire  _T_2540 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 541:62]
  wire  _T_2541 = io_dec_tlu_flush_lower_wb & _T_2540; // @[el2_ifu_mem_ctl.scala 541:60]
  wire  _T_2542 = _T_2541 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 541:88]
  wire  _T_2543 = _T_2542 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 541:115]
  wire  _GEN_51 = _T_2539 & _T_2497; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_2522 ? _T_2533 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_2522 | _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2495 ? _T_2513 : _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_2495 | _GEN_56; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2490 ? _T_2494 : _GEN_58; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2555 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 558:64]
  wire  _T_2557 = _T_2555 & _T_2587; // @[el2_ifu_mem_ctl.scala 558:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2559 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 558:133]
  wire  _T_2560 = _T_2559 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 558:164]
  wire  _T_2561 = _T_2560 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 558:184]
  wire  _T_2562 = _T_2561 & miss_pending; // @[el2_ifu_mem_ctl.scala 558:204]
  wire  _T_2563 = ~_T_2562; // @[el2_ifu_mem_ctl.scala 558:112]
  wire  ifc_bus_ic_req_ff_in = _T_2557 & _T_2563; // @[el2_ifu_mem_ctl.scala 558:110]
  wire  _T_2564 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 559:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 590:45]
  wire  _T_2581 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 593:35]
  wire  _T_2582 = _T_2581 & miss_pending; // @[el2_ifu_mem_ctl.scala 593:53]
  wire  bus_cmd_sent = _T_2582 & _T_2587; // @[el2_ifu_mem_ctl.scala 593:68]
  wire [2:0] _T_2572 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2574 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2576 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 591:51]
  wire  _T_2602 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 601:73]
  wire  _T_2603 = _T_2588 & _T_2602; // @[el2_ifu_mem_ctl.scala 601:71]
  wire  _T_2605 = last_data_recieved_ff & _T_1339; // @[el2_ifu_mem_ctl.scala 601:114]
  wire  last_data_recieved_in = _T_2603 | _T_2605; // @[el2_ifu_mem_ctl.scala 601:89]
  wire [2:0] _T_2611 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 606:45]
  wire  _T_2614 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 607:81]
  wire  _T_2615 = _T_2614 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 607:97]
  wire  _T_2617 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 609:48]
  wire  _T_2618 = _T_2617 & miss_pending; // @[el2_ifu_mem_ctl.scala 609:68]
  wire  bus_inc_cmd_beat_cnt = _T_2618 & _T_2587; // @[el2_ifu_mem_ctl.scala 609:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 611:57]
  wire  _T_2622 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 612:31]
  wire  _T_2623 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 612:71]
  wire  _T_2624 = _T_2623 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 612:87]
  wire  _T_2625 = ~_T_2624; // @[el2_ifu_mem_ctl.scala 612:55]
  wire  bus_hold_cmd_beat_cnt = _T_2622 & _T_2625; // @[el2_ifu_mem_ctl.scala 612:53]
  wire  _T_2626 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 613:46]
  wire  bus_cmd_beat_en = _T_2626 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 613:62]
  wire [2:0] _T_2629 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 615:46]
  wire [2:0] _T_2631 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2632 = bus_inc_cmd_beat_cnt ? _T_2629 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2633 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2635 = _T_2631 | _T_2632; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2635 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2639 = _T_2615 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 616:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 627:62]
  wire  _T_2667 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 632:50]
  wire  _T_2668 = io_ifc_dma_access_ok & _T_2667; // @[el2_ifu_mem_ctl.scala 632:47]
  wire  _T_2669 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 632:70]
  wire  ifc_dma_access_ok_d = _T_2668 & _T_2669; // @[el2_ifu_mem_ctl.scala 632:68]
  wire  _T_2673 = _T_2668 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 633:72]
  wire  _T_2674 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 633:111]
  wire  _T_2675 = _T_2673 & _T_2674; // @[el2_ifu_mem_ctl.scala 633:97]
  wire  ifc_dma_access_q_ok = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 633:127]
  wire  _T_2678 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 636:40]
  wire  _T_2679 = _T_2678 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 636:58]
  wire  _T_2682 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 637:60]
  wire  _T_2683 = _T_2678 & _T_2682; // @[el2_ifu_mem_ctl.scala 637:58]
  wire  _T_2684 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 637:104]
  wire [2:0] _T_2689 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2795 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2804 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2795}; // @[el2_lib.scala 268:22]
  wire  _T_2805 = ^_T_2804; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2813 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2822 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2813}; // @[el2_lib.scala 268:39]
  wire  _T_2823 = ^_T_2822; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2831 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2840 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2831}; // @[el2_lib.scala 268:56]
  wire  _T_2841 = ^_T_2840; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2847 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2855 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2847}; // @[el2_lib.scala 268:73]
  wire  _T_2856 = ^_T_2855; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2870 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2847}; // @[el2_lib.scala 268:90]
  wire  _T_2871 = ^_T_2870; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2876 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2877 = ^_T_2876; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2882 = {_T_2805,_T_2823,_T_2841,_T_2856,_T_2871,_T_2877}; // @[Cat.scala 29:58]
  wire  _T_2883 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2884 = ^_T_2882; // @[el2_lib.scala 269:23]
  wire  _T_2885 = _T_2883 ^ _T_2884; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2991 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_3000 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2991}; // @[el2_lib.scala 268:22]
  wire  _T_3001 = ^_T_3000; // @[el2_lib.scala 268:29]
  wire [8:0] _T_3009 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_3018 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_3009}; // @[el2_lib.scala 268:39]
  wire  _T_3019 = ^_T_3018; // @[el2_lib.scala 268:46]
  wire [8:0] _T_3027 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_3036 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_3027}; // @[el2_lib.scala 268:56]
  wire  _T_3037 = ^_T_3036; // @[el2_lib.scala 268:63]
  wire [6:0] _T_3043 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_3051 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_3043}; // @[el2_lib.scala 268:73]
  wire  _T_3052 = ^_T_3051; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3066 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_3043}; // @[el2_lib.scala 268:90]
  wire  _T_3067 = ^_T_3066; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3072 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3073 = ^_T_3072; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3078 = {_T_3001,_T_3019,_T_3037,_T_3052,_T_3067,_T_3073}; // @[Cat.scala 29:58]
  wire  _T_3079 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3080 = ^_T_3078; // @[el2_lib.scala 269:23]
  wire  _T_3081 = _T_3079 ^ _T_3080; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3082 = {_T_3081,_T_3001,_T_3019,_T_3037,_T_3052,_T_3067,_T_3073}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2885,_T_2805,_T_2823,_T_2841,_T_2856,_T_2871,_T_2877,_T_3082}; // @[Cat.scala 29:58]
  wire  _T_3084 = ~_T_2678; // @[el2_ifu_mem_ctl.scala 642:45]
  wire  _T_3085 = iccm_correct_ecc & _T_3084; // @[el2_ifu_mem_ctl.scala 642:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3086 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3093 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 656:53]
  wire  _T_3425 = _T_3337[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3423 = _T_3337[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3421 = _T_3337[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3419 = _T_3337[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3417 = _T_3337[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3415 = _T_3337[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3413 = _T_3337[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3411 = _T_3337[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3409 = _T_3337[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3407 = _T_3337[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3483 = {_T_3425,_T_3423,_T_3421,_T_3419,_T_3417,_T_3415,_T_3413,_T_3411,_T_3409,_T_3407}; // @[el2_lib.scala 310:69]
  wire  _T_3405 = _T_3337[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3403 = _T_3337[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3401 = _T_3337[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3399 = _T_3337[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3397 = _T_3337[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3395 = _T_3337[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3393 = _T_3337[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3391 = _T_3337[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3389 = _T_3337[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3387 = _T_3337[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3474 = {_T_3405,_T_3403,_T_3401,_T_3399,_T_3397,_T_3395,_T_3393,_T_3391,_T_3389,_T_3387}; // @[el2_lib.scala 310:69]
  wire  _T_3385 = _T_3337[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3383 = _T_3337[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3381 = _T_3337[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3379 = _T_3337[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3377 = _T_3337[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3375 = _T_3337[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3373 = _T_3337[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3371 = _T_3337[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3369 = _T_3337[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3367 = _T_3337[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3464 = {_T_3385,_T_3383,_T_3381,_T_3379,_T_3377,_T_3375,_T_3373,_T_3371,_T_3369,_T_3367}; // @[el2_lib.scala 310:69]
  wire  _T_3365 = _T_3337[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3363 = _T_3337[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3361 = _T_3337[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3359 = _T_3337[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3357 = _T_3337[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3355 = _T_3337[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3353 = _T_3337[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3351 = _T_3337[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3349 = _T_3337[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3465 = {_T_3464,_T_3365,_T_3363,_T_3361,_T_3359,_T_3357,_T_3355,_T_3353,_T_3351,_T_3349}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3485 = {_T_3483,_T_3474,_T_3465}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3440 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3446 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3440}; // @[Cat.scala 29:58]
  wire [38:0] _T_3486 = _T_3485 ^ _T_3446; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3487 = _T_3341 ? _T_3486 : _T_3446; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3487[37:32],_T_3487[30:16],_T_3487[14:8],_T_3487[6:4],_T_3487[2]}; // @[Cat.scala 29:58]
  wire  _T_3810 = _T_3722[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3808 = _T_3722[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3806 = _T_3722[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3804 = _T_3722[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3802 = _T_3722[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3800 = _T_3722[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3798 = _T_3722[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3796 = _T_3722[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3794 = _T_3722[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3792 = _T_3722[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3868 = {_T_3810,_T_3808,_T_3806,_T_3804,_T_3802,_T_3800,_T_3798,_T_3796,_T_3794,_T_3792}; // @[el2_lib.scala 310:69]
  wire  _T_3790 = _T_3722[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3788 = _T_3722[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3786 = _T_3722[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3784 = _T_3722[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3782 = _T_3722[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3780 = _T_3722[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3778 = _T_3722[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3776 = _T_3722[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3774 = _T_3722[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3772 = _T_3722[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3859 = {_T_3790,_T_3788,_T_3786,_T_3784,_T_3782,_T_3780,_T_3778,_T_3776,_T_3774,_T_3772}; // @[el2_lib.scala 310:69]
  wire  _T_3770 = _T_3722[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3768 = _T_3722[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3766 = _T_3722[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3764 = _T_3722[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3762 = _T_3722[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3760 = _T_3722[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3758 = _T_3722[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3756 = _T_3722[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3754 = _T_3722[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3752 = _T_3722[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3849 = {_T_3770,_T_3768,_T_3766,_T_3764,_T_3762,_T_3760,_T_3758,_T_3756,_T_3754,_T_3752}; // @[el2_lib.scala 310:69]
  wire  _T_3750 = _T_3722[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3748 = _T_3722[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3746 = _T_3722[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3744 = _T_3722[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3742 = _T_3722[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3740 = _T_3722[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3738 = _T_3722[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3736 = _T_3722[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3734 = _T_3722[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3850 = {_T_3849,_T_3750,_T_3748,_T_3746,_T_3744,_T_3742,_T_3740,_T_3738,_T_3736,_T_3734}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3870 = {_T_3868,_T_3859,_T_3850}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3825 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3831 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3825}; // @[Cat.scala 29:58]
  wire [38:0] _T_3871 = _T_3870 ^ _T_3831; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3872 = _T_3726 ? _T_3871 : _T_3831; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3872[37:32],_T_3872[30:16],_T_3872[14:8],_T_3872[6:4],_T_3872[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 648:35]
  wire  _T_3345 = ~_T_3337[6]; // @[el2_lib.scala 303:55]
  wire  _T_3346 = _T_3339 & _T_3345; // @[el2_lib.scala 303:53]
  wire  _T_3730 = ~_T_3722[6]; // @[el2_lib.scala 303:55]
  wire  _T_3731 = _T_3724 & _T_3730; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3346,_T_3731}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 650:53]
  wire [63:0] _T_3097 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3098 = {iccm_dma_rdata_1_muxed,_T_3487[37:32],_T_3487[30:16],_T_3487[14:8],_T_3487[6:4],_T_3487[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 652:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 653:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 658:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 662:70]
  wire  _T_3103 = _T_2678 & _T_2667; // @[el2_ifu_mem_ctl.scala 665:65]
  wire  _T_3106 = _T_3084 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 666:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3107 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3109 = _T_3106 ? {{1'd0}, _T_3107} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 666:8]
  wire [31:0] _T_3110 = _T_3103 ? io_dma_mem_addr : {{16'd0}, _T_3109}; // @[el2_ifu_mem_ctl.scala 665:25]
  wire  _T_3499 = _T_3337 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3500 = _T_3487[38] ^ _T_3499; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3500,_T_3487[31],_T_3487[15],_T_3487[7],_T_3487[3],_T_3487[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3884 = _T_3722 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3885 = _T_3872[38] ^ _T_3884; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3885,_T_3872[31],_T_3872[15],_T_3872[7],_T_3872[3],_T_3872[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3901 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 678:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 680:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 681:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 689:62]
  wire  _T_3909 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 683:76]
  wire  _T_3910 = io_iccm_rd_ecc_single_err & _T_3909; // @[el2_ifu_mem_ctl.scala 683:74]
  wire  _T_3912 = _T_3910 & _T_317; // @[el2_ifu_mem_ctl.scala 683:104]
  wire  iccm_ecc_write_status = _T_3912 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 683:127]
  wire  _T_3913 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 684:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3913 & _T_317; // @[el2_ifu_mem_ctl.scala 684:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 688:51]
  wire [13:0] _T_3918 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 687:102]
  wire [38:0] _T_3922 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3927 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 692:41]
  wire  _T_3928 = io_ifc_fetch_req_bf & _T_3927; // @[el2_ifu_mem_ctl.scala 692:39]
  wire  _T_3929 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 692:72]
  wire  _T_3930 = _T_3928 & _T_3929; // @[el2_ifu_mem_ctl.scala 692:70]
  wire  _T_3932 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 693:34]
  wire  _T_3933 = _T_2233 & _T_3932; // @[el2_ifu_mem_ctl.scala 693:32]
  wire  _T_3936 = _T_2249 & _T_3932; // @[el2_ifu_mem_ctl.scala 694:37]
  wire  _T_3937 = _T_3933 | _T_3936; // @[el2_ifu_mem_ctl.scala 693:88]
  wire  _T_3938 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 695:19]
  wire  _T_3940 = _T_3938 & _T_3932; // @[el2_ifu_mem_ctl.scala 695:41]
  wire  _T_3941 = _T_3937 | _T_3940; // @[el2_ifu_mem_ctl.scala 694:88]
  wire  _T_3942 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 696:19]
  wire  _T_3944 = _T_3942 & _T_3932; // @[el2_ifu_mem_ctl.scala 696:35]
  wire  _T_3945 = _T_3941 | _T_3944; // @[el2_ifu_mem_ctl.scala 695:88]
  wire  _T_3948 = _T_2248 & _T_3932; // @[el2_ifu_mem_ctl.scala 697:38]
  wire  _T_3949 = _T_3945 | _T_3948; // @[el2_ifu_mem_ctl.scala 696:88]
  wire  _T_3951 = _T_2249 & miss_state_en; // @[el2_ifu_mem_ctl.scala 698:37]
  wire  _T_3952 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 698:71]
  wire  _T_3953 = _T_3951 & _T_3952; // @[el2_ifu_mem_ctl.scala 698:54]
  wire  _T_3954 = _T_3949 | _T_3953; // @[el2_ifu_mem_ctl.scala 697:57]
  wire  _T_3955 = ~_T_3954; // @[el2_ifu_mem_ctl.scala 693:5]
  wire  _T_3956 = _T_3930 & _T_3955; // @[el2_ifu_mem_ctl.scala 692:96]
  wire  _T_3957 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 699:28]
  wire  _T_3959 = _T_3957 & _T_3927; // @[el2_ifu_mem_ctl.scala 699:50]
  wire  _T_3961 = _T_3959 & _T_3929; // @[el2_ifu_mem_ctl.scala 699:81]
  wire [1:0] _T_3964 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10912 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 796:74]
  wire  bus_wren_1 = _T_10912 & miss_pending; // @[el2_ifu_mem_ctl.scala 796:98]
  wire  _T_10911 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 796:74]
  wire  bus_wren_0 = _T_10911 & miss_pending; // @[el2_ifu_mem_ctl.scala 796:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3970 = ~_T_108; // @[el2_ifu_mem_ctl.scala 702:106]
  wire  _T_3971 = _T_2233 & _T_3970; // @[el2_ifu_mem_ctl.scala 702:104]
  wire  _T_3972 = _T_2249 | _T_3971; // @[el2_ifu_mem_ctl.scala 702:77]
  wire  _T_3976 = ~_T_51; // @[el2_ifu_mem_ctl.scala 702:172]
  wire  _T_3977 = _T_3972 & _T_3976; // @[el2_ifu_mem_ctl.scala 702:170]
  wire  _T_3978 = ~_T_3977; // @[el2_ifu_mem_ctl.scala 702:44]
  wire  _T_3982 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 705:64]
  wire  _T_3983 = ~_T_3982; // @[el2_ifu_mem_ctl.scala 705:50]
  wire  _T_3984 = _T_276 & _T_3983; // @[el2_ifu_mem_ctl.scala 705:48]
  wire  _T_3985 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 705:81]
  wire  ic_valid = _T_3984 & _T_3985; // @[el2_ifu_mem_ctl.scala 705:79]
  wire  _T_3987 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 706:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 709:14]
  wire  _T_3990 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 712:74]
  wire  _T_10909 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 795:45]
  wire  way_status_wr_en = _T_10909 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 795:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3990; // @[el2_ifu_mem_ctl.scala 712:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 714:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 791:41]
  wire  way_status_new = _T_10909 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 794:26]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 722:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 724:132]
  wire  _T_4010 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4011 = _T_4010 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4012 = _T_4011 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4015 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4016 = _T_4015 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4017 = _T_4016 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4020 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4021 = _T_4020 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4022 = _T_4021 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4025 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4026 = _T_4025 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4027 = _T_4026 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4030 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4031 = _T_4030 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4032 = _T_4031 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4035 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4036 = _T_4035 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4037 = _T_4036 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4040 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4041 = _T_4040 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4042 = _T_4041 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4045 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 728:100]
  wire  _T_4046 = _T_4045 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 728:108]
  wire  _T_4047 = _T_4046 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4052 = _T_4011 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4057 = _T_4016 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4062 = _T_4021 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4067 = _T_4026 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4072 = _T_4031 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4077 = _T_4036 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4082 = _T_4041 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4087 = _T_4046 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4092 = _T_4011 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4097 = _T_4016 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4102 = _T_4021 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4107 = _T_4026 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4112 = _T_4031 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4117 = _T_4036 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4122 = _T_4041 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4127 = _T_4046 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4132 = _T_4011 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4137 = _T_4016 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4142 = _T_4021 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4147 = _T_4026 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4152 = _T_4031 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4157 = _T_4036 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4162 = _T_4041 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4167 = _T_4046 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4172 = _T_4011 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4177 = _T_4016 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4182 = _T_4021 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4187 = _T_4026 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4192 = _T_4031 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4197 = _T_4036 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4202 = _T_4041 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4207 = _T_4046 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4212 = _T_4011 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4217 = _T_4016 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4222 = _T_4021 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4227 = _T_4026 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4232 = _T_4031 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4237 = _T_4036 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4242 = _T_4041 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4247 = _T_4046 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4252 = _T_4011 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4257 = _T_4016 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4262 = _T_4021 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4267 = _T_4026 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4272 = _T_4031 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4277 = _T_4036 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4282 = _T_4041 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4287 = _T_4046 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4292 = _T_4011 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4297 = _T_4016 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4302 = _T_4021 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4307 = _T_4026 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4312 = _T_4031 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4317 = _T_4036 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4322 = _T_4041 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4327 = _T_4046 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4332 = _T_4011 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4337 = _T_4016 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4342 = _T_4021 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4347 = _T_4026 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4352 = _T_4031 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4357 = _T_4036 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4362 = _T_4041 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4367 = _T_4046 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4372 = _T_4011 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4377 = _T_4016 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4382 = _T_4021 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4387 = _T_4026 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4392 = _T_4031 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4397 = _T_4036 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4402 = _T_4041 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4407 = _T_4046 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4412 = _T_4011 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4417 = _T_4016 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4422 = _T_4021 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4427 = _T_4026 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4432 = _T_4031 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4437 = _T_4036 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4442 = _T_4041 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4447 = _T_4046 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4452 = _T_4011 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4457 = _T_4016 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4462 = _T_4021 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4467 = _T_4026 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4472 = _T_4031 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4477 = _T_4036 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4482 = _T_4041 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4487 = _T_4046 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4492 = _T_4011 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4497 = _T_4016 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4502 = _T_4021 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4507 = _T_4026 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4512 = _T_4031 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4517 = _T_4036 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4522 = _T_4041 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4527 = _T_4046 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4532 = _T_4011 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4537 = _T_4016 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4542 = _T_4021 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4547 = _T_4026 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4552 = _T_4031 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4557 = _T_4036 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4562 = _T_4041 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4567 = _T_4046 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4572 = _T_4011 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4577 = _T_4016 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4582 = _T_4021 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4587 = _T_4026 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4592 = _T_4031 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4597 = _T_4036 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4602 = _T_4041 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4607 = _T_4046 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4612 = _T_4011 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4617 = _T_4016 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4622 = _T_4021 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4627 = _T_4026 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4632 = _T_4031 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4637 = _T_4036 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4642 = _T_4041 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire  _T_4647 = _T_4046 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 728:131]
  wire [9:0] _T_4657 = {way_status_out_127,way_status_out_126,way_status_out_125,way_status_out_124,way_status_out_123,way_status_out_122,way_status_out_121,way_status_out_120,way_status_out_119,way_status_out_118}; // @[Cat.scala 29:58]
  wire [18:0] _T_4666 = {_T_4657,way_status_out_117,way_status_out_116,way_status_out_115,way_status_out_114,way_status_out_113,way_status_out_112,way_status_out_111,way_status_out_110,way_status_out_109}; // @[Cat.scala 29:58]
  wire [27:0] _T_4675 = {_T_4666,way_status_out_108,way_status_out_107,way_status_out_106,way_status_out_105,way_status_out_104,way_status_out_103,way_status_out_102,way_status_out_101,way_status_out_100}; // @[Cat.scala 29:58]
  wire [36:0] _T_4684 = {_T_4675,way_status_out_99,way_status_out_98,way_status_out_97,way_status_out_96,way_status_out_95,way_status_out_94,way_status_out_93,way_status_out_92,way_status_out_91}; // @[Cat.scala 29:58]
  wire [45:0] _T_4693 = {_T_4684,way_status_out_90,way_status_out_89,way_status_out_88,way_status_out_87,way_status_out_86,way_status_out_85,way_status_out_84,way_status_out_83,way_status_out_82}; // @[Cat.scala 29:58]
  wire [54:0] _T_4702 = {_T_4693,way_status_out_81,way_status_out_80,way_status_out_79,way_status_out_78,way_status_out_77,way_status_out_76,way_status_out_75,way_status_out_74,way_status_out_73}; // @[Cat.scala 29:58]
  wire [63:0] _T_4711 = {_T_4702,way_status_out_72,way_status_out_71,way_status_out_70,way_status_out_69,way_status_out_68,way_status_out_67,way_status_out_66,way_status_out_65,way_status_out_64}; // @[Cat.scala 29:58]
  wire [72:0] _T_4720 = {_T_4711,way_status_out_63,way_status_out_62,way_status_out_61,way_status_out_60,way_status_out_59,way_status_out_58,way_status_out_57,way_status_out_56,way_status_out_55}; // @[Cat.scala 29:58]
  wire [81:0] _T_4729 = {_T_4720,way_status_out_54,way_status_out_53,way_status_out_52,way_status_out_51,way_status_out_50,way_status_out_49,way_status_out_48,way_status_out_47,way_status_out_46}; // @[Cat.scala 29:58]
  wire [90:0] _T_4738 = {_T_4729,way_status_out_45,way_status_out_44,way_status_out_43,way_status_out_42,way_status_out_41,way_status_out_40,way_status_out_39,way_status_out_38,way_status_out_37}; // @[Cat.scala 29:58]
  wire [99:0] _T_4747 = {_T_4738,way_status_out_36,way_status_out_35,way_status_out_34,way_status_out_33,way_status_out_32,way_status_out_31,way_status_out_30,way_status_out_29,way_status_out_28}; // @[Cat.scala 29:58]
  wire [108:0] _T_4756 = {_T_4747,way_status_out_27,way_status_out_26,way_status_out_25,way_status_out_24,way_status_out_23,way_status_out_22,way_status_out_21,way_status_out_20,way_status_out_19}; // @[Cat.scala 29:58]
  wire [117:0] _T_4765 = {_T_4756,way_status_out_18,way_status_out_17,way_status_out_16,way_status_out_15,way_status_out_14,way_status_out_13,way_status_out_12,way_status_out_11,way_status_out_10}; // @[Cat.scala 29:58]
  wire [126:0] _T_4774 = {_T_4765,way_status_out_9,way_status_out_8,way_status_out_7,way_status_out_6,way_status_out_5,way_status_out_4,way_status_out_3,way_status_out_2,way_status_out_1}; // @[Cat.scala 29:58]
  wire [9:0] _T_4783 = {way_status_clken_15,way_status_clken_14,way_status_clken_13,way_status_clken_12,way_status_clken_11,way_status_clken_10,way_status_clken_9,way_status_clken_8,way_status_clken_7,way_status_clken_6}; // @[Cat.scala 29:58]
  wire [14:0] _T_4788 = {_T_4783,way_status_clken_5,way_status_clken_4,way_status_clken_3,way_status_clken_2,way_status_clken_1}; // @[Cat.scala 29:58]
  wire  _T_10915 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 798:84]
  wire  _T_10916 = _T_10915 & miss_pending; // @[el2_ifu_mem_ctl.scala 798:108]
  wire  bus_wren_last_1 = _T_10916 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 798:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 799:84]
  wire  _T_10918 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 800:73]
  wire  _T_10913 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 798:84]
  wire  _T_10914 = _T_10913 & miss_pending; // @[el2_ifu_mem_ctl.scala 798:108]
  wire  bus_wren_last_0 = _T_10914 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 798:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 799:84]
  wire  _T_10917 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 800:73]
  wire [1:0] ifu_tag_wren = {_T_10918,_T_10917}; // @[Cat.scala 29:58]
  wire [1:0] _T_10953 = _T_3990 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10953 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 834:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 741:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 743:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 747:14]
  wire  _T_5436 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 751:78]
  wire  _T_5438 = _T_5436 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5440 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 752:70]
  wire  _T_5442 = _T_5440 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5443 = _T_5438 | _T_5442; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5444 = _T_5443 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire  _T_5448 = _T_5436 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5452 = _T_5440 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5453 = _T_5448 | _T_5452; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5454 = _T_5453 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire [1:0] tag_valid_clken_0 = {_T_5454,_T_5444}; // @[Cat.scala 29:58]
  wire  _T_5456 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 751:78]
  wire  _T_5458 = _T_5456 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5460 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 752:70]
  wire  _T_5462 = _T_5460 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5463 = _T_5458 | _T_5462; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5464 = _T_5463 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire  _T_5468 = _T_5456 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5472 = _T_5460 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5473 = _T_5468 | _T_5472; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5474 = _T_5473 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire [1:0] tag_valid_clken_1 = {_T_5474,_T_5464}; // @[Cat.scala 29:58]
  wire  _T_5476 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 751:78]
  wire  _T_5478 = _T_5476 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5480 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 752:70]
  wire  _T_5482 = _T_5480 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5483 = _T_5478 | _T_5482; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5484 = _T_5483 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire  _T_5488 = _T_5476 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5492 = _T_5480 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5493 = _T_5488 | _T_5492; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5494 = _T_5493 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire [1:0] tag_valid_clken_2 = {_T_5494,_T_5484}; // @[Cat.scala 29:58]
  wire  _T_5496 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 751:78]
  wire  _T_5498 = _T_5496 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5500 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 752:70]
  wire  _T_5502 = _T_5500 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5503 = _T_5498 | _T_5502; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5504 = _T_5503 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire  _T_5508 = _T_5496 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 751:87]
  wire  _T_5512 = _T_5500 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 752:79]
  wire  _T_5513 = _T_5508 | _T_5512; // @[el2_ifu_mem_ctl.scala 751:109]
  wire  _T_5514 = _T_5513 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 752:102]
  wire [1:0] tag_valid_clken_3 = {_T_5514,_T_5504}; // @[Cat.scala 29:58]
  wire [9:0] _T_5523 = {ic_tag_valid_out_1_127,ic_tag_valid_out_1_126,ic_tag_valid_out_1_125,ic_tag_valid_out_1_124,ic_tag_valid_out_1_123,ic_tag_valid_out_1_122,ic_tag_valid_out_1_121,ic_tag_valid_out_1_120,ic_tag_valid_out_1_119,ic_tag_valid_out_1_118}; // @[Cat.scala 29:58]
  wire [18:0] _T_5532 = {_T_5523,ic_tag_valid_out_1_117,ic_tag_valid_out_1_116,ic_tag_valid_out_1_115,ic_tag_valid_out_1_114,ic_tag_valid_out_1_113,ic_tag_valid_out_1_112,ic_tag_valid_out_1_111,ic_tag_valid_out_1_110,ic_tag_valid_out_1_109}; // @[Cat.scala 29:58]
  wire [27:0] _T_5541 = {_T_5532,ic_tag_valid_out_1_108,ic_tag_valid_out_1_107,ic_tag_valid_out_1_106,ic_tag_valid_out_1_105,ic_tag_valid_out_1_104,ic_tag_valid_out_1_103,ic_tag_valid_out_1_102,ic_tag_valid_out_1_101,ic_tag_valid_out_1_100}; // @[Cat.scala 29:58]
  wire [36:0] _T_5550 = {_T_5541,ic_tag_valid_out_1_99,ic_tag_valid_out_1_98,ic_tag_valid_out_1_97,ic_tag_valid_out_1_96,ic_tag_valid_out_1_95,ic_tag_valid_out_1_94,ic_tag_valid_out_1_93,ic_tag_valid_out_1_92,ic_tag_valid_out_1_91}; // @[Cat.scala 29:58]
  wire [45:0] _T_5559 = {_T_5550,ic_tag_valid_out_1_90,ic_tag_valid_out_1_89,ic_tag_valid_out_1_88,ic_tag_valid_out_1_87,ic_tag_valid_out_1_86,ic_tag_valid_out_1_85,ic_tag_valid_out_1_84,ic_tag_valid_out_1_83,ic_tag_valid_out_1_82}; // @[Cat.scala 29:58]
  wire [54:0] _T_5568 = {_T_5559,ic_tag_valid_out_1_81,ic_tag_valid_out_1_80,ic_tag_valid_out_1_79,ic_tag_valid_out_1_78,ic_tag_valid_out_1_77,ic_tag_valid_out_1_76,ic_tag_valid_out_1_75,ic_tag_valid_out_1_74,ic_tag_valid_out_1_73}; // @[Cat.scala 29:58]
  wire [63:0] _T_5577 = {_T_5568,ic_tag_valid_out_1_72,ic_tag_valid_out_1_71,ic_tag_valid_out_1_70,ic_tag_valid_out_1_69,ic_tag_valid_out_1_68,ic_tag_valid_out_1_67,ic_tag_valid_out_1_66,ic_tag_valid_out_1_65,ic_tag_valid_out_1_64}; // @[Cat.scala 29:58]
  wire [72:0] _T_5586 = {_T_5577,ic_tag_valid_out_1_63,ic_tag_valid_out_1_62,ic_tag_valid_out_1_61,ic_tag_valid_out_1_60,ic_tag_valid_out_1_59,ic_tag_valid_out_1_58,ic_tag_valid_out_1_57,ic_tag_valid_out_1_56,ic_tag_valid_out_1_55}; // @[Cat.scala 29:58]
  wire [81:0] _T_5595 = {_T_5586,ic_tag_valid_out_1_54,ic_tag_valid_out_1_53,ic_tag_valid_out_1_52,ic_tag_valid_out_1_51,ic_tag_valid_out_1_50,ic_tag_valid_out_1_49,ic_tag_valid_out_1_48,ic_tag_valid_out_1_47,ic_tag_valid_out_1_46}; // @[Cat.scala 29:58]
  wire [90:0] _T_5604 = {_T_5595,ic_tag_valid_out_1_45,ic_tag_valid_out_1_44,ic_tag_valid_out_1_43,ic_tag_valid_out_1_42,ic_tag_valid_out_1_41,ic_tag_valid_out_1_40,ic_tag_valid_out_1_39,ic_tag_valid_out_1_38,ic_tag_valid_out_1_37}; // @[Cat.scala 29:58]
  wire [99:0] _T_5613 = {_T_5604,ic_tag_valid_out_1_36,ic_tag_valid_out_1_35,ic_tag_valid_out_1_34,ic_tag_valid_out_1_33,ic_tag_valid_out_1_32,ic_tag_valid_out_1_31,ic_tag_valid_out_1_30,ic_tag_valid_out_1_29,ic_tag_valid_out_1_28}; // @[Cat.scala 29:58]
  wire [108:0] _T_5622 = {_T_5613,ic_tag_valid_out_1_27,ic_tag_valid_out_1_26,ic_tag_valid_out_1_25,ic_tag_valid_out_1_24,ic_tag_valid_out_1_23,ic_tag_valid_out_1_22,ic_tag_valid_out_1_21,ic_tag_valid_out_1_20,ic_tag_valid_out_1_19}; // @[Cat.scala 29:58]
  wire [117:0] _T_5631 = {_T_5622,ic_tag_valid_out_1_18,ic_tag_valid_out_1_17,ic_tag_valid_out_1_16,ic_tag_valid_out_1_15,ic_tag_valid_out_1_14,ic_tag_valid_out_1_13,ic_tag_valid_out_1_12,ic_tag_valid_out_1_11,ic_tag_valid_out_1_10}; // @[Cat.scala 29:58]
  wire [126:0] _T_5640 = {_T_5631,ic_tag_valid_out_1_9,ic_tag_valid_out_1_8,ic_tag_valid_out_1_7,ic_tag_valid_out_1_6,ic_tag_valid_out_1_5,ic_tag_valid_out_1_4,ic_tag_valid_out_1_3,ic_tag_valid_out_1_2,ic_tag_valid_out_1_1}; // @[Cat.scala 29:58]
  wire [127:0] _T_5641 = {_T_5640,ic_tag_valid_out_1_0}; // @[Cat.scala 29:58]
  wire [9:0] _T_5650 = {ic_tag_valid_out_0_127,ic_tag_valid_out_0_126,ic_tag_valid_out_0_125,ic_tag_valid_out_0_124,ic_tag_valid_out_0_123,ic_tag_valid_out_0_122,ic_tag_valid_out_0_121,ic_tag_valid_out_0_120,ic_tag_valid_out_0_119,ic_tag_valid_out_0_118}; // @[Cat.scala 29:58]
  wire [18:0] _T_5659 = {_T_5650,ic_tag_valid_out_0_117,ic_tag_valid_out_0_116,ic_tag_valid_out_0_115,ic_tag_valid_out_0_114,ic_tag_valid_out_0_113,ic_tag_valid_out_0_112,ic_tag_valid_out_0_111,ic_tag_valid_out_0_110,ic_tag_valid_out_0_109}; // @[Cat.scala 29:58]
  wire [27:0] _T_5668 = {_T_5659,ic_tag_valid_out_0_108,ic_tag_valid_out_0_107,ic_tag_valid_out_0_106,ic_tag_valid_out_0_105,ic_tag_valid_out_0_104,ic_tag_valid_out_0_103,ic_tag_valid_out_0_102,ic_tag_valid_out_0_101,ic_tag_valid_out_0_100}; // @[Cat.scala 29:58]
  wire [36:0] _T_5677 = {_T_5668,ic_tag_valid_out_0_99,ic_tag_valid_out_0_98,ic_tag_valid_out_0_97,ic_tag_valid_out_0_96,ic_tag_valid_out_0_95,ic_tag_valid_out_0_94,ic_tag_valid_out_0_93,ic_tag_valid_out_0_92,ic_tag_valid_out_0_91}; // @[Cat.scala 29:58]
  wire [45:0] _T_5686 = {_T_5677,ic_tag_valid_out_0_90,ic_tag_valid_out_0_89,ic_tag_valid_out_0_88,ic_tag_valid_out_0_87,ic_tag_valid_out_0_86,ic_tag_valid_out_0_85,ic_tag_valid_out_0_84,ic_tag_valid_out_0_83,ic_tag_valid_out_0_82}; // @[Cat.scala 29:58]
  wire [54:0] _T_5695 = {_T_5686,ic_tag_valid_out_0_81,ic_tag_valid_out_0_80,ic_tag_valid_out_0_79,ic_tag_valid_out_0_78,ic_tag_valid_out_0_77,ic_tag_valid_out_0_76,ic_tag_valid_out_0_75,ic_tag_valid_out_0_74,ic_tag_valid_out_0_73}; // @[Cat.scala 29:58]
  wire [63:0] _T_5704 = {_T_5695,ic_tag_valid_out_0_72,ic_tag_valid_out_0_71,ic_tag_valid_out_0_70,ic_tag_valid_out_0_69,ic_tag_valid_out_0_68,ic_tag_valid_out_0_67,ic_tag_valid_out_0_66,ic_tag_valid_out_0_65,ic_tag_valid_out_0_64}; // @[Cat.scala 29:58]
  wire [72:0] _T_5713 = {_T_5704,ic_tag_valid_out_0_63,ic_tag_valid_out_0_62,ic_tag_valid_out_0_61,ic_tag_valid_out_0_60,ic_tag_valid_out_0_59,ic_tag_valid_out_0_58,ic_tag_valid_out_0_57,ic_tag_valid_out_0_56,ic_tag_valid_out_0_55}; // @[Cat.scala 29:58]
  wire [81:0] _T_5722 = {_T_5713,ic_tag_valid_out_0_54,ic_tag_valid_out_0_53,ic_tag_valid_out_0_52,ic_tag_valid_out_0_51,ic_tag_valid_out_0_50,ic_tag_valid_out_0_49,ic_tag_valid_out_0_48,ic_tag_valid_out_0_47,ic_tag_valid_out_0_46}; // @[Cat.scala 29:58]
  wire [90:0] _T_5731 = {_T_5722,ic_tag_valid_out_0_45,ic_tag_valid_out_0_44,ic_tag_valid_out_0_43,ic_tag_valid_out_0_42,ic_tag_valid_out_0_41,ic_tag_valid_out_0_40,ic_tag_valid_out_0_39,ic_tag_valid_out_0_38,ic_tag_valid_out_0_37}; // @[Cat.scala 29:58]
  wire [99:0] _T_5740 = {_T_5731,ic_tag_valid_out_0_36,ic_tag_valid_out_0_35,ic_tag_valid_out_0_34,ic_tag_valid_out_0_33,ic_tag_valid_out_0_32,ic_tag_valid_out_0_31,ic_tag_valid_out_0_30,ic_tag_valid_out_0_29,ic_tag_valid_out_0_28}; // @[Cat.scala 29:58]
  wire [108:0] _T_5749 = {_T_5740,ic_tag_valid_out_0_27,ic_tag_valid_out_0_26,ic_tag_valid_out_0_25,ic_tag_valid_out_0_24,ic_tag_valid_out_0_23,ic_tag_valid_out_0_22,ic_tag_valid_out_0_21,ic_tag_valid_out_0_20,ic_tag_valid_out_0_19}; // @[Cat.scala 29:58]
  wire [117:0] _T_5758 = {_T_5749,ic_tag_valid_out_0_18,ic_tag_valid_out_0_17,ic_tag_valid_out_0_16,ic_tag_valid_out_0_15,ic_tag_valid_out_0_14,ic_tag_valid_out_0_13,ic_tag_valid_out_0_12,ic_tag_valid_out_0_11,ic_tag_valid_out_0_10}; // @[Cat.scala 29:58]
  wire [126:0] _T_5767 = {_T_5758,ic_tag_valid_out_0_9,ic_tag_valid_out_0_8,ic_tag_valid_out_0_7,ic_tag_valid_out_0_6,ic_tag_valid_out_0_5,ic_tag_valid_out_0_4,ic_tag_valid_out_0_3,ic_tag_valid_out_0_2,ic_tag_valid_out_0_1}; // @[Cat.scala 29:58]
  wire [127:0] _T_5768 = {_T_5767,ic_tag_valid_out_0_0}; // @[Cat.scala 29:58]
  wire  _T_5772 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 760:66]
  wire  _T_5773 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 760:93]
  wire  _T_5774 = _T_5772 & _T_5773; // @[el2_ifu_mem_ctl.scala 760:91]
  wire  _T_5777 = _T_4789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5778 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5780 = _T_5778 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5781 = _T_5777 | _T_5780; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5782 = _T_5781 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5784 = _T_5782 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5794 = _T_4793 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5795 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5797 = _T_5795 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5798 = _T_5794 | _T_5797; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5799 = _T_5798 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5801 = _T_5799 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5811 = _T_4797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5812 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5814 = _T_5812 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5815 = _T_5811 | _T_5814; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5816 = _T_5815 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5818 = _T_5816 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5828 = _T_4801 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5829 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5831 = _T_5829 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5832 = _T_5828 | _T_5831; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5833 = _T_5832 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5835 = _T_5833 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5845 = _T_4805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5846 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5848 = _T_5846 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5849 = _T_5845 | _T_5848; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5850 = _T_5849 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5852 = _T_5850 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5862 = _T_4809 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5863 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5865 = _T_5863 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5866 = _T_5862 | _T_5865; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5867 = _T_5866 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5869 = _T_5867 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5879 = _T_4813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5880 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5882 = _T_5880 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5883 = _T_5879 | _T_5882; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5884 = _T_5883 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5886 = _T_5884 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5896 = _T_4817 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5897 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5899 = _T_5897 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5900 = _T_5896 | _T_5899; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5901 = _T_5900 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5903 = _T_5901 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5913 = _T_4821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5914 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5916 = _T_5914 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5917 = _T_5913 | _T_5916; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5918 = _T_5917 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5920 = _T_5918 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5930 = _T_4825 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5931 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5933 = _T_5931 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5934 = _T_5930 | _T_5933; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5935 = _T_5934 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5937 = _T_5935 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5947 = _T_4829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5948 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5950 = _T_5948 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5951 = _T_5947 | _T_5950; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5952 = _T_5951 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5954 = _T_5952 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5964 = _T_4833 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5965 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5967 = _T_5965 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5968 = _T_5964 | _T_5967; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5969 = _T_5968 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5971 = _T_5969 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5981 = _T_4837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5982 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_5984 = _T_5982 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_5985 = _T_5981 | _T_5984; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_5986 = _T_5985 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_5988 = _T_5986 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_5998 = _T_4841 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_5999 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6001 = _T_5999 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6002 = _T_5998 | _T_6001; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6003 = _T_6002 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6005 = _T_6003 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6015 = _T_4845 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6016 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6018 = _T_6016 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6019 = _T_6015 | _T_6018; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6020 = _T_6019 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6022 = _T_6020 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6032 = _T_4849 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6033 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6035 = _T_6033 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6036 = _T_6032 | _T_6035; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6037 = _T_6036 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6039 = _T_6037 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6049 = _T_4853 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6050 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6052 = _T_6050 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6053 = _T_6049 | _T_6052; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6054 = _T_6053 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6056 = _T_6054 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6066 = _T_4857 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6067 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6069 = _T_6067 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6070 = _T_6066 | _T_6069; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6071 = _T_6070 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6073 = _T_6071 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6083 = _T_4861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6084 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6086 = _T_6084 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6087 = _T_6083 | _T_6086; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6088 = _T_6087 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6090 = _T_6088 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6100 = _T_4865 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6101 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6103 = _T_6101 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6104 = _T_6100 | _T_6103; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6105 = _T_6104 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6107 = _T_6105 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6117 = _T_4869 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6118 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6120 = _T_6118 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6121 = _T_6117 | _T_6120; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6122 = _T_6121 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6124 = _T_6122 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6134 = _T_4873 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6135 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6137 = _T_6135 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6138 = _T_6134 | _T_6137; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6139 = _T_6138 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6141 = _T_6139 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6151 = _T_4877 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6152 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6154 = _T_6152 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6155 = _T_6151 | _T_6154; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6156 = _T_6155 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6158 = _T_6156 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6168 = _T_4881 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6169 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6171 = _T_6169 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6172 = _T_6168 | _T_6171; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6173 = _T_6172 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6175 = _T_6173 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6185 = _T_4885 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6186 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6188 = _T_6186 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6189 = _T_6185 | _T_6188; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6190 = _T_6189 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6192 = _T_6190 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6202 = _T_4889 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6203 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6205 = _T_6203 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6206 = _T_6202 | _T_6205; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6207 = _T_6206 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6209 = _T_6207 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6219 = _T_4893 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6220 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6222 = _T_6220 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6223 = _T_6219 | _T_6222; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6224 = _T_6223 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6226 = _T_6224 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6236 = _T_4897 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6237 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6239 = _T_6237 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6240 = _T_6236 | _T_6239; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6241 = _T_6240 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6243 = _T_6241 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6253 = _T_4901 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6254 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6256 = _T_6254 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6257 = _T_6253 | _T_6256; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6258 = _T_6257 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6260 = _T_6258 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6270 = _T_4905 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6271 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6273 = _T_6271 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6274 = _T_6270 | _T_6273; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6275 = _T_6274 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6277 = _T_6275 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6287 = _T_4909 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6288 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6290 = _T_6288 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6291 = _T_6287 | _T_6290; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6292 = _T_6291 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6294 = _T_6292 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6304 = _T_4913 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6305 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6307 = _T_6305 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6308 = _T_6304 | _T_6307; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6309 = _T_6308 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6311 = _T_6309 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6321 = _T_4789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6324 = _T_5778 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6325 = _T_6321 | _T_6324; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6326 = _T_6325 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6328 = _T_6326 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6338 = _T_4793 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6341 = _T_5795 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6342 = _T_6338 | _T_6341; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6343 = _T_6342 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6345 = _T_6343 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6355 = _T_4797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6358 = _T_5812 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6359 = _T_6355 | _T_6358; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6360 = _T_6359 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6362 = _T_6360 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6372 = _T_4801 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6375 = _T_5829 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6376 = _T_6372 | _T_6375; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6377 = _T_6376 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6379 = _T_6377 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6389 = _T_4805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6392 = _T_5846 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6393 = _T_6389 | _T_6392; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6394 = _T_6393 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6396 = _T_6394 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6406 = _T_4809 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6409 = _T_5863 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6410 = _T_6406 | _T_6409; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6411 = _T_6410 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6413 = _T_6411 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6423 = _T_4813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6426 = _T_5880 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6427 = _T_6423 | _T_6426; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6428 = _T_6427 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6430 = _T_6428 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6440 = _T_4817 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6443 = _T_5897 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6444 = _T_6440 | _T_6443; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6445 = _T_6444 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6447 = _T_6445 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6457 = _T_4821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6460 = _T_5914 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6461 = _T_6457 | _T_6460; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6462 = _T_6461 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6464 = _T_6462 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6474 = _T_4825 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6477 = _T_5931 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6478 = _T_6474 | _T_6477; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6479 = _T_6478 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6481 = _T_6479 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6491 = _T_4829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6494 = _T_5948 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6495 = _T_6491 | _T_6494; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6496 = _T_6495 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6498 = _T_6496 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6508 = _T_4833 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6511 = _T_5965 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6512 = _T_6508 | _T_6511; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6513 = _T_6512 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6515 = _T_6513 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6525 = _T_4837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6528 = _T_5982 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6529 = _T_6525 | _T_6528; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6530 = _T_6529 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6532 = _T_6530 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6542 = _T_4841 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6545 = _T_5999 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6546 = _T_6542 | _T_6545; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6547 = _T_6546 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6549 = _T_6547 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6559 = _T_4845 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6562 = _T_6016 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6563 = _T_6559 | _T_6562; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6564 = _T_6563 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6566 = _T_6564 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6576 = _T_4849 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6579 = _T_6033 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6580 = _T_6576 | _T_6579; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6581 = _T_6580 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6583 = _T_6581 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6593 = _T_4853 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6596 = _T_6050 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6597 = _T_6593 | _T_6596; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6598 = _T_6597 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6600 = _T_6598 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6610 = _T_4857 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6613 = _T_6067 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6614 = _T_6610 | _T_6613; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6615 = _T_6614 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6617 = _T_6615 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6627 = _T_4861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6630 = _T_6084 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6631 = _T_6627 | _T_6630; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6632 = _T_6631 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6634 = _T_6632 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6644 = _T_4865 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6647 = _T_6101 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6648 = _T_6644 | _T_6647; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6649 = _T_6648 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6651 = _T_6649 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6661 = _T_4869 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6664 = _T_6118 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6665 = _T_6661 | _T_6664; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6666 = _T_6665 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6668 = _T_6666 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6678 = _T_4873 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6681 = _T_6135 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6682 = _T_6678 | _T_6681; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6683 = _T_6682 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6685 = _T_6683 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6695 = _T_4877 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6698 = _T_6152 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6699 = _T_6695 | _T_6698; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6700 = _T_6699 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6702 = _T_6700 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6712 = _T_4881 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6715 = _T_6169 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6716 = _T_6712 | _T_6715; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6717 = _T_6716 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6719 = _T_6717 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6729 = _T_4885 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6732 = _T_6186 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6733 = _T_6729 | _T_6732; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6734 = _T_6733 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6736 = _T_6734 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6746 = _T_4889 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6749 = _T_6203 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6750 = _T_6746 | _T_6749; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6751 = _T_6750 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6753 = _T_6751 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6763 = _T_4893 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6766 = _T_6220 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6767 = _T_6763 | _T_6766; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6768 = _T_6767 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6770 = _T_6768 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6780 = _T_4897 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6783 = _T_6237 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6784 = _T_6780 | _T_6783; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6785 = _T_6784 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6787 = _T_6785 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6797 = _T_4901 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6800 = _T_6254 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6801 = _T_6797 | _T_6800; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6802 = _T_6801 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6804 = _T_6802 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6814 = _T_4905 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6817 = _T_6271 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6818 = _T_6814 | _T_6817; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6819 = _T_6818 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6821 = _T_6819 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6831 = _T_4909 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6834 = _T_6288 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6835 = _T_6831 | _T_6834; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6836 = _T_6835 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6838 = _T_6836 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6848 = _T_4913 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6851 = _T_6305 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6852 = _T_6848 | _T_6851; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6853 = _T_6852 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6855 = _T_6853 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6865 = _T_4917 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6866 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6868 = _T_6866 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6869 = _T_6865 | _T_6868; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6870 = _T_6869 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6872 = _T_6870 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6882 = _T_4921 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6883 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6885 = _T_6883 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6886 = _T_6882 | _T_6885; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6887 = _T_6886 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6889 = _T_6887 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6899 = _T_4925 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6900 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6902 = _T_6900 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6903 = _T_6899 | _T_6902; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6904 = _T_6903 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6906 = _T_6904 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6916 = _T_4929 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6917 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6919 = _T_6917 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6920 = _T_6916 | _T_6919; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6921 = _T_6920 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6923 = _T_6921 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6933 = _T_4933 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6934 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6936 = _T_6934 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6937 = _T_6933 | _T_6936; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6938 = _T_6937 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6940 = _T_6938 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6950 = _T_4937 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6951 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6953 = _T_6951 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6954 = _T_6950 | _T_6953; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6955 = _T_6954 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6957 = _T_6955 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6967 = _T_4941 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6968 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6970 = _T_6968 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6971 = _T_6967 | _T_6970; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6972 = _T_6971 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6974 = _T_6972 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_6984 = _T_4945 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_6985 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_6987 = _T_6985 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_6988 = _T_6984 | _T_6987; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_6989 = _T_6988 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_6991 = _T_6989 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7001 = _T_4949 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7002 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7004 = _T_7002 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7005 = _T_7001 | _T_7004; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7006 = _T_7005 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7008 = _T_7006 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7018 = _T_4953 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7019 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7021 = _T_7019 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7022 = _T_7018 | _T_7021; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7023 = _T_7022 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7025 = _T_7023 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7035 = _T_4957 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7036 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7038 = _T_7036 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7039 = _T_7035 | _T_7038; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7040 = _T_7039 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7042 = _T_7040 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7052 = _T_4961 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7053 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7055 = _T_7053 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7056 = _T_7052 | _T_7055; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7057 = _T_7056 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7059 = _T_7057 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7069 = _T_4965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7070 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7072 = _T_7070 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7073 = _T_7069 | _T_7072; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7074 = _T_7073 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7076 = _T_7074 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7086 = _T_4969 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7087 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7089 = _T_7087 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7090 = _T_7086 | _T_7089; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7091 = _T_7090 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7093 = _T_7091 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7103 = _T_4973 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7104 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7106 = _T_7104 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7107 = _T_7103 | _T_7106; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7108 = _T_7107 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7110 = _T_7108 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7120 = _T_4977 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7121 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7123 = _T_7121 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7124 = _T_7120 | _T_7123; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7125 = _T_7124 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7127 = _T_7125 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7137 = _T_4981 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7138 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7140 = _T_7138 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7141 = _T_7137 | _T_7140; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7142 = _T_7141 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7144 = _T_7142 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7154 = _T_4985 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7155 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7157 = _T_7155 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7158 = _T_7154 | _T_7157; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7159 = _T_7158 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7161 = _T_7159 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7171 = _T_4989 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7172 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7174 = _T_7172 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7175 = _T_7171 | _T_7174; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7176 = _T_7175 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7178 = _T_7176 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7188 = _T_4993 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7189 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7191 = _T_7189 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7192 = _T_7188 | _T_7191; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7193 = _T_7192 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7195 = _T_7193 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7205 = _T_4997 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7206 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7208 = _T_7206 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7209 = _T_7205 | _T_7208; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7210 = _T_7209 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7212 = _T_7210 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7222 = _T_5001 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7223 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7225 = _T_7223 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7226 = _T_7222 | _T_7225; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7227 = _T_7226 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7229 = _T_7227 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7239 = _T_5005 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7240 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7242 = _T_7240 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7243 = _T_7239 | _T_7242; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7244 = _T_7243 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7246 = _T_7244 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7256 = _T_5009 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7257 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7259 = _T_7257 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7260 = _T_7256 | _T_7259; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7261 = _T_7260 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7263 = _T_7261 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7273 = _T_5013 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7274 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7276 = _T_7274 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7277 = _T_7273 | _T_7276; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7278 = _T_7277 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7280 = _T_7278 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7290 = _T_5017 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7291 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7293 = _T_7291 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7294 = _T_7290 | _T_7293; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7295 = _T_7294 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7297 = _T_7295 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7307 = _T_5021 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7308 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7310 = _T_7308 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7311 = _T_7307 | _T_7310; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7312 = _T_7311 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7314 = _T_7312 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7324 = _T_5025 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7325 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7327 = _T_7325 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7328 = _T_7324 | _T_7327; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7329 = _T_7328 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7331 = _T_7329 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7341 = _T_5029 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7342 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7344 = _T_7342 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7345 = _T_7341 | _T_7344; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7346 = _T_7345 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7348 = _T_7346 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7358 = _T_5033 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7359 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7361 = _T_7359 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7362 = _T_7358 | _T_7361; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7363 = _T_7362 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7365 = _T_7363 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7375 = _T_5037 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7376 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7378 = _T_7376 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7379 = _T_7375 | _T_7378; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7380 = _T_7379 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7382 = _T_7380 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7392 = _T_5041 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7393 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7395 = _T_7393 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7396 = _T_7392 | _T_7395; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7397 = _T_7396 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7399 = _T_7397 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7409 = _T_4917 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7412 = _T_6866 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7413 = _T_7409 | _T_7412; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7414 = _T_7413 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7416 = _T_7414 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7426 = _T_4921 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7429 = _T_6883 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7430 = _T_7426 | _T_7429; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7431 = _T_7430 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7433 = _T_7431 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7443 = _T_4925 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7446 = _T_6900 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7447 = _T_7443 | _T_7446; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7448 = _T_7447 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7450 = _T_7448 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7460 = _T_4929 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7463 = _T_6917 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7464 = _T_7460 | _T_7463; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7465 = _T_7464 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7467 = _T_7465 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7477 = _T_4933 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7480 = _T_6934 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7481 = _T_7477 | _T_7480; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7482 = _T_7481 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7484 = _T_7482 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7494 = _T_4937 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7497 = _T_6951 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7498 = _T_7494 | _T_7497; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7499 = _T_7498 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7501 = _T_7499 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7511 = _T_4941 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7514 = _T_6968 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7515 = _T_7511 | _T_7514; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7516 = _T_7515 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7518 = _T_7516 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7528 = _T_4945 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7531 = _T_6985 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7532 = _T_7528 | _T_7531; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7533 = _T_7532 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7535 = _T_7533 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7545 = _T_4949 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7548 = _T_7002 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7549 = _T_7545 | _T_7548; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7550 = _T_7549 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7552 = _T_7550 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7562 = _T_4953 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7565 = _T_7019 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7566 = _T_7562 | _T_7565; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7567 = _T_7566 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7569 = _T_7567 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7579 = _T_4957 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7582 = _T_7036 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7583 = _T_7579 | _T_7582; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7584 = _T_7583 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7586 = _T_7584 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7596 = _T_4961 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7599 = _T_7053 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7600 = _T_7596 | _T_7599; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7601 = _T_7600 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7603 = _T_7601 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7613 = _T_4965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7616 = _T_7070 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7617 = _T_7613 | _T_7616; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7618 = _T_7617 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7620 = _T_7618 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7630 = _T_4969 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7633 = _T_7087 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7634 = _T_7630 | _T_7633; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7635 = _T_7634 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7637 = _T_7635 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7647 = _T_4973 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7650 = _T_7104 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7651 = _T_7647 | _T_7650; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7652 = _T_7651 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7654 = _T_7652 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7664 = _T_4977 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7667 = _T_7121 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7668 = _T_7664 | _T_7667; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7669 = _T_7668 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7671 = _T_7669 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7681 = _T_4981 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7684 = _T_7138 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7685 = _T_7681 | _T_7684; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7686 = _T_7685 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7688 = _T_7686 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7698 = _T_4985 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7701 = _T_7155 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7702 = _T_7698 | _T_7701; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7703 = _T_7702 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7705 = _T_7703 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7715 = _T_4989 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7718 = _T_7172 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7719 = _T_7715 | _T_7718; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7720 = _T_7719 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7722 = _T_7720 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7732 = _T_4993 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7735 = _T_7189 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7736 = _T_7732 | _T_7735; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7737 = _T_7736 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7739 = _T_7737 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7749 = _T_4997 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7752 = _T_7206 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7753 = _T_7749 | _T_7752; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7754 = _T_7753 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7756 = _T_7754 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7766 = _T_5001 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7769 = _T_7223 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7770 = _T_7766 | _T_7769; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7771 = _T_7770 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7773 = _T_7771 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7783 = _T_5005 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7786 = _T_7240 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7787 = _T_7783 | _T_7786; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7788 = _T_7787 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7790 = _T_7788 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7800 = _T_5009 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7803 = _T_7257 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7804 = _T_7800 | _T_7803; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7805 = _T_7804 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7807 = _T_7805 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7817 = _T_5013 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7820 = _T_7274 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7821 = _T_7817 | _T_7820; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7822 = _T_7821 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7824 = _T_7822 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7834 = _T_5017 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7837 = _T_7291 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7838 = _T_7834 | _T_7837; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7839 = _T_7838 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7841 = _T_7839 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7851 = _T_5021 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7854 = _T_7308 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7855 = _T_7851 | _T_7854; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7856 = _T_7855 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7858 = _T_7856 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7868 = _T_5025 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7871 = _T_7325 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7872 = _T_7868 | _T_7871; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7873 = _T_7872 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7875 = _T_7873 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7885 = _T_5029 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7888 = _T_7342 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7889 = _T_7885 | _T_7888; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7890 = _T_7889 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7892 = _T_7890 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7902 = _T_5033 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7905 = _T_7359 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7906 = _T_7902 | _T_7905; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7907 = _T_7906 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7909 = _T_7907 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7919 = _T_5037 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7922 = _T_7376 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7923 = _T_7919 | _T_7922; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7924 = _T_7923 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7926 = _T_7924 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7936 = _T_5041 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7939 = _T_7393 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7940 = _T_7936 | _T_7939; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7941 = _T_7940 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7943 = _T_7941 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7953 = _T_5045 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7954 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7956 = _T_7954 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7957 = _T_7953 | _T_7956; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7958 = _T_7957 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7960 = _T_7958 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7970 = _T_5049 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7971 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7973 = _T_7971 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7974 = _T_7970 | _T_7973; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7975 = _T_7974 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7977 = _T_7975 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_7987 = _T_5053 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_7988 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_7990 = _T_7988 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_7991 = _T_7987 | _T_7990; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_7992 = _T_7991 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_7994 = _T_7992 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8004 = _T_5057 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8005 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8007 = _T_8005 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8008 = _T_8004 | _T_8007; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8009 = _T_8008 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8011 = _T_8009 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8021 = _T_5061 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8022 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8024 = _T_8022 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8025 = _T_8021 | _T_8024; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8026 = _T_8025 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8028 = _T_8026 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8038 = _T_5065 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8039 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8041 = _T_8039 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8042 = _T_8038 | _T_8041; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8043 = _T_8042 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8045 = _T_8043 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8055 = _T_5069 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8056 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8058 = _T_8056 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8059 = _T_8055 | _T_8058; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8060 = _T_8059 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8062 = _T_8060 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8072 = _T_5073 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8073 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8075 = _T_8073 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8076 = _T_8072 | _T_8075; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8077 = _T_8076 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8079 = _T_8077 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8089 = _T_5077 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8090 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8092 = _T_8090 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8093 = _T_8089 | _T_8092; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8094 = _T_8093 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8096 = _T_8094 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8106 = _T_5081 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8107 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8109 = _T_8107 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8110 = _T_8106 | _T_8109; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8111 = _T_8110 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8113 = _T_8111 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8123 = _T_5085 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8124 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8126 = _T_8124 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8127 = _T_8123 | _T_8126; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8128 = _T_8127 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8130 = _T_8128 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8140 = _T_5089 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8141 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8143 = _T_8141 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8144 = _T_8140 | _T_8143; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8145 = _T_8144 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8147 = _T_8145 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8157 = _T_5093 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8158 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8160 = _T_8158 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8161 = _T_8157 | _T_8160; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8162 = _T_8161 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8164 = _T_8162 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8174 = _T_5097 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8175 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8177 = _T_8175 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8178 = _T_8174 | _T_8177; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8179 = _T_8178 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8181 = _T_8179 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8191 = _T_5101 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8192 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8194 = _T_8192 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8195 = _T_8191 | _T_8194; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8196 = _T_8195 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8198 = _T_8196 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8208 = _T_5105 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8209 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8211 = _T_8209 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8212 = _T_8208 | _T_8211; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8213 = _T_8212 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8215 = _T_8213 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8225 = _T_5109 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8226 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8228 = _T_8226 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8229 = _T_8225 | _T_8228; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8230 = _T_8229 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8232 = _T_8230 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8242 = _T_5113 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8243 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8245 = _T_8243 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8246 = _T_8242 | _T_8245; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8247 = _T_8246 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8249 = _T_8247 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8259 = _T_5117 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8260 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8262 = _T_8260 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8263 = _T_8259 | _T_8262; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8264 = _T_8263 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8266 = _T_8264 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8276 = _T_5121 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8277 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8279 = _T_8277 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8280 = _T_8276 | _T_8279; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8281 = _T_8280 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8283 = _T_8281 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8293 = _T_5125 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8294 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8296 = _T_8294 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8297 = _T_8293 | _T_8296; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8298 = _T_8297 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8300 = _T_8298 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8310 = _T_5129 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8311 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8313 = _T_8311 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8314 = _T_8310 | _T_8313; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8315 = _T_8314 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8317 = _T_8315 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8327 = _T_5133 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8328 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8330 = _T_8328 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8331 = _T_8327 | _T_8330; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8332 = _T_8331 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8334 = _T_8332 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8344 = _T_5137 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8345 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8347 = _T_8345 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8348 = _T_8344 | _T_8347; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8349 = _T_8348 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8351 = _T_8349 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8361 = _T_5141 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8362 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8364 = _T_8362 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8365 = _T_8361 | _T_8364; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8366 = _T_8365 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8368 = _T_8366 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8378 = _T_5145 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8379 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8381 = _T_8379 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8382 = _T_8378 | _T_8381; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8383 = _T_8382 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8385 = _T_8383 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8395 = _T_5149 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8396 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8398 = _T_8396 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8399 = _T_8395 | _T_8398; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8400 = _T_8399 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8402 = _T_8400 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8412 = _T_5153 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8413 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8415 = _T_8413 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8416 = _T_8412 | _T_8415; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8417 = _T_8416 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8419 = _T_8417 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8429 = _T_5157 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8430 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8432 = _T_8430 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8433 = _T_8429 | _T_8432; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8434 = _T_8433 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8436 = _T_8434 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8446 = _T_5161 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8447 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8449 = _T_8447 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8450 = _T_8446 | _T_8449; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8451 = _T_8450 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8453 = _T_8451 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8463 = _T_5165 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8464 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8466 = _T_8464 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8467 = _T_8463 | _T_8466; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8468 = _T_8467 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8470 = _T_8468 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8480 = _T_5169 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8481 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_8483 = _T_8481 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8484 = _T_8480 | _T_8483; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8485 = _T_8484 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8487 = _T_8485 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8497 = _T_5045 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8500 = _T_7954 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8501 = _T_8497 | _T_8500; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8502 = _T_8501 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8504 = _T_8502 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8514 = _T_5049 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8517 = _T_7971 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8518 = _T_8514 | _T_8517; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8519 = _T_8518 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8521 = _T_8519 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8531 = _T_5053 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8534 = _T_7988 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8535 = _T_8531 | _T_8534; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8536 = _T_8535 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8538 = _T_8536 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8548 = _T_5057 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8551 = _T_8005 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8552 = _T_8548 | _T_8551; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8553 = _T_8552 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8555 = _T_8553 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8565 = _T_5061 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8568 = _T_8022 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8569 = _T_8565 | _T_8568; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8570 = _T_8569 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8572 = _T_8570 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8582 = _T_5065 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8585 = _T_8039 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8586 = _T_8582 | _T_8585; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8587 = _T_8586 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8589 = _T_8587 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8599 = _T_5069 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8602 = _T_8056 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8603 = _T_8599 | _T_8602; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8604 = _T_8603 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8606 = _T_8604 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8616 = _T_5073 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8619 = _T_8073 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8620 = _T_8616 | _T_8619; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8621 = _T_8620 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8623 = _T_8621 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8633 = _T_5077 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8636 = _T_8090 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8637 = _T_8633 | _T_8636; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8638 = _T_8637 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8640 = _T_8638 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8650 = _T_5081 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8653 = _T_8107 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8654 = _T_8650 | _T_8653; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8655 = _T_8654 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8657 = _T_8655 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8667 = _T_5085 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8670 = _T_8124 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8671 = _T_8667 | _T_8670; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8672 = _T_8671 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8674 = _T_8672 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8684 = _T_5089 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8687 = _T_8141 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8688 = _T_8684 | _T_8687; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8689 = _T_8688 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8691 = _T_8689 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8701 = _T_5093 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8704 = _T_8158 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8705 = _T_8701 | _T_8704; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8706 = _T_8705 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8708 = _T_8706 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8718 = _T_5097 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8721 = _T_8175 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8722 = _T_8718 | _T_8721; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8723 = _T_8722 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8725 = _T_8723 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8735 = _T_5101 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8738 = _T_8192 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8739 = _T_8735 | _T_8738; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8740 = _T_8739 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8742 = _T_8740 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8752 = _T_5105 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8755 = _T_8209 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8756 = _T_8752 | _T_8755; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8757 = _T_8756 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8759 = _T_8757 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8769 = _T_5109 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8772 = _T_8226 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8773 = _T_8769 | _T_8772; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8774 = _T_8773 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8776 = _T_8774 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8786 = _T_5113 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8789 = _T_8243 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8790 = _T_8786 | _T_8789; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8791 = _T_8790 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8793 = _T_8791 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8803 = _T_5117 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8806 = _T_8260 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8807 = _T_8803 | _T_8806; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8808 = _T_8807 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8810 = _T_8808 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8820 = _T_5121 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8823 = _T_8277 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8824 = _T_8820 | _T_8823; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8825 = _T_8824 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8827 = _T_8825 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8837 = _T_5125 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8840 = _T_8294 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8841 = _T_8837 | _T_8840; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8842 = _T_8841 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8844 = _T_8842 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8854 = _T_5129 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8857 = _T_8311 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8858 = _T_8854 | _T_8857; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8859 = _T_8858 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8861 = _T_8859 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8871 = _T_5133 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8874 = _T_8328 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8875 = _T_8871 | _T_8874; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8876 = _T_8875 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8878 = _T_8876 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8888 = _T_5137 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8891 = _T_8345 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8892 = _T_8888 | _T_8891; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8893 = _T_8892 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8895 = _T_8893 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8905 = _T_5141 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8908 = _T_8362 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8909 = _T_8905 | _T_8908; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8910 = _T_8909 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8912 = _T_8910 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8922 = _T_5145 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8925 = _T_8379 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8926 = _T_8922 | _T_8925; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8927 = _T_8926 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8929 = _T_8927 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8939 = _T_5149 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8942 = _T_8396 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8943 = _T_8939 | _T_8942; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8944 = _T_8943 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8946 = _T_8944 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8956 = _T_5153 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8959 = _T_8413 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8960 = _T_8956 | _T_8959; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8961 = _T_8960 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8963 = _T_8961 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8973 = _T_5157 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8976 = _T_8430 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8977 = _T_8973 | _T_8976; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8978 = _T_8977 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8980 = _T_8978 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_8990 = _T_5161 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_8993 = _T_8447 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_8994 = _T_8990 | _T_8993; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_8995 = _T_8994 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_8997 = _T_8995 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9007 = _T_5165 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9010 = _T_8464 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9011 = _T_9007 | _T_9010; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9012 = _T_9011 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9014 = _T_9012 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9024 = _T_5169 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9027 = _T_8481 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9028 = _T_9024 | _T_9027; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9029 = _T_9028 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9031 = _T_9029 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9041 = _T_5173 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9042 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9044 = _T_9042 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9045 = _T_9041 | _T_9044; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9046 = _T_9045 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9048 = _T_9046 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9058 = _T_5177 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9059 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9061 = _T_9059 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9062 = _T_9058 | _T_9061; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9063 = _T_9062 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9065 = _T_9063 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9075 = _T_5181 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9076 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9078 = _T_9076 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9079 = _T_9075 | _T_9078; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9080 = _T_9079 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9082 = _T_9080 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9092 = _T_5185 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9093 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9095 = _T_9093 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9096 = _T_9092 | _T_9095; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9097 = _T_9096 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9099 = _T_9097 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9109 = _T_5189 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9110 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9112 = _T_9110 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9113 = _T_9109 | _T_9112; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9114 = _T_9113 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9116 = _T_9114 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9126 = _T_5193 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9127 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9129 = _T_9127 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9130 = _T_9126 | _T_9129; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9131 = _T_9130 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9133 = _T_9131 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9143 = _T_5197 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9144 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9146 = _T_9144 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9147 = _T_9143 | _T_9146; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9148 = _T_9147 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9150 = _T_9148 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9160 = _T_5201 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9161 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9163 = _T_9161 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9164 = _T_9160 | _T_9163; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9165 = _T_9164 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9167 = _T_9165 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9177 = _T_5205 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9178 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9180 = _T_9178 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9181 = _T_9177 | _T_9180; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9182 = _T_9181 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9184 = _T_9182 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9194 = _T_5209 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9195 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9197 = _T_9195 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9198 = _T_9194 | _T_9197; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9199 = _T_9198 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9201 = _T_9199 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9211 = _T_5213 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9212 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9214 = _T_9212 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9215 = _T_9211 | _T_9214; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9216 = _T_9215 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9218 = _T_9216 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9228 = _T_5217 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9229 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9231 = _T_9229 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9232 = _T_9228 | _T_9231; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9233 = _T_9232 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9235 = _T_9233 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9245 = _T_5221 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9246 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9248 = _T_9246 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9249 = _T_9245 | _T_9248; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9250 = _T_9249 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9252 = _T_9250 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9262 = _T_5225 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9263 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9265 = _T_9263 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9266 = _T_9262 | _T_9265; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9267 = _T_9266 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9269 = _T_9267 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9279 = _T_5229 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9280 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9282 = _T_9280 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9283 = _T_9279 | _T_9282; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9284 = _T_9283 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9286 = _T_9284 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9296 = _T_5233 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9297 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9299 = _T_9297 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9300 = _T_9296 | _T_9299; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9301 = _T_9300 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9303 = _T_9301 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9313 = _T_5237 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9314 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9316 = _T_9314 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9317 = _T_9313 | _T_9316; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9318 = _T_9317 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9320 = _T_9318 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9330 = _T_5241 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9331 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9333 = _T_9331 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9334 = _T_9330 | _T_9333; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9335 = _T_9334 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9337 = _T_9335 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9347 = _T_5245 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9348 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9350 = _T_9348 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9351 = _T_9347 | _T_9350; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9352 = _T_9351 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9354 = _T_9352 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9364 = _T_5249 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9365 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9367 = _T_9365 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9368 = _T_9364 | _T_9367; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9369 = _T_9368 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9371 = _T_9369 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9381 = _T_5253 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9382 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9384 = _T_9382 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9385 = _T_9381 | _T_9384; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9386 = _T_9385 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9388 = _T_9386 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9398 = _T_5257 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9399 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9401 = _T_9399 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9402 = _T_9398 | _T_9401; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9403 = _T_9402 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9405 = _T_9403 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9415 = _T_5261 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9416 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9418 = _T_9416 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9419 = _T_9415 | _T_9418; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9420 = _T_9419 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9422 = _T_9420 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9432 = _T_5265 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9433 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9435 = _T_9433 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9436 = _T_9432 | _T_9435; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9437 = _T_9436 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9439 = _T_9437 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9449 = _T_5269 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9450 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9452 = _T_9450 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9453 = _T_9449 | _T_9452; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9454 = _T_9453 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9456 = _T_9454 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9466 = _T_5273 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9467 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9469 = _T_9467 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9470 = _T_9466 | _T_9469; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9471 = _T_9470 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9473 = _T_9471 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9483 = _T_5277 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9484 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9486 = _T_9484 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9487 = _T_9483 | _T_9486; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9488 = _T_9487 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9490 = _T_9488 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9500 = _T_5281 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9501 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9503 = _T_9501 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9504 = _T_9500 | _T_9503; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9505 = _T_9504 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9507 = _T_9505 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9517 = _T_5285 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9518 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9520 = _T_9518 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9521 = _T_9517 | _T_9520; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9522 = _T_9521 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9524 = _T_9522 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9534 = _T_5289 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9535 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9537 = _T_9535 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9538 = _T_9534 | _T_9537; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9539 = _T_9538 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9541 = _T_9539 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9551 = _T_5293 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9552 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9554 = _T_9552 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9555 = _T_9551 | _T_9554; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9556 = _T_9555 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9558 = _T_9556 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9568 = _T_5297 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9569 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 761:102]
  wire  _T_9571 = _T_9569 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9572 = _T_9568 | _T_9571; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9573 = _T_9572 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9575 = _T_9573 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9585 = _T_5173 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9588 = _T_9042 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9589 = _T_9585 | _T_9588; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9590 = _T_9589 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9592 = _T_9590 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9602 = _T_5177 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9605 = _T_9059 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9606 = _T_9602 | _T_9605; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9607 = _T_9606 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9609 = _T_9607 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9619 = _T_5181 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9622 = _T_9076 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9623 = _T_9619 | _T_9622; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9624 = _T_9623 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9626 = _T_9624 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9636 = _T_5185 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9639 = _T_9093 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9640 = _T_9636 | _T_9639; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9641 = _T_9640 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9643 = _T_9641 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9653 = _T_5189 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9656 = _T_9110 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9657 = _T_9653 | _T_9656; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9658 = _T_9657 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9660 = _T_9658 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9670 = _T_5193 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9673 = _T_9127 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9674 = _T_9670 | _T_9673; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9675 = _T_9674 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9677 = _T_9675 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9687 = _T_5197 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9690 = _T_9144 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9691 = _T_9687 | _T_9690; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9692 = _T_9691 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9694 = _T_9692 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9704 = _T_5201 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9707 = _T_9161 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9708 = _T_9704 | _T_9707; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9709 = _T_9708 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9711 = _T_9709 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9721 = _T_5205 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9724 = _T_9178 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9725 = _T_9721 | _T_9724; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9726 = _T_9725 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9728 = _T_9726 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9738 = _T_5209 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9741 = _T_9195 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9742 = _T_9738 | _T_9741; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9743 = _T_9742 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9745 = _T_9743 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9755 = _T_5213 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9758 = _T_9212 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9759 = _T_9755 | _T_9758; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9760 = _T_9759 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9762 = _T_9760 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9772 = _T_5217 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9775 = _T_9229 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9776 = _T_9772 | _T_9775; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9777 = _T_9776 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9779 = _T_9777 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9789 = _T_5221 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9792 = _T_9246 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9793 = _T_9789 | _T_9792; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9794 = _T_9793 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9796 = _T_9794 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9806 = _T_5225 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9809 = _T_9263 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9810 = _T_9806 | _T_9809; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9811 = _T_9810 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9813 = _T_9811 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9823 = _T_5229 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9826 = _T_9280 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9827 = _T_9823 | _T_9826; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9828 = _T_9827 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9830 = _T_9828 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9840 = _T_5233 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9843 = _T_9297 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9844 = _T_9840 | _T_9843; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9845 = _T_9844 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9847 = _T_9845 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9857 = _T_5237 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9860 = _T_9314 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9861 = _T_9857 | _T_9860; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9862 = _T_9861 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9864 = _T_9862 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9874 = _T_5241 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9877 = _T_9331 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9878 = _T_9874 | _T_9877; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9879 = _T_9878 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9881 = _T_9879 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9891 = _T_5245 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9894 = _T_9348 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9895 = _T_9891 | _T_9894; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9896 = _T_9895 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9898 = _T_9896 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9908 = _T_5249 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9911 = _T_9365 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9912 = _T_9908 | _T_9911; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9913 = _T_9912 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9915 = _T_9913 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9925 = _T_5253 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9928 = _T_9382 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9929 = _T_9925 | _T_9928; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9930 = _T_9929 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9932 = _T_9930 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9942 = _T_5257 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9945 = _T_9399 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9946 = _T_9942 | _T_9945; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9947 = _T_9946 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9949 = _T_9947 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9959 = _T_5261 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9962 = _T_9416 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9963 = _T_9959 | _T_9962; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9964 = _T_9963 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9966 = _T_9964 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9976 = _T_5265 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9979 = _T_9433 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9980 = _T_9976 | _T_9979; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9981 = _T_9980 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_9983 = _T_9981 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_9993 = _T_5269 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_9996 = _T_9450 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_9997 = _T_9993 | _T_9996; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_9998 = _T_9997 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10000 = _T_9998 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10010 = _T_5273 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_10013 = _T_9467 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_10014 = _T_10010 | _T_10013; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_10015 = _T_10014 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10017 = _T_10015 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10027 = _T_5277 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_10030 = _T_9484 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_10031 = _T_10027 | _T_10030; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_10032 = _T_10031 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10034 = _T_10032 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10044 = _T_5281 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_10047 = _T_9501 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_10048 = _T_10044 | _T_10047; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_10049 = _T_10048 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10051 = _T_10049 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10061 = _T_5285 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_10064 = _T_9518 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_10065 = _T_10061 | _T_10064; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_10066 = _T_10065 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10068 = _T_10066 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10078 = _T_5289 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_10081 = _T_9535 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_10082 = _T_10078 | _T_10081; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_10083 = _T_10082 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10085 = _T_10083 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10095 = _T_5293 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_10098 = _T_9552 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_10099 = _T_10095 | _T_10098; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_10100 = _T_10099 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10102 = _T_10100 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10112 = _T_5297 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 761:59]
  wire  _T_10115 = _T_9569 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 761:124]
  wire  _T_10116 = _T_10112 | _T_10115; // @[el2_ifu_mem_ctl.scala 761:81]
  wire  _T_10117 = _T_10116 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 761:147]
  wire  _T_10119 = _T_10117 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 761:165]
  wire  _T_10921 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 816:63]
  wire  _T_10922 = _T_10921 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 816:85]
  wire [1:0] _T_10924 = _T_10922 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10931; // @[el2_ifu_mem_ctl.scala 821:57]
  reg  _T_10932; // @[el2_ifu_mem_ctl.scala 822:56]
  reg  _T_10933; // @[el2_ifu_mem_ctl.scala 823:59]
  wire  _T_10934 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 824:80]
  wire  _T_10935 = ifu_bus_arvalid_ff & _T_10934; // @[el2_ifu_mem_ctl.scala 824:78]
  wire  _T_10936 = _T_10935 & miss_pending; // @[el2_ifu_mem_ctl.scala 824:100]
  reg  _T_10937; // @[el2_ifu_mem_ctl.scala 824:58]
  reg  _T_10938; // @[el2_ifu_mem_ctl.scala 825:58]
  wire  _T_10941 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 832:71]
  wire  _T_10943 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 832:124]
  wire  _T_10945 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 833:50]
  wire  _T_10947 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 833:103]
  wire [3:0] _T_10950 = {_T_10941,_T_10943,_T_10945,_T_10947}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 835:53]
  reg  _T_10961; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 332:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 331:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 196:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3978; // @[el2_ifu_mem_ctl.scala 702:21]
  assign io_ifu_pmu_ic_miss = _T_10931; // @[el2_ifu_mem_ctl.scala 821:22]
  assign io_ifu_pmu_ic_hit = _T_10932; // @[el2_ifu_mem_ctl.scala 822:21]
  assign io_ifu_pmu_bus_error = _T_10933; // @[el2_ifu_mem_ctl.scala 823:24]
  assign io_ifu_pmu_bus_busy = _T_10937; // @[el2_ifu_mem_ctl.scala 824:23]
  assign io_ifu_pmu_bus_trxn = _T_10938; // @[el2_ifu_mem_ctl.scala 825:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 146:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 145:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 144:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 142:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 153:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 155:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 148:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 141:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 138:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 147:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 156:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 151:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 564:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2572; // @[el2_ifu_mem_ctl.scala 565:19]
  assign io_ifu_axi_araddr = _T_2574 & _T_2576; // @[el2_ifu_mem_ctl.scala 566:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 569:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 152:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 567:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 570:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 143:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 568:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 154:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 149:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 571:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 661:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 659:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 663:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 654:20]
  assign io_iccm_ready = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 634:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 341:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3964; // @[el2_ifu_mem_ctl.scala 701:15]
  assign io_ic_rd_en = _T_3956 | _T_3961; // @[el2_ifu_mem_ctl.scala 692:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 348:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 348:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 349:23]
  assign io_ifu_ic_debug_rd_data = _T_1209; // @[el2_ifu_mem_ctl.scala 357:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 828:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 830:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 831:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 829:25]
  assign io_ic_debug_way = _T_10950[1:0]; // @[el2_ifu_mem_ctl.scala 832:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10924; // @[el2_ifu_mem_ctl.scala 816:19]
  assign io_iccm_rw_addr = _T_3110[14:0]; // @[el2_ifu_mem_ctl.scala 665:19]
  assign io_iccm_wren = _T_2679 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 636:16]
  assign io_iccm_rden = _T_2683 | _T_2684; // @[el2_ifu_mem_ctl.scala 637:16]
  assign io_iccm_wr_data = _T_3085 ? _T_3086 : _T_3093; // @[el2_ifu_mem_ctl.scala 642:19]
  assign io_iccm_wr_size = _T_2689 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 639:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 293:15]
  assign io_ic_access_fault_f = _T_2457 & _T_317; // @[el2_ifu_mem_ctl.scala 389:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1271; // @[el2_ifu_mem_ctl.scala 390:29]
  assign io_iccm_rd_ecc_single_err = _T_3901 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 678:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 679:29]
  assign io_ic_error_start = _T_1197 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 351:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 195:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 194:24]
  assign io_ic_fetch_val_f = {_T_1279,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 393:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 386:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 383:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 384:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10961; // @[el2_ifu_mem_ctl.scala 839:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2462; // @[el2_ifu_mem_ctl.scala 483:27]
  assign io_iccm_correction_state = _T_2490 ? 1'h0 : _GEN_60; // @[el2_ifu_mem_ctl.scala 518:28 el2_ifu_mem_ctl.scala 531:32 el2_ifu_mem_ctl.scala 538:32 el2_ifu_mem_ctl.scala 545:32]
  assign io_valids = {_T_5641,_T_5768}; // @[el2_ifu_mem_ctl.scala 756:15]
  assign io_tagv_mb_in = scnd_miss_req ? _T_290 : _T_296; // @[el2_ifu_mem_ctl.scala 854:17]
  assign io_test = _T_3990 ? io_ic_debug_wr_data[4] : way_status_new; // @[el2_ifu_mem_ctl.scala 720:11]
  assign io_test_way_status_out = {_T_4774,way_status_out_0}; // @[el2_ifu_mem_ctl.scala 730:26]
  assign io_test_way_status_clken = {_T_4788,way_status_clken_0}; // @[el2_ifu_mem_ctl.scala 732:28]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_127 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_126 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_125 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_124 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_123 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_122 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_121 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_120 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_119 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_118 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_117 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_116 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_115 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_114 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_113 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_112 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_111 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_110 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_109 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_108 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_107 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_106 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_105 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_104 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_103 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_102 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_101 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_100 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_99 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_98 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_97 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_96 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_95 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_94 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_93 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_92 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_91 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_90 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_89 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_88 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_87 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_86 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_85 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_84 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_83 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_82 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_81 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_80 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_79 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_78 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_77 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_76 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_75 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_74 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_73 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_72 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_71 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_70 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_69 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_68 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_67 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_66 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_65 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_64 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_63 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_62 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_61 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_60 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_59 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_58 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_57 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_56 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_55 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_54 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_53 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_52 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_51 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_50 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_49 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_48 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_47 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_46 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_45 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_44 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_43 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_42 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_41 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_40 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_39 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_38 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_37 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_36 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_35 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_34 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_33 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_32 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_31 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_30 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_29 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_28 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_27 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_26 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_25 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_24 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_23 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_22 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_21 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_20 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_19 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_18 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_17 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_16 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_15 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_14 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_13 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_12 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_11 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_10 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_9 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_8 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_7 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_6 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_5 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_4 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_3 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_2 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_0 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1209 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_443[6:0];
  _RAND_444 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_446[2:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_449[0:0];
  _RAND_450 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_450[38:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_453[2:0];
  _RAND_454 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_454[0:0];
  _RAND_455 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_455[63:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_456[13:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_458[13:0];
  _RAND_459 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_459[6:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way_status_new_ff = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  ic_valid_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10931 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10932 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10933 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10937 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10938 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_10961 = _RAND_469[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4647) begin
      way_status_out_127 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4642) begin
      way_status_out_126 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4637) begin
      way_status_out_125 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4632) begin
      way_status_out_124 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4627) begin
      way_status_out_123 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4622) begin
      way_status_out_122 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4617) begin
      way_status_out_121 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4612) begin
      way_status_out_120 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4607) begin
      way_status_out_119 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4602) begin
      way_status_out_118 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4597) begin
      way_status_out_117 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4592) begin
      way_status_out_116 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4587) begin
      way_status_out_115 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4582) begin
      way_status_out_114 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4577) begin
      way_status_out_113 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4572) begin
      way_status_out_112 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4567) begin
      way_status_out_111 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4562) begin
      way_status_out_110 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4557) begin
      way_status_out_109 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4552) begin
      way_status_out_108 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4547) begin
      way_status_out_107 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4542) begin
      way_status_out_106 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4537) begin
      way_status_out_105 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4532) begin
      way_status_out_104 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4527) begin
      way_status_out_103 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4522) begin
      way_status_out_102 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4517) begin
      way_status_out_101 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4512) begin
      way_status_out_100 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4507) begin
      way_status_out_99 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4502) begin
      way_status_out_98 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4497) begin
      way_status_out_97 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4492) begin
      way_status_out_96 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4487) begin
      way_status_out_95 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4482) begin
      way_status_out_94 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4477) begin
      way_status_out_93 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4472) begin
      way_status_out_92 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4467) begin
      way_status_out_91 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4462) begin
      way_status_out_90 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4457) begin
      way_status_out_89 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4452) begin
      way_status_out_88 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4447) begin
      way_status_out_87 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4442) begin
      way_status_out_86 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4437) begin
      way_status_out_85 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4432) begin
      way_status_out_84 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4427) begin
      way_status_out_83 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4422) begin
      way_status_out_82 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4417) begin
      way_status_out_81 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4412) begin
      way_status_out_80 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4407) begin
      way_status_out_79 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4402) begin
      way_status_out_78 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4397) begin
      way_status_out_77 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4392) begin
      way_status_out_76 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4387) begin
      way_status_out_75 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4382) begin
      way_status_out_74 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4377) begin
      way_status_out_73 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4372) begin
      way_status_out_72 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4367) begin
      way_status_out_71 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4362) begin
      way_status_out_70 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4357) begin
      way_status_out_69 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4352) begin
      way_status_out_68 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4347) begin
      way_status_out_67 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4342) begin
      way_status_out_66 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4337) begin
      way_status_out_65 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4332) begin
      way_status_out_64 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4327) begin
      way_status_out_63 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4322) begin
      way_status_out_62 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4317) begin
      way_status_out_61 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4312) begin
      way_status_out_60 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4307) begin
      way_status_out_59 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4302) begin
      way_status_out_58 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4297) begin
      way_status_out_57 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4292) begin
      way_status_out_56 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4287) begin
      way_status_out_55 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4282) begin
      way_status_out_54 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4277) begin
      way_status_out_53 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4272) begin
      way_status_out_52 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4267) begin
      way_status_out_51 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4262) begin
      way_status_out_50 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4257) begin
      way_status_out_49 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4252) begin
      way_status_out_48 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4247) begin
      way_status_out_47 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4242) begin
      way_status_out_46 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4237) begin
      way_status_out_45 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4232) begin
      way_status_out_44 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4227) begin
      way_status_out_43 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4222) begin
      way_status_out_42 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4217) begin
      way_status_out_41 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4212) begin
      way_status_out_40 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4207) begin
      way_status_out_39 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4202) begin
      way_status_out_38 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4197) begin
      way_status_out_37 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4192) begin
      way_status_out_36 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4187) begin
      way_status_out_35 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4182) begin
      way_status_out_34 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4177) begin
      way_status_out_33 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4172) begin
      way_status_out_32 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4167) begin
      way_status_out_31 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4162) begin
      way_status_out_30 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4157) begin
      way_status_out_29 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4152) begin
      way_status_out_28 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4147) begin
      way_status_out_27 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4142) begin
      way_status_out_26 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4137) begin
      way_status_out_25 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4132) begin
      way_status_out_24 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4127) begin
      way_status_out_23 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4122) begin
      way_status_out_22 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4117) begin
      way_status_out_21 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4112) begin
      way_status_out_20 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4107) begin
      way_status_out_19 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4102) begin
      way_status_out_18 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4097) begin
      way_status_out_17 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4092) begin
      way_status_out_16 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4087) begin
      way_status_out_15 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4082) begin
      way_status_out_14 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4077) begin
      way_status_out_13 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4072) begin
      way_status_out_12 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4067) begin
      way_status_out_11 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4062) begin
      way_status_out_10 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4057) begin
      way_status_out_9 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4052) begin
      way_status_out_8 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4047) begin
      way_status_out_7 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4042) begin
      way_status_out_6 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4037) begin
      way_status_out_5 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4032) begin
      way_status_out_4 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4027) begin
      way_status_out_3 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_4022) begin
      way_status_out_2 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_4017) begin
      way_status_out_1 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_4012) begin
      way_status_out_0 <= way_status_new_ff;
    end
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2615) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2611;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_6328) begin
      ic_tag_valid_out_1_0 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_6345) begin
      ic_tag_valid_out_1_1 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_6362) begin
      ic_tag_valid_out_1_2 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_6379) begin
      ic_tag_valid_out_1_3 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_6396) begin
      ic_tag_valid_out_1_4 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_6413) begin
      ic_tag_valid_out_1_5 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_6430) begin
      ic_tag_valid_out_1_6 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_6447) begin
      ic_tag_valid_out_1_7 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_6464) begin
      ic_tag_valid_out_1_8 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_6481) begin
      ic_tag_valid_out_1_9 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_6498) begin
      ic_tag_valid_out_1_10 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_6515) begin
      ic_tag_valid_out_1_11 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_6532) begin
      ic_tag_valid_out_1_12 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_6549) begin
      ic_tag_valid_out_1_13 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_6566) begin
      ic_tag_valid_out_1_14 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_6583) begin
      ic_tag_valid_out_1_15 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_6600) begin
      ic_tag_valid_out_1_16 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_6617) begin
      ic_tag_valid_out_1_17 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6634) begin
      ic_tag_valid_out_1_18 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6651) begin
      ic_tag_valid_out_1_19 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6668) begin
      ic_tag_valid_out_1_20 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6685) begin
      ic_tag_valid_out_1_21 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6702) begin
      ic_tag_valid_out_1_22 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6719) begin
      ic_tag_valid_out_1_23 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6736) begin
      ic_tag_valid_out_1_24 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6753) begin
      ic_tag_valid_out_1_25 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6770) begin
      ic_tag_valid_out_1_26 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6787) begin
      ic_tag_valid_out_1_27 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6804) begin
      ic_tag_valid_out_1_28 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6821) begin
      ic_tag_valid_out_1_29 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6838) begin
      ic_tag_valid_out_1_30 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6855) begin
      ic_tag_valid_out_1_31 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_7416) begin
      ic_tag_valid_out_1_32 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_7433) begin
      ic_tag_valid_out_1_33 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_7450) begin
      ic_tag_valid_out_1_34 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_7467) begin
      ic_tag_valid_out_1_35 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_7484) begin
      ic_tag_valid_out_1_36 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_7501) begin
      ic_tag_valid_out_1_37 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_7518) begin
      ic_tag_valid_out_1_38 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_7535) begin
      ic_tag_valid_out_1_39 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_7552) begin
      ic_tag_valid_out_1_40 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_7569) begin
      ic_tag_valid_out_1_41 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_7586) begin
      ic_tag_valid_out_1_42 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_7603) begin
      ic_tag_valid_out_1_43 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_7620) begin
      ic_tag_valid_out_1_44 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_7637) begin
      ic_tag_valid_out_1_45 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_7654) begin
      ic_tag_valid_out_1_46 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_7671) begin
      ic_tag_valid_out_1_47 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7688) begin
      ic_tag_valid_out_1_48 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7705) begin
      ic_tag_valid_out_1_49 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7722) begin
      ic_tag_valid_out_1_50 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7739) begin
      ic_tag_valid_out_1_51 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7756) begin
      ic_tag_valid_out_1_52 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7773) begin
      ic_tag_valid_out_1_53 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7790) begin
      ic_tag_valid_out_1_54 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7807) begin
      ic_tag_valid_out_1_55 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7824) begin
      ic_tag_valid_out_1_56 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7841) begin
      ic_tag_valid_out_1_57 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7858) begin
      ic_tag_valid_out_1_58 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7875) begin
      ic_tag_valid_out_1_59 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7892) begin
      ic_tag_valid_out_1_60 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7909) begin
      ic_tag_valid_out_1_61 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7926) begin
      ic_tag_valid_out_1_62 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7943) begin
      ic_tag_valid_out_1_63 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_8504) begin
      ic_tag_valid_out_1_64 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_8521) begin
      ic_tag_valid_out_1_65 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_8538) begin
      ic_tag_valid_out_1_66 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_8555) begin
      ic_tag_valid_out_1_67 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_8572) begin
      ic_tag_valid_out_1_68 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_8589) begin
      ic_tag_valid_out_1_69 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_8606) begin
      ic_tag_valid_out_1_70 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_8623) begin
      ic_tag_valid_out_1_71 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_8640) begin
      ic_tag_valid_out_1_72 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_8657) begin
      ic_tag_valid_out_1_73 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_8674) begin
      ic_tag_valid_out_1_74 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_8691) begin
      ic_tag_valid_out_1_75 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_8708) begin
      ic_tag_valid_out_1_76 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_8725) begin
      ic_tag_valid_out_1_77 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_8742) begin
      ic_tag_valid_out_1_78 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8759) begin
      ic_tag_valid_out_1_79 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8776) begin
      ic_tag_valid_out_1_80 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8793) begin
      ic_tag_valid_out_1_81 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8810) begin
      ic_tag_valid_out_1_82 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8827) begin
      ic_tag_valid_out_1_83 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8844) begin
      ic_tag_valid_out_1_84 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8861) begin
      ic_tag_valid_out_1_85 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8878) begin
      ic_tag_valid_out_1_86 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8895) begin
      ic_tag_valid_out_1_87 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8912) begin
      ic_tag_valid_out_1_88 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8929) begin
      ic_tag_valid_out_1_89 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8946) begin
      ic_tag_valid_out_1_90 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8963) begin
      ic_tag_valid_out_1_91 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8980) begin
      ic_tag_valid_out_1_92 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8997) begin
      ic_tag_valid_out_1_93 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_9014) begin
      ic_tag_valid_out_1_94 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_9031) begin
      ic_tag_valid_out_1_95 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_9592) begin
      ic_tag_valid_out_1_96 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_9609) begin
      ic_tag_valid_out_1_97 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_9626) begin
      ic_tag_valid_out_1_98 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_9643) begin
      ic_tag_valid_out_1_99 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_9660) begin
      ic_tag_valid_out_1_100 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_9677) begin
      ic_tag_valid_out_1_101 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_9694) begin
      ic_tag_valid_out_1_102 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_9711) begin
      ic_tag_valid_out_1_103 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_9728) begin
      ic_tag_valid_out_1_104 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_9745) begin
      ic_tag_valid_out_1_105 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_9762) begin
      ic_tag_valid_out_1_106 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_9779) begin
      ic_tag_valid_out_1_107 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_9796) begin
      ic_tag_valid_out_1_108 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9813) begin
      ic_tag_valid_out_1_109 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9830) begin
      ic_tag_valid_out_1_110 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9847) begin
      ic_tag_valid_out_1_111 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9864) begin
      ic_tag_valid_out_1_112 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9881) begin
      ic_tag_valid_out_1_113 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9898) begin
      ic_tag_valid_out_1_114 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9915) begin
      ic_tag_valid_out_1_115 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9932) begin
      ic_tag_valid_out_1_116 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9949) begin
      ic_tag_valid_out_1_117 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9966) begin
      ic_tag_valid_out_1_118 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9983) begin
      ic_tag_valid_out_1_119 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_10000) begin
      ic_tag_valid_out_1_120 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_10017) begin
      ic_tag_valid_out_1_121 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_10034) begin
      ic_tag_valid_out_1_122 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_10051) begin
      ic_tag_valid_out_1_123 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_10068) begin
      ic_tag_valid_out_1_124 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_10085) begin
      ic_tag_valid_out_1_125 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_10102) begin
      ic_tag_valid_out_1_126 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_10119) begin
      ic_tag_valid_out_1_127 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5784) begin
      ic_tag_valid_out_0_0 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5801) begin
      ic_tag_valid_out_0_1 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5818) begin
      ic_tag_valid_out_0_2 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5835) begin
      ic_tag_valid_out_0_3 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5852) begin
      ic_tag_valid_out_0_4 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5869) begin
      ic_tag_valid_out_0_5 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5886) begin
      ic_tag_valid_out_0_6 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5903) begin
      ic_tag_valid_out_0_7 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5920) begin
      ic_tag_valid_out_0_8 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5937) begin
      ic_tag_valid_out_0_9 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5954) begin
      ic_tag_valid_out_0_10 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5971) begin
      ic_tag_valid_out_0_11 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5988) begin
      ic_tag_valid_out_0_12 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_6005) begin
      ic_tag_valid_out_0_13 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_6022) begin
      ic_tag_valid_out_0_14 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_6039) begin
      ic_tag_valid_out_0_15 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_6056) begin
      ic_tag_valid_out_0_16 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_6073) begin
      ic_tag_valid_out_0_17 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_6090) begin
      ic_tag_valid_out_0_18 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_6107) begin
      ic_tag_valid_out_0_19 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_6124) begin
      ic_tag_valid_out_0_20 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_6141) begin
      ic_tag_valid_out_0_21 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_6158) begin
      ic_tag_valid_out_0_22 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_6175) begin
      ic_tag_valid_out_0_23 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_6192) begin
      ic_tag_valid_out_0_24 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_6209) begin
      ic_tag_valid_out_0_25 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_6226) begin
      ic_tag_valid_out_0_26 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_6243) begin
      ic_tag_valid_out_0_27 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_6260) begin
      ic_tag_valid_out_0_28 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_6277) begin
      ic_tag_valid_out_0_29 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_6294) begin
      ic_tag_valid_out_0_30 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_6311) begin
      ic_tag_valid_out_0_31 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6872) begin
      ic_tag_valid_out_0_32 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6889) begin
      ic_tag_valid_out_0_33 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6906) begin
      ic_tag_valid_out_0_34 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6923) begin
      ic_tag_valid_out_0_35 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6940) begin
      ic_tag_valid_out_0_36 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6957) begin
      ic_tag_valid_out_0_37 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6974) begin
      ic_tag_valid_out_0_38 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6991) begin
      ic_tag_valid_out_0_39 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_7008) begin
      ic_tag_valid_out_0_40 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_7025) begin
      ic_tag_valid_out_0_41 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_7042) begin
      ic_tag_valid_out_0_42 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_7059) begin
      ic_tag_valid_out_0_43 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_7076) begin
      ic_tag_valid_out_0_44 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_7093) begin
      ic_tag_valid_out_0_45 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_7110) begin
      ic_tag_valid_out_0_46 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_7127) begin
      ic_tag_valid_out_0_47 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_7144) begin
      ic_tag_valid_out_0_48 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_7161) begin
      ic_tag_valid_out_0_49 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_7178) begin
      ic_tag_valid_out_0_50 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_7195) begin
      ic_tag_valid_out_0_51 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_7212) begin
      ic_tag_valid_out_0_52 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_7229) begin
      ic_tag_valid_out_0_53 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_7246) begin
      ic_tag_valid_out_0_54 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_7263) begin
      ic_tag_valid_out_0_55 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_7280) begin
      ic_tag_valid_out_0_56 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_7297) begin
      ic_tag_valid_out_0_57 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_7314) begin
      ic_tag_valid_out_0_58 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_7331) begin
      ic_tag_valid_out_0_59 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_7348) begin
      ic_tag_valid_out_0_60 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_7365) begin
      ic_tag_valid_out_0_61 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_7382) begin
      ic_tag_valid_out_0_62 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_7399) begin
      ic_tag_valid_out_0_63 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7960) begin
      ic_tag_valid_out_0_64 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7977) begin
      ic_tag_valid_out_0_65 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7994) begin
      ic_tag_valid_out_0_66 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_8011) begin
      ic_tag_valid_out_0_67 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_8028) begin
      ic_tag_valid_out_0_68 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_8045) begin
      ic_tag_valid_out_0_69 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_8062) begin
      ic_tag_valid_out_0_70 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_8079) begin
      ic_tag_valid_out_0_71 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_8096) begin
      ic_tag_valid_out_0_72 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_8113) begin
      ic_tag_valid_out_0_73 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_8130) begin
      ic_tag_valid_out_0_74 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_8147) begin
      ic_tag_valid_out_0_75 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_8164) begin
      ic_tag_valid_out_0_76 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_8181) begin
      ic_tag_valid_out_0_77 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_8198) begin
      ic_tag_valid_out_0_78 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_8215) begin
      ic_tag_valid_out_0_79 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_8232) begin
      ic_tag_valid_out_0_80 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_8249) begin
      ic_tag_valid_out_0_81 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_8266) begin
      ic_tag_valid_out_0_82 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_8283) begin
      ic_tag_valid_out_0_83 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_8300) begin
      ic_tag_valid_out_0_84 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_8317) begin
      ic_tag_valid_out_0_85 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_8334) begin
      ic_tag_valid_out_0_86 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_8351) begin
      ic_tag_valid_out_0_87 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_8368) begin
      ic_tag_valid_out_0_88 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_8385) begin
      ic_tag_valid_out_0_89 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_8402) begin
      ic_tag_valid_out_0_90 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_8419) begin
      ic_tag_valid_out_0_91 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_8436) begin
      ic_tag_valid_out_0_92 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_8453) begin
      ic_tag_valid_out_0_93 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_8470) begin
      ic_tag_valid_out_0_94 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_8487) begin
      ic_tag_valid_out_0_95 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_9048) begin
      ic_tag_valid_out_0_96 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_9065) begin
      ic_tag_valid_out_0_97 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_9082) begin
      ic_tag_valid_out_0_98 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_9099) begin
      ic_tag_valid_out_0_99 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_9116) begin
      ic_tag_valid_out_0_100 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_9133) begin
      ic_tag_valid_out_0_101 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_9150) begin
      ic_tag_valid_out_0_102 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_9167) begin
      ic_tag_valid_out_0_103 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_9184) begin
      ic_tag_valid_out_0_104 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_9201) begin
      ic_tag_valid_out_0_105 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_9218) begin
      ic_tag_valid_out_0_106 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_9235) begin
      ic_tag_valid_out_0_107 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_9252) begin
      ic_tag_valid_out_0_108 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_9269) begin
      ic_tag_valid_out_0_109 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_9286) begin
      ic_tag_valid_out_0_110 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_9303) begin
      ic_tag_valid_out_0_111 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_9320) begin
      ic_tag_valid_out_0_112 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_9337) begin
      ic_tag_valid_out_0_113 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_9354) begin
      ic_tag_valid_out_0_114 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_9371) begin
      ic_tag_valid_out_0_115 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_9388) begin
      ic_tag_valid_out_0_116 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_9405) begin
      ic_tag_valid_out_0_117 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_9422) begin
      ic_tag_valid_out_0_118 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_9439) begin
      ic_tag_valid_out_0_119 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_9456) begin
      ic_tag_valid_out_0_120 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_9473) begin
      ic_tag_valid_out_0_121 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_9490) begin
      ic_tag_valid_out_0_122 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_9507) begin
      ic_tag_valid_out_0_123 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_9524) begin
      ic_tag_valid_out_0_124 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_9541) begin
      ic_tag_valid_out_0_125 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_9558) begin
      ic_tag_valid_out_0_126 <= _T_5774;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_9575) begin
      ic_tag_valid_out_0_127 <= _T_5774;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1209 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_1209 <= {{5'd0}, _T_1208};
      end else begin
        _T_1209 <= io_ic_debug_rd_data;
      end
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2564) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2639) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2683;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2465) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2467) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2477) begin
        perr_state <= 3'h0;
      end else if (_T_2480) begin
        if (_T_2482) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2486) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2490) begin
        err_stop_state <= 2'h1;
      end else if (_T_2495) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (_T_2518) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2522) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2539) begin
        if (_T_2543) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1368;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3987) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1408;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3922;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3097;
    end else begin
      iccm_dma_rdata <= _T_3098;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3918;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3987) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_3990) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_10909) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3990) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10961 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10961 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10931 <= 1'h0;
    end else begin
      _T_10931 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10932 <= 1'h0;
    end else begin
      _T_10932 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10933 <= 1'h0;
    end else begin
      _T_10933 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10937 <= 1'h0;
    end else begin
      _T_10937 <= _T_10936;
    end
    if (reset) begin
      _T_10938 <= 1'h0;
    end else begin
      _T_10938 <= bus_cmd_sent;
    end
  end
endmodule
