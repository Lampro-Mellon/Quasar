module el2_lsu_trigger(
  input         clock,
  input         reset,
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input         io_trigger_pkt_any_0_execute,
  input         io_trigger_pkt_any_0_m,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input         io_trigger_pkt_any_1_execute,
  input         io_trigger_pkt_any_1_m,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input         io_trigger_pkt_any_2_execute,
  input         io_trigger_pkt_any_2_m,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input         io_trigger_pkt_any_3_execute,
  input         io_trigger_pkt_any_3_m,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_lsu_pkt_m_fast_int,
  input         io_lsu_pkt_m_by,
  input         io_lsu_pkt_m_half,
  input         io_lsu_pkt_m_word,
  input         io_lsu_pkt_m_dword,
  input         io_lsu_pkt_m_load,
  input         io_lsu_pkt_m_store,
  input         io_lsu_pkt_m_unsign,
  input         io_lsu_pkt_m_dma,
  input         io_lsu_pkt_m_store_data_bypass_d,
  input         io_lsu_pkt_m_load_ldst_bypass_d,
  input         io_lsu_pkt_m_store_data_bypass_m,
  input         io_lsu_pkt_m_valid,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_store_data_m,
  output [3:0]  io_lsu_trigger_match_m
);
  wire [15:0] _T_1 = io_lsu_pkt_m_word ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_3 = _T_1 & io_store_data_m[31:16]; // @[el2_lsu_trigger.scala 18:61]
  wire  _T_4 = io_lsu_pkt_m_half | io_lsu_pkt_m_word; // @[el2_lsu_trigger.scala 18:114]
  wire [7:0] _T_6 = _T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_8 = _T_6 & io_store_data_m[15:8]; // @[el2_lsu_trigger.scala 18:136]
  wire [31:0] store_data_trigger_m = {_T_3,_T_8,io_store_data_m[7:0]}; // @[Cat.scala 29:58]
  wire  _T_11 = ~io_trigger_pkt_any_0_select; // @[el2_lsu_trigger.scala 20:57]
  wire [31:0] _T_13 = _T_11 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_14 = _T_13 & io_lsu_addr_m; // @[el2_lsu_trigger.scala 20:88]
  wire [31:0] _T_16 = io_trigger_pkt_any_0_select ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _GEN_0 = {{31'd0}, io_trigger_pkt_any_0_store}; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_17 = _T_16 & _GEN_0; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_18 = _T_17 & store_data_trigger_m; // @[el2_lsu_trigger.scala 20:179]
  wire [31:0] lsu_match_data_0 = _T_14 | _T_18; // @[el2_lsu_trigger.scala 20:105]
  wire  _T_20 = ~io_trigger_pkt_any_1_select; // @[el2_lsu_trigger.scala 20:57]
  wire [31:0] _T_22 = _T_20 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_23 = _T_22 & io_lsu_addr_m; // @[el2_lsu_trigger.scala 20:88]
  wire [31:0] _T_25 = io_trigger_pkt_any_1_select ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _GEN_1 = {{31'd0}, io_trigger_pkt_any_1_store}; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_26 = _T_25 & _GEN_1; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_27 = _T_26 & store_data_trigger_m; // @[el2_lsu_trigger.scala 20:179]
  wire [31:0] lsu_match_data_1 = _T_23 | _T_27; // @[el2_lsu_trigger.scala 20:105]
  wire  _T_29 = ~io_trigger_pkt_any_2_select; // @[el2_lsu_trigger.scala 20:57]
  wire [31:0] _T_31 = _T_29 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_32 = _T_31 & io_lsu_addr_m; // @[el2_lsu_trigger.scala 20:88]
  wire [31:0] _T_34 = io_trigger_pkt_any_2_select ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _GEN_2 = {{31'd0}, io_trigger_pkt_any_2_store}; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_35 = _T_34 & _GEN_2; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_36 = _T_35 & store_data_trigger_m; // @[el2_lsu_trigger.scala 20:179]
  wire [31:0] lsu_match_data_2 = _T_32 | _T_36; // @[el2_lsu_trigger.scala 20:105]
  wire  _T_38 = ~io_trigger_pkt_any_3_select; // @[el2_lsu_trigger.scala 20:57]
  wire [31:0] _T_40 = _T_38 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_41 = _T_40 & io_lsu_addr_m; // @[el2_lsu_trigger.scala 20:88]
  wire [31:0] _T_43 = io_trigger_pkt_any_3_select ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _GEN_3 = {{31'd0}, io_trigger_pkt_any_3_store}; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_44 = _T_43 & _GEN_3; // @[el2_lsu_trigger.scala 20:148]
  wire [31:0] _T_45 = _T_44 & store_data_trigger_m; // @[el2_lsu_trigger.scala 20:179]
  wire [31:0] lsu_match_data_3 = _T_41 | _T_45; // @[el2_lsu_trigger.scala 20:105]
  wire  _T_48 = ~io_lsu_pkt_m_dma; // @[el2_lsu_trigger.scala 21:71]
  wire  _T_49 = io_lsu_pkt_m_valid & _T_48; // @[el2_lsu_trigger.scala 21:69]
  wire  _T_50 = io_trigger_pkt_any_0_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 21:120]
  wire  _T_51 = _T_49 & _T_50; // @[el2_lsu_trigger.scala 21:89]
  wire  _T_52 = io_trigger_pkt_any_0_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 22:33]
  wire  _T_54 = _T_52 & _T_11; // @[el2_lsu_trigger.scala 22:53]
  wire  _T_57 = &io_trigger_pkt_any_0_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_58 = ~_T_57; // @[el2_lib.scala 194:39]
  wire  _T_59 = io_trigger_pkt_any_0_match_ & _T_58; // @[el2_lib.scala 194:37]
  wire  _T_62 = io_trigger_pkt_any_0_tdata2[0] == lsu_match_data_0[0]; // @[el2_lib.scala 195:52]
  wire  _T_63 = _T_59 | _T_62; // @[el2_lib.scala 195:41]
  wire  _T_65 = &io_trigger_pkt_any_0_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_66 = _T_65 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_69 = io_trigger_pkt_any_0_tdata2[1] == lsu_match_data_0[1]; // @[el2_lib.scala 197:80]
  wire  _T_70 = _T_66 | _T_69; // @[el2_lib.scala 197:25]
  wire  _T_72 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_73 = _T_72 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_76 = io_trigger_pkt_any_0_tdata2[2] == lsu_match_data_0[2]; // @[el2_lib.scala 197:80]
  wire  _T_77 = _T_73 | _T_76; // @[el2_lib.scala 197:25]
  wire  _T_79 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_80 = _T_79 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_83 = io_trigger_pkt_any_0_tdata2[3] == lsu_match_data_0[3]; // @[el2_lib.scala 197:80]
  wire  _T_84 = _T_80 | _T_83; // @[el2_lib.scala 197:25]
  wire  _T_86 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_87 = _T_86 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_90 = io_trigger_pkt_any_0_tdata2[4] == lsu_match_data_0[4]; // @[el2_lib.scala 197:80]
  wire  _T_91 = _T_87 | _T_90; // @[el2_lib.scala 197:25]
  wire  _T_93 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_94 = _T_93 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_97 = io_trigger_pkt_any_0_tdata2[5] == lsu_match_data_0[5]; // @[el2_lib.scala 197:80]
  wire  _T_98 = _T_94 | _T_97; // @[el2_lib.scala 197:25]
  wire  _T_100 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_101 = _T_100 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_104 = io_trigger_pkt_any_0_tdata2[6] == lsu_match_data_0[6]; // @[el2_lib.scala 197:80]
  wire  _T_105 = _T_101 | _T_104; // @[el2_lib.scala 197:25]
  wire  _T_107 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_108 = _T_107 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_111 = io_trigger_pkt_any_0_tdata2[7] == lsu_match_data_0[7]; // @[el2_lib.scala 197:80]
  wire  _T_112 = _T_108 | _T_111; // @[el2_lib.scala 197:25]
  wire  _T_114 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_115 = _T_114 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_118 = io_trigger_pkt_any_0_tdata2[8] == lsu_match_data_0[8]; // @[el2_lib.scala 197:80]
  wire  _T_119 = _T_115 | _T_118; // @[el2_lib.scala 197:25]
  wire  _T_121 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_122 = _T_121 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_125 = io_trigger_pkt_any_0_tdata2[9] == lsu_match_data_0[9]; // @[el2_lib.scala 197:80]
  wire  _T_126 = _T_122 | _T_125; // @[el2_lib.scala 197:25]
  wire  _T_128 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_129 = _T_128 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_132 = io_trigger_pkt_any_0_tdata2[10] == lsu_match_data_0[10]; // @[el2_lib.scala 197:80]
  wire  _T_133 = _T_129 | _T_132; // @[el2_lib.scala 197:25]
  wire  _T_135 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_136 = _T_135 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_139 = io_trigger_pkt_any_0_tdata2[11] == lsu_match_data_0[11]; // @[el2_lib.scala 197:80]
  wire  _T_140 = _T_136 | _T_139; // @[el2_lib.scala 197:25]
  wire  _T_142 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_143 = _T_142 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_146 = io_trigger_pkt_any_0_tdata2[12] == lsu_match_data_0[12]; // @[el2_lib.scala 197:80]
  wire  _T_147 = _T_143 | _T_146; // @[el2_lib.scala 197:25]
  wire  _T_149 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_150 = _T_149 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_153 = io_trigger_pkt_any_0_tdata2[13] == lsu_match_data_0[13]; // @[el2_lib.scala 197:80]
  wire  _T_154 = _T_150 | _T_153; // @[el2_lib.scala 197:25]
  wire  _T_156 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_157 = _T_156 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_160 = io_trigger_pkt_any_0_tdata2[14] == lsu_match_data_0[14]; // @[el2_lib.scala 197:80]
  wire  _T_161 = _T_157 | _T_160; // @[el2_lib.scala 197:25]
  wire  _T_163 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_164 = _T_163 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_167 = io_trigger_pkt_any_0_tdata2[15] == lsu_match_data_0[15]; // @[el2_lib.scala 197:80]
  wire  _T_168 = _T_164 | _T_167; // @[el2_lib.scala 197:25]
  wire  _T_170 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_171 = _T_170 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_174 = io_trigger_pkt_any_0_tdata2[16] == lsu_match_data_0[16]; // @[el2_lib.scala 197:80]
  wire  _T_175 = _T_171 | _T_174; // @[el2_lib.scala 197:25]
  wire  _T_177 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_178 = _T_177 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_181 = io_trigger_pkt_any_0_tdata2[17] == lsu_match_data_0[17]; // @[el2_lib.scala 197:80]
  wire  _T_182 = _T_178 | _T_181; // @[el2_lib.scala 197:25]
  wire  _T_184 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_185 = _T_184 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_188 = io_trigger_pkt_any_0_tdata2[18] == lsu_match_data_0[18]; // @[el2_lib.scala 197:80]
  wire  _T_189 = _T_185 | _T_188; // @[el2_lib.scala 197:25]
  wire  _T_191 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_192 = _T_191 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_195 = io_trigger_pkt_any_0_tdata2[19] == lsu_match_data_0[19]; // @[el2_lib.scala 197:80]
  wire  _T_196 = _T_192 | _T_195; // @[el2_lib.scala 197:25]
  wire  _T_198 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_199 = _T_198 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_202 = io_trigger_pkt_any_0_tdata2[20] == lsu_match_data_0[20]; // @[el2_lib.scala 197:80]
  wire  _T_203 = _T_199 | _T_202; // @[el2_lib.scala 197:25]
  wire  _T_205 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_206 = _T_205 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_209 = io_trigger_pkt_any_0_tdata2[21] == lsu_match_data_0[21]; // @[el2_lib.scala 197:80]
  wire  _T_210 = _T_206 | _T_209; // @[el2_lib.scala 197:25]
  wire  _T_212 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_213 = _T_212 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_216 = io_trigger_pkt_any_0_tdata2[22] == lsu_match_data_0[22]; // @[el2_lib.scala 197:80]
  wire  _T_217 = _T_213 | _T_216; // @[el2_lib.scala 197:25]
  wire  _T_219 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_220 = _T_219 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_223 = io_trigger_pkt_any_0_tdata2[23] == lsu_match_data_0[23]; // @[el2_lib.scala 197:80]
  wire  _T_224 = _T_220 | _T_223; // @[el2_lib.scala 197:25]
  wire  _T_226 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_227 = _T_226 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_230 = io_trigger_pkt_any_0_tdata2[24] == lsu_match_data_0[24]; // @[el2_lib.scala 197:80]
  wire  _T_231 = _T_227 | _T_230; // @[el2_lib.scala 197:25]
  wire  _T_233 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_234 = _T_233 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_237 = io_trigger_pkt_any_0_tdata2[25] == lsu_match_data_0[25]; // @[el2_lib.scala 197:80]
  wire  _T_238 = _T_234 | _T_237; // @[el2_lib.scala 197:25]
  wire  _T_240 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_241 = _T_240 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_244 = io_trigger_pkt_any_0_tdata2[26] == lsu_match_data_0[26]; // @[el2_lib.scala 197:80]
  wire  _T_245 = _T_241 | _T_244; // @[el2_lib.scala 197:25]
  wire  _T_247 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_248 = _T_247 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_251 = io_trigger_pkt_any_0_tdata2[27] == lsu_match_data_0[27]; // @[el2_lib.scala 197:80]
  wire  _T_252 = _T_248 | _T_251; // @[el2_lib.scala 197:25]
  wire  _T_254 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_255 = _T_254 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_258 = io_trigger_pkt_any_0_tdata2[28] == lsu_match_data_0[28]; // @[el2_lib.scala 197:80]
  wire  _T_259 = _T_255 | _T_258; // @[el2_lib.scala 197:25]
  wire  _T_261 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_262 = _T_261 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_265 = io_trigger_pkt_any_0_tdata2[29] == lsu_match_data_0[29]; // @[el2_lib.scala 197:80]
  wire  _T_266 = _T_262 | _T_265; // @[el2_lib.scala 197:25]
  wire  _T_268 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_269 = _T_268 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_272 = io_trigger_pkt_any_0_tdata2[30] == lsu_match_data_0[30]; // @[el2_lib.scala 197:80]
  wire  _T_273 = _T_269 | _T_272; // @[el2_lib.scala 197:25]
  wire  _T_275 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_276 = _T_275 & _T_59; // @[el2_lib.scala 197:43]
  wire  _T_279 = io_trigger_pkt_any_0_tdata2[31] == lsu_match_data_0[31]; // @[el2_lib.scala 197:80]
  wire  _T_280 = _T_276 | _T_279; // @[el2_lib.scala 197:25]
  wire [7:0] _T_287 = {_T_112,_T_105,_T_98,_T_91,_T_84,_T_77,_T_70,_T_63}; // @[el2_lib.scala 198:14]
  wire [15:0] _T_295 = {_T_168,_T_161,_T_154,_T_147,_T_140,_T_133,_T_126,_T_119,_T_287}; // @[el2_lib.scala 198:14]
  wire [7:0] _T_302 = {_T_224,_T_217,_T_210,_T_203,_T_196,_T_189,_T_182,_T_175}; // @[el2_lib.scala 198:14]
  wire [31:0] _T_311 = {_T_280,_T_273,_T_266,_T_259,_T_252,_T_245,_T_238,_T_231,_T_302,_T_295}; // @[el2_lib.scala 198:14]
  wire [31:0] _GEN_4 = {{31'd0}, _T_54}; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _T_312 = _GEN_4 & _T_311; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _GEN_5 = {{31'd0}, _T_51}; // @[el2_lsu_trigger.scala 21:141]
  wire [31:0] _T_313 = _GEN_5 | _T_312; // @[el2_lsu_trigger.scala 21:141]
  wire  _T_316 = io_trigger_pkt_any_1_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 21:120]
  wire  _T_317 = _T_49 & _T_316; // @[el2_lsu_trigger.scala 21:89]
  wire  _T_318 = io_trigger_pkt_any_1_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 22:33]
  wire  _T_320 = _T_318 & _T_20; // @[el2_lsu_trigger.scala 22:53]
  wire  _T_323 = &io_trigger_pkt_any_1_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_324 = ~_T_323; // @[el2_lib.scala 194:39]
  wire  _T_325 = io_trigger_pkt_any_1_match_ & _T_324; // @[el2_lib.scala 194:37]
  wire  _T_328 = io_trigger_pkt_any_1_tdata2[0] == lsu_match_data_1[0]; // @[el2_lib.scala 195:52]
  wire  _T_329 = _T_325 | _T_328; // @[el2_lib.scala 195:41]
  wire  _T_331 = &io_trigger_pkt_any_1_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_332 = _T_331 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_335 = io_trigger_pkt_any_1_tdata2[1] == lsu_match_data_1[1]; // @[el2_lib.scala 197:80]
  wire  _T_336 = _T_332 | _T_335; // @[el2_lib.scala 197:25]
  wire  _T_338 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_339 = _T_338 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_342 = io_trigger_pkt_any_1_tdata2[2] == lsu_match_data_1[2]; // @[el2_lib.scala 197:80]
  wire  _T_343 = _T_339 | _T_342; // @[el2_lib.scala 197:25]
  wire  _T_345 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_346 = _T_345 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_349 = io_trigger_pkt_any_1_tdata2[3] == lsu_match_data_1[3]; // @[el2_lib.scala 197:80]
  wire  _T_350 = _T_346 | _T_349; // @[el2_lib.scala 197:25]
  wire  _T_352 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_353 = _T_352 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_356 = io_trigger_pkt_any_1_tdata2[4] == lsu_match_data_1[4]; // @[el2_lib.scala 197:80]
  wire  _T_357 = _T_353 | _T_356; // @[el2_lib.scala 197:25]
  wire  _T_359 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_360 = _T_359 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_363 = io_trigger_pkt_any_1_tdata2[5] == lsu_match_data_1[5]; // @[el2_lib.scala 197:80]
  wire  _T_364 = _T_360 | _T_363; // @[el2_lib.scala 197:25]
  wire  _T_366 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_367 = _T_366 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_370 = io_trigger_pkt_any_1_tdata2[6] == lsu_match_data_1[6]; // @[el2_lib.scala 197:80]
  wire  _T_371 = _T_367 | _T_370; // @[el2_lib.scala 197:25]
  wire  _T_373 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_374 = _T_373 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_377 = io_trigger_pkt_any_1_tdata2[7] == lsu_match_data_1[7]; // @[el2_lib.scala 197:80]
  wire  _T_378 = _T_374 | _T_377; // @[el2_lib.scala 197:25]
  wire  _T_380 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_381 = _T_380 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_384 = io_trigger_pkt_any_1_tdata2[8] == lsu_match_data_1[8]; // @[el2_lib.scala 197:80]
  wire  _T_385 = _T_381 | _T_384; // @[el2_lib.scala 197:25]
  wire  _T_387 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_388 = _T_387 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_391 = io_trigger_pkt_any_1_tdata2[9] == lsu_match_data_1[9]; // @[el2_lib.scala 197:80]
  wire  _T_392 = _T_388 | _T_391; // @[el2_lib.scala 197:25]
  wire  _T_394 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_395 = _T_394 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_398 = io_trigger_pkt_any_1_tdata2[10] == lsu_match_data_1[10]; // @[el2_lib.scala 197:80]
  wire  _T_399 = _T_395 | _T_398; // @[el2_lib.scala 197:25]
  wire  _T_401 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_402 = _T_401 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_405 = io_trigger_pkt_any_1_tdata2[11] == lsu_match_data_1[11]; // @[el2_lib.scala 197:80]
  wire  _T_406 = _T_402 | _T_405; // @[el2_lib.scala 197:25]
  wire  _T_408 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_409 = _T_408 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_412 = io_trigger_pkt_any_1_tdata2[12] == lsu_match_data_1[12]; // @[el2_lib.scala 197:80]
  wire  _T_413 = _T_409 | _T_412; // @[el2_lib.scala 197:25]
  wire  _T_415 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_416 = _T_415 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_419 = io_trigger_pkt_any_1_tdata2[13] == lsu_match_data_1[13]; // @[el2_lib.scala 197:80]
  wire  _T_420 = _T_416 | _T_419; // @[el2_lib.scala 197:25]
  wire  _T_422 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_423 = _T_422 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_426 = io_trigger_pkt_any_1_tdata2[14] == lsu_match_data_1[14]; // @[el2_lib.scala 197:80]
  wire  _T_427 = _T_423 | _T_426; // @[el2_lib.scala 197:25]
  wire  _T_429 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_430 = _T_429 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_433 = io_trigger_pkt_any_1_tdata2[15] == lsu_match_data_1[15]; // @[el2_lib.scala 197:80]
  wire  _T_434 = _T_430 | _T_433; // @[el2_lib.scala 197:25]
  wire  _T_436 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_437 = _T_436 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_440 = io_trigger_pkt_any_1_tdata2[16] == lsu_match_data_1[16]; // @[el2_lib.scala 197:80]
  wire  _T_441 = _T_437 | _T_440; // @[el2_lib.scala 197:25]
  wire  _T_443 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_444 = _T_443 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_447 = io_trigger_pkt_any_1_tdata2[17] == lsu_match_data_1[17]; // @[el2_lib.scala 197:80]
  wire  _T_448 = _T_444 | _T_447; // @[el2_lib.scala 197:25]
  wire  _T_450 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_451 = _T_450 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_454 = io_trigger_pkt_any_1_tdata2[18] == lsu_match_data_1[18]; // @[el2_lib.scala 197:80]
  wire  _T_455 = _T_451 | _T_454; // @[el2_lib.scala 197:25]
  wire  _T_457 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_458 = _T_457 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_461 = io_trigger_pkt_any_1_tdata2[19] == lsu_match_data_1[19]; // @[el2_lib.scala 197:80]
  wire  _T_462 = _T_458 | _T_461; // @[el2_lib.scala 197:25]
  wire  _T_464 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_465 = _T_464 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_468 = io_trigger_pkt_any_1_tdata2[20] == lsu_match_data_1[20]; // @[el2_lib.scala 197:80]
  wire  _T_469 = _T_465 | _T_468; // @[el2_lib.scala 197:25]
  wire  _T_471 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_472 = _T_471 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_475 = io_trigger_pkt_any_1_tdata2[21] == lsu_match_data_1[21]; // @[el2_lib.scala 197:80]
  wire  _T_476 = _T_472 | _T_475; // @[el2_lib.scala 197:25]
  wire  _T_478 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_479 = _T_478 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_482 = io_trigger_pkt_any_1_tdata2[22] == lsu_match_data_1[22]; // @[el2_lib.scala 197:80]
  wire  _T_483 = _T_479 | _T_482; // @[el2_lib.scala 197:25]
  wire  _T_485 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_486 = _T_485 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_489 = io_trigger_pkt_any_1_tdata2[23] == lsu_match_data_1[23]; // @[el2_lib.scala 197:80]
  wire  _T_490 = _T_486 | _T_489; // @[el2_lib.scala 197:25]
  wire  _T_492 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_493 = _T_492 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_496 = io_trigger_pkt_any_1_tdata2[24] == lsu_match_data_1[24]; // @[el2_lib.scala 197:80]
  wire  _T_497 = _T_493 | _T_496; // @[el2_lib.scala 197:25]
  wire  _T_499 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_500 = _T_499 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_503 = io_trigger_pkt_any_1_tdata2[25] == lsu_match_data_1[25]; // @[el2_lib.scala 197:80]
  wire  _T_504 = _T_500 | _T_503; // @[el2_lib.scala 197:25]
  wire  _T_506 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_507 = _T_506 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_510 = io_trigger_pkt_any_1_tdata2[26] == lsu_match_data_1[26]; // @[el2_lib.scala 197:80]
  wire  _T_511 = _T_507 | _T_510; // @[el2_lib.scala 197:25]
  wire  _T_513 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_514 = _T_513 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_517 = io_trigger_pkt_any_1_tdata2[27] == lsu_match_data_1[27]; // @[el2_lib.scala 197:80]
  wire  _T_518 = _T_514 | _T_517; // @[el2_lib.scala 197:25]
  wire  _T_520 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_521 = _T_520 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_524 = io_trigger_pkt_any_1_tdata2[28] == lsu_match_data_1[28]; // @[el2_lib.scala 197:80]
  wire  _T_525 = _T_521 | _T_524; // @[el2_lib.scala 197:25]
  wire  _T_527 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_528 = _T_527 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_531 = io_trigger_pkt_any_1_tdata2[29] == lsu_match_data_1[29]; // @[el2_lib.scala 197:80]
  wire  _T_532 = _T_528 | _T_531; // @[el2_lib.scala 197:25]
  wire  _T_534 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_535 = _T_534 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_538 = io_trigger_pkt_any_1_tdata2[30] == lsu_match_data_1[30]; // @[el2_lib.scala 197:80]
  wire  _T_539 = _T_535 | _T_538; // @[el2_lib.scala 197:25]
  wire  _T_541 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_542 = _T_541 & _T_325; // @[el2_lib.scala 197:43]
  wire  _T_545 = io_trigger_pkt_any_1_tdata2[31] == lsu_match_data_1[31]; // @[el2_lib.scala 197:80]
  wire  _T_546 = _T_542 | _T_545; // @[el2_lib.scala 197:25]
  wire [7:0] _T_553 = {_T_378,_T_371,_T_364,_T_357,_T_350,_T_343,_T_336,_T_329}; // @[el2_lib.scala 198:14]
  wire [15:0] _T_561 = {_T_434,_T_427,_T_420,_T_413,_T_406,_T_399,_T_392,_T_385,_T_553}; // @[el2_lib.scala 198:14]
  wire [7:0] _T_568 = {_T_490,_T_483,_T_476,_T_469,_T_462,_T_455,_T_448,_T_441}; // @[el2_lib.scala 198:14]
  wire [31:0] _T_577 = {_T_546,_T_539,_T_532,_T_525,_T_518,_T_511,_T_504,_T_497,_T_568,_T_561}; // @[el2_lib.scala 198:14]
  wire [31:0] _GEN_6 = {{31'd0}, _T_320}; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _T_578 = _GEN_6 & _T_577; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _GEN_7 = {{31'd0}, _T_317}; // @[el2_lsu_trigger.scala 21:141]
  wire [31:0] _T_579 = _GEN_7 | _T_578; // @[el2_lsu_trigger.scala 21:141]
  wire  _T_582 = io_trigger_pkt_any_2_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 21:120]
  wire  _T_583 = _T_49 & _T_582; // @[el2_lsu_trigger.scala 21:89]
  wire  _T_584 = io_trigger_pkt_any_2_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 22:33]
  wire  _T_586 = _T_584 & _T_29; // @[el2_lsu_trigger.scala 22:53]
  wire  _T_589 = &io_trigger_pkt_any_2_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_590 = ~_T_589; // @[el2_lib.scala 194:39]
  wire  _T_591 = io_trigger_pkt_any_2_match_ & _T_590; // @[el2_lib.scala 194:37]
  wire  _T_594 = io_trigger_pkt_any_2_tdata2[0] == lsu_match_data_2[0]; // @[el2_lib.scala 195:52]
  wire  _T_595 = _T_591 | _T_594; // @[el2_lib.scala 195:41]
  wire  _T_597 = &io_trigger_pkt_any_2_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_598 = _T_597 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_601 = io_trigger_pkt_any_2_tdata2[1] == lsu_match_data_2[1]; // @[el2_lib.scala 197:80]
  wire  _T_602 = _T_598 | _T_601; // @[el2_lib.scala 197:25]
  wire  _T_604 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_605 = _T_604 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_608 = io_trigger_pkt_any_2_tdata2[2] == lsu_match_data_2[2]; // @[el2_lib.scala 197:80]
  wire  _T_609 = _T_605 | _T_608; // @[el2_lib.scala 197:25]
  wire  _T_611 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_612 = _T_611 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_615 = io_trigger_pkt_any_2_tdata2[3] == lsu_match_data_2[3]; // @[el2_lib.scala 197:80]
  wire  _T_616 = _T_612 | _T_615; // @[el2_lib.scala 197:25]
  wire  _T_618 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_619 = _T_618 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_622 = io_trigger_pkt_any_2_tdata2[4] == lsu_match_data_2[4]; // @[el2_lib.scala 197:80]
  wire  _T_623 = _T_619 | _T_622; // @[el2_lib.scala 197:25]
  wire  _T_625 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_626 = _T_625 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_629 = io_trigger_pkt_any_2_tdata2[5] == lsu_match_data_2[5]; // @[el2_lib.scala 197:80]
  wire  _T_630 = _T_626 | _T_629; // @[el2_lib.scala 197:25]
  wire  _T_632 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_633 = _T_632 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_636 = io_trigger_pkt_any_2_tdata2[6] == lsu_match_data_2[6]; // @[el2_lib.scala 197:80]
  wire  _T_637 = _T_633 | _T_636; // @[el2_lib.scala 197:25]
  wire  _T_639 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_640 = _T_639 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_643 = io_trigger_pkt_any_2_tdata2[7] == lsu_match_data_2[7]; // @[el2_lib.scala 197:80]
  wire  _T_644 = _T_640 | _T_643; // @[el2_lib.scala 197:25]
  wire  _T_646 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_647 = _T_646 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_650 = io_trigger_pkt_any_2_tdata2[8] == lsu_match_data_2[8]; // @[el2_lib.scala 197:80]
  wire  _T_651 = _T_647 | _T_650; // @[el2_lib.scala 197:25]
  wire  _T_653 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_654 = _T_653 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_657 = io_trigger_pkt_any_2_tdata2[9] == lsu_match_data_2[9]; // @[el2_lib.scala 197:80]
  wire  _T_658 = _T_654 | _T_657; // @[el2_lib.scala 197:25]
  wire  _T_660 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_661 = _T_660 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_664 = io_trigger_pkt_any_2_tdata2[10] == lsu_match_data_2[10]; // @[el2_lib.scala 197:80]
  wire  _T_665 = _T_661 | _T_664; // @[el2_lib.scala 197:25]
  wire  _T_667 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_668 = _T_667 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_671 = io_trigger_pkt_any_2_tdata2[11] == lsu_match_data_2[11]; // @[el2_lib.scala 197:80]
  wire  _T_672 = _T_668 | _T_671; // @[el2_lib.scala 197:25]
  wire  _T_674 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_675 = _T_674 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_678 = io_trigger_pkt_any_2_tdata2[12] == lsu_match_data_2[12]; // @[el2_lib.scala 197:80]
  wire  _T_679 = _T_675 | _T_678; // @[el2_lib.scala 197:25]
  wire  _T_681 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_682 = _T_681 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_685 = io_trigger_pkt_any_2_tdata2[13] == lsu_match_data_2[13]; // @[el2_lib.scala 197:80]
  wire  _T_686 = _T_682 | _T_685; // @[el2_lib.scala 197:25]
  wire  _T_688 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_689 = _T_688 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_692 = io_trigger_pkt_any_2_tdata2[14] == lsu_match_data_2[14]; // @[el2_lib.scala 197:80]
  wire  _T_693 = _T_689 | _T_692; // @[el2_lib.scala 197:25]
  wire  _T_695 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_696 = _T_695 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_699 = io_trigger_pkt_any_2_tdata2[15] == lsu_match_data_2[15]; // @[el2_lib.scala 197:80]
  wire  _T_700 = _T_696 | _T_699; // @[el2_lib.scala 197:25]
  wire  _T_702 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_703 = _T_702 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_706 = io_trigger_pkt_any_2_tdata2[16] == lsu_match_data_2[16]; // @[el2_lib.scala 197:80]
  wire  _T_707 = _T_703 | _T_706; // @[el2_lib.scala 197:25]
  wire  _T_709 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_710 = _T_709 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_713 = io_trigger_pkt_any_2_tdata2[17] == lsu_match_data_2[17]; // @[el2_lib.scala 197:80]
  wire  _T_714 = _T_710 | _T_713; // @[el2_lib.scala 197:25]
  wire  _T_716 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_717 = _T_716 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_720 = io_trigger_pkt_any_2_tdata2[18] == lsu_match_data_2[18]; // @[el2_lib.scala 197:80]
  wire  _T_721 = _T_717 | _T_720; // @[el2_lib.scala 197:25]
  wire  _T_723 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_724 = _T_723 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_727 = io_trigger_pkt_any_2_tdata2[19] == lsu_match_data_2[19]; // @[el2_lib.scala 197:80]
  wire  _T_728 = _T_724 | _T_727; // @[el2_lib.scala 197:25]
  wire  _T_730 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_731 = _T_730 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_734 = io_trigger_pkt_any_2_tdata2[20] == lsu_match_data_2[20]; // @[el2_lib.scala 197:80]
  wire  _T_735 = _T_731 | _T_734; // @[el2_lib.scala 197:25]
  wire  _T_737 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_738 = _T_737 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_741 = io_trigger_pkt_any_2_tdata2[21] == lsu_match_data_2[21]; // @[el2_lib.scala 197:80]
  wire  _T_742 = _T_738 | _T_741; // @[el2_lib.scala 197:25]
  wire  _T_744 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_745 = _T_744 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_748 = io_trigger_pkt_any_2_tdata2[22] == lsu_match_data_2[22]; // @[el2_lib.scala 197:80]
  wire  _T_749 = _T_745 | _T_748; // @[el2_lib.scala 197:25]
  wire  _T_751 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_752 = _T_751 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_755 = io_trigger_pkt_any_2_tdata2[23] == lsu_match_data_2[23]; // @[el2_lib.scala 197:80]
  wire  _T_756 = _T_752 | _T_755; // @[el2_lib.scala 197:25]
  wire  _T_758 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_759 = _T_758 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_762 = io_trigger_pkt_any_2_tdata2[24] == lsu_match_data_2[24]; // @[el2_lib.scala 197:80]
  wire  _T_763 = _T_759 | _T_762; // @[el2_lib.scala 197:25]
  wire  _T_765 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_766 = _T_765 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_769 = io_trigger_pkt_any_2_tdata2[25] == lsu_match_data_2[25]; // @[el2_lib.scala 197:80]
  wire  _T_770 = _T_766 | _T_769; // @[el2_lib.scala 197:25]
  wire  _T_772 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_773 = _T_772 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_776 = io_trigger_pkt_any_2_tdata2[26] == lsu_match_data_2[26]; // @[el2_lib.scala 197:80]
  wire  _T_777 = _T_773 | _T_776; // @[el2_lib.scala 197:25]
  wire  _T_779 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_780 = _T_779 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_783 = io_trigger_pkt_any_2_tdata2[27] == lsu_match_data_2[27]; // @[el2_lib.scala 197:80]
  wire  _T_784 = _T_780 | _T_783; // @[el2_lib.scala 197:25]
  wire  _T_786 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_787 = _T_786 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_790 = io_trigger_pkt_any_2_tdata2[28] == lsu_match_data_2[28]; // @[el2_lib.scala 197:80]
  wire  _T_791 = _T_787 | _T_790; // @[el2_lib.scala 197:25]
  wire  _T_793 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_794 = _T_793 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_797 = io_trigger_pkt_any_2_tdata2[29] == lsu_match_data_2[29]; // @[el2_lib.scala 197:80]
  wire  _T_798 = _T_794 | _T_797; // @[el2_lib.scala 197:25]
  wire  _T_800 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_801 = _T_800 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_804 = io_trigger_pkt_any_2_tdata2[30] == lsu_match_data_2[30]; // @[el2_lib.scala 197:80]
  wire  _T_805 = _T_801 | _T_804; // @[el2_lib.scala 197:25]
  wire  _T_807 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_808 = _T_807 & _T_591; // @[el2_lib.scala 197:43]
  wire  _T_811 = io_trigger_pkt_any_2_tdata2[31] == lsu_match_data_2[31]; // @[el2_lib.scala 197:80]
  wire  _T_812 = _T_808 | _T_811; // @[el2_lib.scala 197:25]
  wire [7:0] _T_819 = {_T_644,_T_637,_T_630,_T_623,_T_616,_T_609,_T_602,_T_595}; // @[el2_lib.scala 198:14]
  wire [15:0] _T_827 = {_T_700,_T_693,_T_686,_T_679,_T_672,_T_665,_T_658,_T_651,_T_819}; // @[el2_lib.scala 198:14]
  wire [7:0] _T_834 = {_T_756,_T_749,_T_742,_T_735,_T_728,_T_721,_T_714,_T_707}; // @[el2_lib.scala 198:14]
  wire [31:0] _T_843 = {_T_812,_T_805,_T_798,_T_791,_T_784,_T_777,_T_770,_T_763,_T_834,_T_827}; // @[el2_lib.scala 198:14]
  wire [31:0] _GEN_8 = {{31'd0}, _T_586}; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _T_844 = _GEN_8 & _T_843; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _GEN_9 = {{31'd0}, _T_583}; // @[el2_lsu_trigger.scala 21:141]
  wire [31:0] _T_845 = _GEN_9 | _T_844; // @[el2_lsu_trigger.scala 21:141]
  wire  _T_848 = io_trigger_pkt_any_3_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 21:120]
  wire  _T_849 = _T_49 & _T_848; // @[el2_lsu_trigger.scala 21:89]
  wire  _T_850 = io_trigger_pkt_any_3_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 22:33]
  wire  _T_852 = _T_850 & _T_38; // @[el2_lsu_trigger.scala 22:53]
  wire  _T_855 = &io_trigger_pkt_any_3_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_856 = ~_T_855; // @[el2_lib.scala 194:39]
  wire  _T_857 = io_trigger_pkt_any_3_match_ & _T_856; // @[el2_lib.scala 194:37]
  wire  _T_860 = io_trigger_pkt_any_3_tdata2[0] == lsu_match_data_3[0]; // @[el2_lib.scala 195:52]
  wire  _T_861 = _T_857 | _T_860; // @[el2_lib.scala 195:41]
  wire  _T_863 = &io_trigger_pkt_any_3_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_864 = _T_863 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_867 = io_trigger_pkt_any_3_tdata2[1] == lsu_match_data_3[1]; // @[el2_lib.scala 197:80]
  wire  _T_868 = _T_864 | _T_867; // @[el2_lib.scala 197:25]
  wire  _T_870 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_871 = _T_870 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_874 = io_trigger_pkt_any_3_tdata2[2] == lsu_match_data_3[2]; // @[el2_lib.scala 197:80]
  wire  _T_875 = _T_871 | _T_874; // @[el2_lib.scala 197:25]
  wire  _T_877 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_878 = _T_877 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_881 = io_trigger_pkt_any_3_tdata2[3] == lsu_match_data_3[3]; // @[el2_lib.scala 197:80]
  wire  _T_882 = _T_878 | _T_881; // @[el2_lib.scala 197:25]
  wire  _T_884 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_885 = _T_884 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_888 = io_trigger_pkt_any_3_tdata2[4] == lsu_match_data_3[4]; // @[el2_lib.scala 197:80]
  wire  _T_889 = _T_885 | _T_888; // @[el2_lib.scala 197:25]
  wire  _T_891 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_892 = _T_891 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_895 = io_trigger_pkt_any_3_tdata2[5] == lsu_match_data_3[5]; // @[el2_lib.scala 197:80]
  wire  _T_896 = _T_892 | _T_895; // @[el2_lib.scala 197:25]
  wire  _T_898 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_899 = _T_898 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_902 = io_trigger_pkt_any_3_tdata2[6] == lsu_match_data_3[6]; // @[el2_lib.scala 197:80]
  wire  _T_903 = _T_899 | _T_902; // @[el2_lib.scala 197:25]
  wire  _T_905 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_906 = _T_905 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_909 = io_trigger_pkt_any_3_tdata2[7] == lsu_match_data_3[7]; // @[el2_lib.scala 197:80]
  wire  _T_910 = _T_906 | _T_909; // @[el2_lib.scala 197:25]
  wire  _T_912 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_913 = _T_912 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_916 = io_trigger_pkt_any_3_tdata2[8] == lsu_match_data_3[8]; // @[el2_lib.scala 197:80]
  wire  _T_917 = _T_913 | _T_916; // @[el2_lib.scala 197:25]
  wire  _T_919 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_920 = _T_919 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_923 = io_trigger_pkt_any_3_tdata2[9] == lsu_match_data_3[9]; // @[el2_lib.scala 197:80]
  wire  _T_924 = _T_920 | _T_923; // @[el2_lib.scala 197:25]
  wire  _T_926 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_927 = _T_926 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_930 = io_trigger_pkt_any_3_tdata2[10] == lsu_match_data_3[10]; // @[el2_lib.scala 197:80]
  wire  _T_931 = _T_927 | _T_930; // @[el2_lib.scala 197:25]
  wire  _T_933 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_934 = _T_933 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_937 = io_trigger_pkt_any_3_tdata2[11] == lsu_match_data_3[11]; // @[el2_lib.scala 197:80]
  wire  _T_938 = _T_934 | _T_937; // @[el2_lib.scala 197:25]
  wire  _T_940 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_941 = _T_940 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_944 = io_trigger_pkt_any_3_tdata2[12] == lsu_match_data_3[12]; // @[el2_lib.scala 197:80]
  wire  _T_945 = _T_941 | _T_944; // @[el2_lib.scala 197:25]
  wire  _T_947 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_948 = _T_947 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_951 = io_trigger_pkt_any_3_tdata2[13] == lsu_match_data_3[13]; // @[el2_lib.scala 197:80]
  wire  _T_952 = _T_948 | _T_951; // @[el2_lib.scala 197:25]
  wire  _T_954 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_955 = _T_954 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_958 = io_trigger_pkt_any_3_tdata2[14] == lsu_match_data_3[14]; // @[el2_lib.scala 197:80]
  wire  _T_959 = _T_955 | _T_958; // @[el2_lib.scala 197:25]
  wire  _T_961 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_962 = _T_961 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_965 = io_trigger_pkt_any_3_tdata2[15] == lsu_match_data_3[15]; // @[el2_lib.scala 197:80]
  wire  _T_966 = _T_962 | _T_965; // @[el2_lib.scala 197:25]
  wire  _T_968 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_969 = _T_968 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_972 = io_trigger_pkt_any_3_tdata2[16] == lsu_match_data_3[16]; // @[el2_lib.scala 197:80]
  wire  _T_973 = _T_969 | _T_972; // @[el2_lib.scala 197:25]
  wire  _T_975 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_976 = _T_975 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_979 = io_trigger_pkt_any_3_tdata2[17] == lsu_match_data_3[17]; // @[el2_lib.scala 197:80]
  wire  _T_980 = _T_976 | _T_979; // @[el2_lib.scala 197:25]
  wire  _T_982 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_983 = _T_982 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_986 = io_trigger_pkt_any_3_tdata2[18] == lsu_match_data_3[18]; // @[el2_lib.scala 197:80]
  wire  _T_987 = _T_983 | _T_986; // @[el2_lib.scala 197:25]
  wire  _T_989 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_990 = _T_989 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_993 = io_trigger_pkt_any_3_tdata2[19] == lsu_match_data_3[19]; // @[el2_lib.scala 197:80]
  wire  _T_994 = _T_990 | _T_993; // @[el2_lib.scala 197:25]
  wire  _T_996 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_997 = _T_996 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1000 = io_trigger_pkt_any_3_tdata2[20] == lsu_match_data_3[20]; // @[el2_lib.scala 197:80]
  wire  _T_1001 = _T_997 | _T_1000; // @[el2_lib.scala 197:25]
  wire  _T_1003 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_1004 = _T_1003 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1007 = io_trigger_pkt_any_3_tdata2[21] == lsu_match_data_3[21]; // @[el2_lib.scala 197:80]
  wire  _T_1008 = _T_1004 | _T_1007; // @[el2_lib.scala 197:25]
  wire  _T_1010 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_1011 = _T_1010 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1014 = io_trigger_pkt_any_3_tdata2[22] == lsu_match_data_3[22]; // @[el2_lib.scala 197:80]
  wire  _T_1015 = _T_1011 | _T_1014; // @[el2_lib.scala 197:25]
  wire  _T_1017 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_1018 = _T_1017 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1021 = io_trigger_pkt_any_3_tdata2[23] == lsu_match_data_3[23]; // @[el2_lib.scala 197:80]
  wire  _T_1022 = _T_1018 | _T_1021; // @[el2_lib.scala 197:25]
  wire  _T_1024 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_1025 = _T_1024 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1028 = io_trigger_pkt_any_3_tdata2[24] == lsu_match_data_3[24]; // @[el2_lib.scala 197:80]
  wire  _T_1029 = _T_1025 | _T_1028; // @[el2_lib.scala 197:25]
  wire  _T_1031 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_1032 = _T_1031 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1035 = io_trigger_pkt_any_3_tdata2[25] == lsu_match_data_3[25]; // @[el2_lib.scala 197:80]
  wire  _T_1036 = _T_1032 | _T_1035; // @[el2_lib.scala 197:25]
  wire  _T_1038 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_1039 = _T_1038 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1042 = io_trigger_pkt_any_3_tdata2[26] == lsu_match_data_3[26]; // @[el2_lib.scala 197:80]
  wire  _T_1043 = _T_1039 | _T_1042; // @[el2_lib.scala 197:25]
  wire  _T_1045 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_1046 = _T_1045 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1049 = io_trigger_pkt_any_3_tdata2[27] == lsu_match_data_3[27]; // @[el2_lib.scala 197:80]
  wire  _T_1050 = _T_1046 | _T_1049; // @[el2_lib.scala 197:25]
  wire  _T_1052 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_1053 = _T_1052 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1056 = io_trigger_pkt_any_3_tdata2[28] == lsu_match_data_3[28]; // @[el2_lib.scala 197:80]
  wire  _T_1057 = _T_1053 | _T_1056; // @[el2_lib.scala 197:25]
  wire  _T_1059 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_1060 = _T_1059 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1063 = io_trigger_pkt_any_3_tdata2[29] == lsu_match_data_3[29]; // @[el2_lib.scala 197:80]
  wire  _T_1064 = _T_1060 | _T_1063; // @[el2_lib.scala 197:25]
  wire  _T_1066 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_1067 = _T_1066 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1070 = io_trigger_pkt_any_3_tdata2[30] == lsu_match_data_3[30]; // @[el2_lib.scala 197:80]
  wire  _T_1071 = _T_1067 | _T_1070; // @[el2_lib.scala 197:25]
  wire  _T_1073 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_1074 = _T_1073 & _T_857; // @[el2_lib.scala 197:43]
  wire  _T_1077 = io_trigger_pkt_any_3_tdata2[31] == lsu_match_data_3[31]; // @[el2_lib.scala 197:80]
  wire  _T_1078 = _T_1074 | _T_1077; // @[el2_lib.scala 197:25]
  wire [7:0] _T_1085 = {_T_910,_T_903,_T_896,_T_889,_T_882,_T_875,_T_868,_T_861}; // @[el2_lib.scala 198:14]
  wire [15:0] _T_1093 = {_T_966,_T_959,_T_952,_T_945,_T_938,_T_931,_T_924,_T_917,_T_1085}; // @[el2_lib.scala 198:14]
  wire [7:0] _T_1100 = {_T_1022,_T_1015,_T_1008,_T_1001,_T_994,_T_987,_T_980,_T_973}; // @[el2_lib.scala 198:14]
  wire [31:0] _T_1109 = {_T_1078,_T_1071,_T_1064,_T_1057,_T_1050,_T_1043,_T_1036,_T_1029,_T_1100,_T_1093}; // @[el2_lib.scala 198:14]
  wire [31:0] _GEN_10 = {{31'd0}, _T_852}; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _T_1110 = _GEN_10 & _T_1109; // @[el2_lsu_trigger.scala 22:86]
  wire [31:0] _GEN_11 = {{31'd0}, _T_849}; // @[el2_lsu_trigger.scala 21:141]
  wire [31:0] _T_1111 = _GEN_11 | _T_1110; // @[el2_lsu_trigger.scala 21:141]
  wire [127:0] _T_1114 = {_T_1111,_T_845,_T_579,_T_313}; // @[Cat.scala 29:58]
  assign io_lsu_trigger_match_m = _T_1114[3:0]; // @[el2_lsu_trigger.scala 16:25 el2_lsu_trigger.scala 21:26]
endmodule
