module el2_ifu_compress_ctl(
  input         clock,
  input         reset,
  input  [15:0] io_din,
  output [31:0] io_dout,
  output [31:0] io_l1,
  output [31:0] io_l2,
  output [31:0] io_l3,
  output        io_legal,
  output [31:0] io_o,
  output [19:0] io_sluimmd,
  output [5:0]  io_uimm5d,
  output [5:0]  io_ulwspimm7d,
  output [4:0]  io_ulwimm6d,
  output [5:0]  io_simm9d,
  output [7:0]  io_uimm9d,
  output [5:0]  io_simm5d,
  output [19:0] io_sjald,
  output [11:0] io_l2_31
);
  wire  _T_2 = ~io_din[14]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_4 = ~io_din[13]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_7 = ~io_din[6]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_9 = ~io_din[5]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_11 = io_din[15] & _T_2; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_12 = _T_11 & _T_4; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_13 = _T_12 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_14 = _T_13 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_15 = _T_14 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_16 = _T_15 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_23 = ~io_din[11]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_28 = _T_12 & _T_23; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_29 = _T_28 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_30 = _T_29 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  out_30 = _T_16 | _T_30; // @[el2_ifu_compress_ctl.scala 32:53]
  wire  _T_38 = ~io_din[10]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_40 = ~io_din[9]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_42 = ~io_din[8]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_44 = ~io_din[7]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_50 = ~io_din[4]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_52 = ~io_din[3]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_54 = ~io_din[2]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_56 = _T_2 & io_din[12]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_57 = _T_56 & _T_23; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_58 = _T_57 & _T_38; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_59 = _T_58 & _T_40; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_60 = _T_59 & _T_42; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_61 = _T_60 & _T_44; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_62 = _T_61 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_63 = _T_62 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_64 = _T_63 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_65 = _T_64 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_66 = _T_65 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  out_20 = _T_66 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_79 = _T_28 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_90 = _T_12 & _T_38; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_91 = _T_90 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_92 = _T_79 | _T_91; // @[el2_ifu_compress_ctl.scala 34:46]
  wire  _T_102 = _T_12 & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_103 = _T_102 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_104 = _T_92 | _T_103; // @[el2_ifu_compress_ctl.scala 34:80]
  wire  _T_114 = _T_12 & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_115 = _T_114 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  out_14 = _T_104 | _T_115; // @[el2_ifu_compress_ctl.scala 34:113]
  wire  _T_128 = _T_12 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_129 = _T_128 & _T_38; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_130 = _T_129 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_142 = _T_128 & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_143 = _T_142 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_144 = _T_130 | _T_143; // @[el2_ifu_compress_ctl.scala 36:50]
  wire  _T_147 = ~io_din[0]; // @[el2_ifu_compress_ctl.scala 36:101]
  wire  _T_148 = io_din[14] & _T_147; // @[el2_ifu_compress_ctl.scala 36:99]
  wire  out_13 = _T_144 | _T_148; // @[el2_ifu_compress_ctl.scala 36:86]
  wire  _T_161 = _T_102 & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_162 = _T_161 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_175 = _T_162 | _T_79; // @[el2_ifu_compress_ctl.scala 37:47]
  wire  _T_188 = _T_175 | _T_91; // @[el2_ifu_compress_ctl.scala 37:81]
  wire  _T_190 = ~io_din[15]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_194 = _T_190 & _T_2; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_195 = _T_194 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_196 = _T_188 | _T_195; // @[el2_ifu_compress_ctl.scala 37:115]
  wire  _T_200 = io_din[15] & io_din[14]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_201 = _T_200 & io_din[13]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  out_12 = _T_196 | _T_201; // @[el2_ifu_compress_ctl.scala 38:26]
  wire  _T_217 = _T_11 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_218 = _T_217 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_219 = _T_218 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_220 = _T_219 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_221 = _T_220 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_224 = _T_221 & _T_147; // @[el2_ifu_compress_ctl.scala 39:53]
  wire  _T_228 = _T_2 & io_din[13]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_229 = _T_224 | _T_228; // @[el2_ifu_compress_ctl.scala 39:67]
  wire  _T_234 = _T_200 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  out_6 = _T_229 | _T_234; // @[el2_ifu_compress_ctl.scala 39:88]
  wire  _T_239 = io_din[15] & _T_147; // @[el2_ifu_compress_ctl.scala 41:24]
  wire  _T_243 = io_din[15] & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_244 = _T_243 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_245 = _T_239 | _T_244; // @[el2_ifu_compress_ctl.scala 41:39]
  wire  _T_249 = io_din[13] & _T_42; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_250 = _T_245 | _T_249; // @[el2_ifu_compress_ctl.scala 41:63]
  wire  _T_253 = io_din[13] & io_din[7]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_254 = _T_250 | _T_253; // @[el2_ifu_compress_ctl.scala 41:83]
  wire  _T_257 = io_din[13] & io_din[9]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_258 = _T_254 | _T_257; // @[el2_ifu_compress_ctl.scala 41:102]
  wire  _T_261 = io_din[13] & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_262 = _T_258 | _T_261; // @[el2_ifu_compress_ctl.scala 42:22]
  wire  _T_265 = io_din[13] & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_266 = _T_262 | _T_265; // @[el2_ifu_compress_ctl.scala 42:42]
  wire  _T_271 = _T_266 | _T_228; // @[el2_ifu_compress_ctl.scala 42:62]
  wire  out_5 = _T_271 | _T_200; // @[el2_ifu_compress_ctl.scala 42:83]
  wire  _T_288 = _T_2 & _T_23; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_289 = _T_288 & _T_38; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_290 = _T_289 & _T_40; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_291 = _T_290 & _T_42; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_292 = _T_291 & _T_44; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_295 = _T_292 & _T_147; // @[el2_ifu_compress_ctl.scala 45:50]
  wire  _T_303 = _T_194 & _T_147; // @[el2_ifu_compress_ctl.scala 45:87]
  wire  _T_304 = _T_295 | _T_303; // @[el2_ifu_compress_ctl.scala 45:65]
  wire  _T_308 = _T_2 & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_311 = _T_308 & _T_147; // @[el2_ifu_compress_ctl.scala 46:23]
  wire  _T_312 = _T_304 | _T_311; // @[el2_ifu_compress_ctl.scala 45:102]
  wire  _T_317 = _T_190 & io_din[14]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_318 = _T_317 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_319 = _T_312 | _T_318; // @[el2_ifu_compress_ctl.scala 46:38]
  wire  _T_323 = _T_2 & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_326 = _T_323 & _T_147; // @[el2_ifu_compress_ctl.scala 46:82]
  wire  _T_327 = _T_319 | _T_326; // @[el2_ifu_compress_ctl.scala 46:62]
  wire  _T_331 = _T_2 & io_din[4]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_334 = _T_331 & _T_147; // @[el2_ifu_compress_ctl.scala 47:23]
  wire  _T_335 = _T_327 | _T_334; // @[el2_ifu_compress_ctl.scala 46:97]
  wire  _T_339 = _T_2 & io_din[3]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_342 = _T_339 & _T_147; // @[el2_ifu_compress_ctl.scala 47:58]
  wire  _T_343 = _T_335 | _T_342; // @[el2_ifu_compress_ctl.scala 47:38]
  wire  _T_347 = _T_2 & io_din[2]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_350 = _T_347 & _T_147; // @[el2_ifu_compress_ctl.scala 47:93]
  wire  _T_351 = _T_343 | _T_350; // @[el2_ifu_compress_ctl.scala 47:73]
  wire  _T_357 = _T_2 & _T_4; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_358 = _T_357 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  out_4 = _T_351 | _T_358; // @[el2_ifu_compress_ctl.scala 47:108]
  wire  _T_380 = _T_56 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_381 = _T_380 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_382 = _T_381 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_383 = _T_382 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_384 = _T_383 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_385 = _T_384 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_386 = _T_385 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_403 = _T_56 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_404 = _T_403 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_405 = _T_404 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_406 = _T_405 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_407 = _T_406 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_408 = _T_407 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_409 = _T_408 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_410 = _T_386 | _T_409; // @[el2_ifu_compress_ctl.scala 54:59]
  wire  _T_427 = _T_56 & io_din[9]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_428 = _T_427 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_429 = _T_428 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_430 = _T_429 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_431 = _T_430 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_432 = _T_431 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_433 = _T_432 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_434 = _T_410 | _T_433; // @[el2_ifu_compress_ctl.scala 55:59]
  wire  _T_451 = _T_56 & io_din[8]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_452 = _T_451 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_453 = _T_452 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_454 = _T_453 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_455 = _T_454 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_456 = _T_455 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_457 = _T_456 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_458 = _T_434 | _T_457; // @[el2_ifu_compress_ctl.scala 56:58]
  wire  _T_475 = _T_56 & io_din[7]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_476 = _T_475 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_477 = _T_476 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_478 = _T_477 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_479 = _T_478 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_480 = _T_479 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_481 = _T_480 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_482 = _T_458 | _T_481; // @[el2_ifu_compress_ctl.scala 57:55]
  wire  _T_487 = ~io_din[12]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_499 = _T_11 & _T_487; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_500 = _T_499 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_501 = _T_500 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_502 = _T_501 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_503 = _T_502 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_504 = _T_503 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_507 = _T_504 & _T_147; // @[el2_ifu_compress_ctl.scala 59:56]
  wire  _T_508 = _T_482 | _T_507; // @[el2_ifu_compress_ctl.scala 58:57]
  wire  _T_514 = _T_190 & io_din[13]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_515 = _T_514 & _T_42; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_516 = _T_508 | _T_515; // @[el2_ifu_compress_ctl.scala 59:71]
  wire  _T_522 = _T_514 & io_din[7]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_523 = _T_516 | _T_522; // @[el2_ifu_compress_ctl.scala 60:34]
  wire  _T_529 = _T_514 & io_din[9]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_530 = _T_523 | _T_529; // @[el2_ifu_compress_ctl.scala 61:33]
  wire  _T_536 = _T_514 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_537 = _T_530 | _T_536; // @[el2_ifu_compress_ctl.scala 62:33]
  wire  _T_543 = _T_514 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_544 = _T_537 | _T_543; // @[el2_ifu_compress_ctl.scala 63:34]
  wire  out_2 = _T_544 | _T_228; // @[el2_ifu_compress_ctl.scala 64:34]
  wire [4:0] rs2d = io_din[6:2]; // @[el2_ifu_compress_ctl.scala 73:20]
  wire [4:0] rdd = io_din[11:7]; // @[el2_ifu_compress_ctl.scala 74:19]
  wire [4:0] rdpd = {2'h1,io_din[9:7]}; // @[Cat.scala 29:58]
  wire [4:0] rs2pd = {2'h1,io_din[4:2]}; // @[Cat.scala 29:58]
  wire  _T_557 = _T_308 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_564 = _T_317 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_565 = _T_564 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_566 = _T_557 | _T_565; // @[el2_ifu_compress_ctl.scala 78:33]
  wire  _T_572 = _T_323 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_573 = _T_566 | _T_572; // @[el2_ifu_compress_ctl.scala 78:58]
  wire  _T_580 = _T_317 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_581 = _T_580 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_582 = _T_573 | _T_581; // @[el2_ifu_compress_ctl.scala 78:79]
  wire  _T_588 = _T_331 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_589 = _T_582 | _T_588; // @[el2_ifu_compress_ctl.scala 78:104]
  wire  _T_596 = _T_317 & io_din[9]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_597 = _T_596 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_598 = _T_589 | _T_597; // @[el2_ifu_compress_ctl.scala 79:24]
  wire  _T_604 = _T_339 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_605 = _T_598 | _T_604; // @[el2_ifu_compress_ctl.scala 79:48]
  wire  _T_613 = _T_317 & _T_42; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_614 = _T_613 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_615 = _T_605 | _T_614; // @[el2_ifu_compress_ctl.scala 79:69]
  wire  _T_621 = _T_347 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_622 = _T_615 | _T_621; // @[el2_ifu_compress_ctl.scala 79:94]
  wire  _T_629 = _T_317 & io_din[7]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_630 = _T_629 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_631 = _T_622 | _T_630; // @[el2_ifu_compress_ctl.scala 80:22]
  wire  _T_635 = _T_190 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_636 = _T_631 | _T_635; // @[el2_ifu_compress_ctl.scala 80:46]
  wire  _T_642 = _T_190 & _T_4; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_643 = _T_642 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  rdrd = _T_636 | _T_643; // @[el2_ifu_compress_ctl.scala 80:65]
  wire  _T_651 = _T_380 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_659 = _T_403 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_660 = _T_651 | _T_659; // @[el2_ifu_compress_ctl.scala 82:38]
  wire  _T_668 = _T_427 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_669 = _T_660 | _T_668; // @[el2_ifu_compress_ctl.scala 83:28]
  wire  _T_677 = _T_451 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_678 = _T_669 | _T_677; // @[el2_ifu_compress_ctl.scala 84:27]
  wire  _T_686 = _T_475 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_687 = _T_678 | _T_686; // @[el2_ifu_compress_ctl.scala 85:27]
  wire  _T_703 = _T_2 & _T_487; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_704 = _T_703 & _T_7; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_705 = _T_704 & _T_9; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_706 = _T_705 & _T_50; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_707 = _T_706 & _T_52; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_708 = _T_707 & _T_54; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_709 = _T_708 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_710 = _T_687 | _T_709; // @[el2_ifu_compress_ctl.scala 86:27]
  wire  _T_717 = _T_56 & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_718 = _T_717 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_719 = _T_710 | _T_718; // @[el2_ifu_compress_ctl.scala 87:41]
  wire  _T_726 = _T_56 & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_727 = _T_726 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_728 = _T_719 | _T_727; // @[el2_ifu_compress_ctl.scala 88:27]
  wire  _T_735 = _T_56 & io_din[4]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_736 = _T_735 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_737 = _T_728 | _T_736; // @[el2_ifu_compress_ctl.scala 89:27]
  wire  _T_744 = _T_56 & io_din[3]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_745 = _T_744 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_746 = _T_737 | _T_745; // @[el2_ifu_compress_ctl.scala 90:27]
  wire  _T_753 = _T_56 & io_din[2]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_754 = _T_753 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_755 = _T_746 | _T_754; // @[el2_ifu_compress_ctl.scala 91:27]
  wire  _T_764 = _T_194 & _T_4; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_765 = _T_764 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_766 = _T_755 | _T_765; // @[el2_ifu_compress_ctl.scala 92:27]
  wire  rdrs1 = _T_766 | _T_195; // @[el2_ifu_compress_ctl.scala 93:30]
  wire  _T_777 = io_din[15] & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_778 = _T_777 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_782 = io_din[15] & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_783 = _T_782 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_784 = _T_778 | _T_783; // @[el2_ifu_compress_ctl.scala 96:34]
  wire  _T_788 = io_din[15] & io_din[4]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_789 = _T_788 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_790 = _T_784 | _T_789; // @[el2_ifu_compress_ctl.scala 96:54]
  wire  _T_794 = io_din[15] & io_din[3]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_795 = _T_794 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_796 = _T_790 | _T_795; // @[el2_ifu_compress_ctl.scala 96:74]
  wire  _T_800 = io_din[15] & io_din[2]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_801 = _T_800 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_802 = _T_796 | _T_801; // @[el2_ifu_compress_ctl.scala 96:94]
  wire  _T_807 = _T_200 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  rs2rs2 = _T_802 | _T_807; // @[el2_ifu_compress_ctl.scala 96:114]
  wire  rdprd = _T_12 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_820 = io_din[15] & _T_4; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_821 = _T_820 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_827 = _T_821 | _T_234; // @[el2_ifu_compress_ctl.scala 100:36]
  wire  _T_830 = ~io_din[1]; // @[el2_ifu_compress_ctl.scala 29:83]
  wire  _T_831 = io_din[14] & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_834 = _T_831 & _T_147; // @[el2_ifu_compress_ctl.scala 100:76]
  wire  rdprs1 = _T_827 | _T_834; // @[el2_ifu_compress_ctl.scala 100:57]
  wire  _T_846 = _T_128 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_847 = _T_846 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_851 = io_din[15] & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_854 = _T_851 & _T_147; // @[el2_ifu_compress_ctl.scala 102:66]
  wire  rs2prs2 = _T_847 | _T_854; // @[el2_ifu_compress_ctl.scala 102:47]
  wire  _T_859 = _T_190 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  rs2prd = _T_859 & _T_147; // @[el2_ifu_compress_ctl.scala 103:33]
  wire  _T_866 = _T_2 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  uimm9_2 = _T_866 & _T_147; // @[el2_ifu_compress_ctl.scala 104:34]
  wire  _T_875 = _T_317 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  ulwimm6_2 = _T_875 & _T_147; // @[el2_ifu_compress_ctl.scala 105:39]
  wire  ulwspimm7_2 = _T_317 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_897 = _T_317 & io_din[13]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_898 = _T_897 & _T_23; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_899 = _T_898 & _T_38; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_900 = _T_899 & _T_40; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_901 = _T_900 & io_din[8]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  rdeq2 = _T_901 & _T_44; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1027 = _T_194 & io_din[13]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  rdeq1 = _T_482 | _T_1027; // @[el2_ifu_compress_ctl.scala 110:42]
  wire  _T_1050 = io_din[14] & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1051 = rdeq2 | _T_1050; // @[el2_ifu_compress_ctl.scala 111:53]
  wire  rs1eq2 = _T_1051 | uimm9_2; // @[el2_ifu_compress_ctl.scala 111:71]
  wire  _T_1092 = _T_357 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1093 = _T_1092 & _T_38; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1094 = _T_1093 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  simm5_0 = _T_1094 | _T_643; // @[el2_ifu_compress_ctl.scala 114:45]
  wire  _T_1112 = _T_897 & io_din[7]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1121 = _T_897 & _T_42; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1122 = _T_1112 | _T_1121; // @[el2_ifu_compress_ctl.scala 116:44]
  wire  _T_1130 = _T_897 & io_din[9]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1131 = _T_1122 | _T_1130; // @[el2_ifu_compress_ctl.scala 117:29]
  wire  _T_1139 = _T_897 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1140 = _T_1131 | _T_1139; // @[el2_ifu_compress_ctl.scala 118:28]
  wire  _T_1148 = _T_897 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  sluimm17_12 = _T_1140 | _T_1148; // @[el2_ifu_compress_ctl.scala 119:29]
  wire  uimm5_0 = _T_79 | _T_195; // @[el2_ifu_compress_ctl.scala 121:45]
  wire [6:0] l1_6 = {out_6,out_5,out_4,_T_228,out_2,1'h1,1'h1}; // @[Cat.scala 29:58]
  wire [4:0] _T_1192 = rdrd ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1193 = rdprd ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1194 = rs2prd ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1195 = rdeq1 ? 5'h1 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1196 = rdeq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1197 = _T_1192 | _T_1193; // @[Mux.scala 27:72]
  wire [4:0] _T_1198 = _T_1197 | _T_1194; // @[Mux.scala 27:72]
  wire [4:0] _T_1199 = _T_1198 | _T_1195; // @[Mux.scala 27:72]
  wire [4:0] l1_11 = _T_1199 | _T_1196; // @[Mux.scala 27:72]
  wire [4:0] _T_1210 = rdrs1 ? rdd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1211 = rdprs1 ? rdpd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1212 = rs1eq2 ? 5'h2 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1213 = _T_1210 | _T_1211; // @[Mux.scala 27:72]
  wire [4:0] l1_19 = _T_1213 | _T_1212; // @[Mux.scala 27:72]
  wire [4:0] _T_1219 = {3'h0,1'h0,out_20}; // @[Cat.scala 29:58]
  wire [4:0] _T_1222 = rs2rs2 ? rs2d : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1223 = rs2prs2 ? rs2pd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1224 = _T_1222 | _T_1223; // @[Mux.scala 27:72]
  wire [4:0] l1_24 = _T_1219 | _T_1224; // @[el2_ifu_compress_ctl.scala 134:67]
  wire [14:0] _T_1232 = {out_14,out_13,out_12,l1_11,l1_6}; // @[Cat.scala 29:58]
  wire [16:0] _T_1234 = {1'h0,out_30,2'h0,3'h0,l1_24,l1_19}; // @[Cat.scala 29:58]
  wire [31:0] l1 = {1'h0,out_30,2'h0,3'h0,l1_24,l1_19,_T_1232}; // @[Cat.scala 29:58]
  wire [5:0] simm5d = {io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [1:0] _T_1241 = {io_din[5],io_din[6]}; // @[Cat.scala 29:58]
  wire [5:0] _T_1242 = {io_din[10:7],io_din[12:11]}; // @[Cat.scala 29:58]
  wire [1:0] _T_1248 = {io_din[2],io_din[6]}; // @[Cat.scala 29:58]
  wire [3:0] _T_1250 = {io_din[12],io_din[4:3],io_din[5]}; // @[Cat.scala 29:58]
  wire [5:0] simm9d = {io_din[12],io_din[4:3],io_din[5],io_din[2],io_din[6]}; // @[Cat.scala 29:58]
  wire [3:0] _T_1254 = {io_din[5],io_din[12:10]}; // @[Cat.scala 29:58]
  wire [2:0] _T_1258 = {io_din[3:2],io_din[12]}; // @[Cat.scala 29:58]
  wire [10:0] sjald_1 = {io_din[12],io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:4],io_din[3]}; // @[Cat.scala 29:58]
  wire [8:0] sjald_12 = io_din[12] ? 9'h1ff : 9'h0; // @[Bitwise.scala 72:12]
  wire [19:0] sjald = {sjald_12,io_din[12],io_din[8],io_din[10:9],io_din[6],io_din[7],io_din[2],io_din[11],io_din[5:4],io_din[3]}; // @[Cat.scala 29:58]
  wire [14:0] _T_1281 = io_din[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [19:0] sluimmd = {_T_1281,rs2d}; // @[Cat.scala 29:58]
  wire [6:0] _T_1287 = simm5d[5] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_1289 = {_T_1287,simm5d[4:0]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1292 = {2'h0,io_din[10:7],io_din[12:11],io_din[5],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [2:0] _T_1296 = simm9d[5] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_1299 = {_T_1296,simm9d[4:0],4'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1302 = {5'h0,io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1305 = {4'h0,io_din[3:2],io_din[12],io_din[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1307 = {6'h0,io_din[12],rs2d}; // @[Cat.scala 29:58]
  wire [11:0] _T_1312 = {sjald[19],sjald[9:0],sjald[10]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1314 = simm5_0 ? _T_1289 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1315 = uimm9_2 ? _T_1292 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1316 = rdeq2 ? _T_1299 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1317 = ulwimm6_2 ? _T_1302 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1318 = ulwspimm7_2 ? _T_1305 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1319 = uimm5_0 ? _T_1307 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1320 = _T_228 ? _T_1312 : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1321 = sluimm17_12 ? sluimmd[19:8] : 12'h0; // @[Mux.scala 27:72]
  wire [11:0] _T_1322 = _T_1314 | _T_1315; // @[Mux.scala 27:72]
  wire [11:0] _T_1323 = _T_1322 | _T_1316; // @[Mux.scala 27:72]
  wire [11:0] _T_1324 = _T_1323 | _T_1317; // @[Mux.scala 27:72]
  wire [11:0] _T_1325 = _T_1324 | _T_1318; // @[Mux.scala 27:72]
  wire [11:0] _T_1326 = _T_1325 | _T_1319; // @[Mux.scala 27:72]
  wire [11:0] _T_1327 = _T_1326 | _T_1320; // @[Mux.scala 27:72]
  wire [11:0] _T_1328 = _T_1327 | _T_1321; // @[Mux.scala 27:72]
  wire [8:0] _T_1336 = _T_228 ? sjald[19:11] : 9'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_1337 = sluimm17_12 ? sluimmd[7:0] : 8'h0; // @[Mux.scala 27:72]
  wire [8:0] _GEN_0 = {{1'd0}, _T_1337}; // @[Mux.scala 27:72]
  wire [8:0] _T_1338 = _T_1336 | _GEN_0; // @[Mux.scala 27:72]
  wire [8:0] _GEN_1 = {{1'd0}, l1[19:12]}; // @[el2_ifu_compress_ctl.scala 162:25]
  wire [8:0] l2_19 = _GEN_1 | _T_1338; // @[el2_ifu_compress_ctl.scala 162:25]
  wire [32:0] l2 = {io_l2_31,l2_19,l1[11:0]}; // @[Cat.scala 29:58]
  wire [8:0] sbr8d = {io_din[12],io_din[6],io_din[5],io_din[2],io_din[11],io_din[10],io_din[4],io_din[3],1'h0}; // @[Cat.scala 29:58]
  wire [6:0] uswimm6d = {io_din[5],io_din[12:10],io_din[6],2'h0}; // @[Cat.scala 29:58]
  wire [7:0] uswspimm7d = {io_din[8:7],io_din[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [3:0] _T_1369 = sbr8d[8] ? 4'hf : 4'h0; // @[Bitwise.scala 72:12]
  wire [6:0] _T_1371 = {_T_1369,sbr8d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1374 = {5'h0,uswimm6d[6:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1377 = {4'h0,uswspimm7d[7:5]}; // @[Cat.scala 29:58]
  wire [6:0] _T_1378 = _T_234 ? _T_1371 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1379 = _T_854 ? _T_1374 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1380 = _T_807 ? _T_1377 : 7'h0; // @[Mux.scala 27:72]
  wire [6:0] _T_1381 = _T_1378 | _T_1379; // @[Mux.scala 27:72]
  wire [6:0] _T_1382 = _T_1381 | _T_1380; // @[Mux.scala 27:72]
  wire [6:0] l3_31 = l2[31:25] | _T_1382; // @[el2_ifu_compress_ctl.scala 170:25]
  wire [12:0] l3_24 = l2[24:12]; // @[el2_ifu_compress_ctl.scala 173:17]
  wire [4:0] _T_1388 = {sbr8d[4:1],sbr8d[8]}; // @[Cat.scala 29:58]
  wire [4:0] _T_1393 = _T_234 ? _T_1388 : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1394 = _T_854 ? uswimm6d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1395 = _T_807 ? uswspimm7d[4:0] : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_1396 = _T_1393 | _T_1394; // @[Mux.scala 27:72]
  wire [4:0] _T_1397 = _T_1396 | _T_1395; // @[Mux.scala 27:72]
  wire [4:0] l3_11 = l2[11:7] | _T_1397; // @[el2_ifu_compress_ctl.scala 174:24]
  wire [11:0] _T_1400 = {l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire [19:0] _T_1401 = {l3_31,l3_24}; // @[Cat.scala 29:58]
  wire [31:0] l3 = {l3_31,l3_24,l3_11,l2[6:0]}; // @[Cat.scala 29:58]
  wire  _T_1408 = _T_4 & _T_487; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1409 = _T_1408 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1410 = _T_1409 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1413 = _T_1410 & _T_147; // @[el2_ifu_compress_ctl.scala 179:39]
  wire  _T_1421 = _T_1408 & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1422 = _T_1421 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1425 = _T_1422 & _T_147; // @[el2_ifu_compress_ctl.scala 179:79]
  wire  _T_1426 = _T_1413 | _T_1425; // @[el2_ifu_compress_ctl.scala 179:54]
  wire  _T_1435 = _T_642 & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1436 = _T_1435 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1437 = _T_1426 | _T_1436; // @[el2_ifu_compress_ctl.scala 179:94]
  wire  _T_1445 = _T_1408 & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1446 = _T_1445 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1449 = _T_1446 & _T_147; // @[el2_ifu_compress_ctl.scala 180:55]
  wire  _T_1450 = _T_1437 | _T_1449; // @[el2_ifu_compress_ctl.scala 180:30]
  wire  _T_1458 = _T_1408 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1459 = _T_1458 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1462 = _T_1459 & _T_147; // @[el2_ifu_compress_ctl.scala 180:96]
  wire  _T_1463 = _T_1450 | _T_1462; // @[el2_ifu_compress_ctl.scala 180:70]
  wire  _T_1472 = _T_642 & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1473 = _T_1472 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1474 = _T_1463 | _T_1473; // @[el2_ifu_compress_ctl.scala 180:111]
  wire  _T_1481 = io_din[15] & _T_487; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1482 = _T_1481 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1483 = _T_1482 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1484 = _T_1474 | _T_1483; // @[el2_ifu_compress_ctl.scala 181:29]
  wire  _T_1492 = _T_1408 & io_din[9]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1493 = _T_1492 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1496 = _T_1493 & _T_147; // @[el2_ifu_compress_ctl.scala 181:79]
  wire  _T_1497 = _T_1484 | _T_1496; // @[el2_ifu_compress_ctl.scala 181:54]
  wire  _T_1504 = _T_487 & io_din[6]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1505 = _T_1504 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1506 = _T_1505 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1507 = _T_1497 | _T_1506; // @[el2_ifu_compress_ctl.scala 181:94]
  wire  _T_1516 = _T_642 & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1517 = _T_1516 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1518 = _T_1507 | _T_1517; // @[el2_ifu_compress_ctl.scala 181:118]
  wire  _T_1526 = _T_1408 & io_din[8]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1527 = _T_1526 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1530 = _T_1527 & _T_147; // @[el2_ifu_compress_ctl.scala 182:28]
  wire  _T_1531 = _T_1518 | _T_1530; // @[el2_ifu_compress_ctl.scala 181:144]
  wire  _T_1538 = _T_487 & io_din[5]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1539 = _T_1538 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1540 = _T_1539 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1541 = _T_1531 | _T_1540; // @[el2_ifu_compress_ctl.scala 182:43]
  wire  _T_1550 = _T_642 & io_din[10]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1551 = _T_1550 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1552 = _T_1541 | _T_1551; // @[el2_ifu_compress_ctl.scala 182:67]
  wire  _T_1560 = _T_1408 & io_din[7]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1561 = _T_1560 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1564 = _T_1561 & _T_147; // @[el2_ifu_compress_ctl.scala 183:28]
  wire  _T_1565 = _T_1552 | _T_1564; // @[el2_ifu_compress_ctl.scala 182:94]
  wire  _T_1573 = io_din[12] & io_din[11]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1574 = _T_1573 & _T_38; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1575 = _T_1574 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1576 = _T_1575 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1577 = _T_1565 | _T_1576; // @[el2_ifu_compress_ctl.scala 183:43]
  wire  _T_1586 = _T_642 & io_din[9]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1587 = _T_1586 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1588 = _T_1577 | _T_1587; // @[el2_ifu_compress_ctl.scala 183:71]
  wire  _T_1596 = _T_1408 & io_din[4]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1597 = _T_1596 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1600 = _T_1597 & _T_147; // @[el2_ifu_compress_ctl.scala 184:28]
  wire  _T_1601 = _T_1588 | _T_1600; // @[el2_ifu_compress_ctl.scala 183:97]
  wire  _T_1607 = io_din[13] & io_din[12]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1608 = _T_1607 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1609 = _T_1608 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1610 = _T_1601 | _T_1609; // @[el2_ifu_compress_ctl.scala 184:43]
  wire  _T_1619 = _T_642 & io_din[8]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1620 = _T_1619 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1621 = _T_1610 | _T_1620; // @[el2_ifu_compress_ctl.scala 184:67]
  wire  _T_1629 = _T_1408 & io_din[3]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1630 = _T_1629 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1633 = _T_1630 & _T_147; // @[el2_ifu_compress_ctl.scala 185:28]
  wire  _T_1634 = _T_1621 | _T_1633; // @[el2_ifu_compress_ctl.scala 184:93]
  wire  _T_1640 = io_din[13] & io_din[4]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1641 = _T_1640 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1642 = _T_1641 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1643 = _T_1634 | _T_1642; // @[el2_ifu_compress_ctl.scala 185:43]
  wire  _T_1651 = _T_1408 & io_din[2]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1652 = _T_1651 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1655 = _T_1652 & _T_147; // @[el2_ifu_compress_ctl.scala 185:91]
  wire  _T_1656 = _T_1643 | _T_1655; // @[el2_ifu_compress_ctl.scala 185:66]
  wire  _T_1665 = _T_642 & io_din[7]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1666 = _T_1665 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1667 = _T_1656 | _T_1666; // @[el2_ifu_compress_ctl.scala 185:106]
  wire  _T_1673 = io_din[13] & io_din[3]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1674 = _T_1673 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1675 = _T_1674 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1676 = _T_1667 | _T_1675; // @[el2_ifu_compress_ctl.scala 186:29]
  wire  _T_1682 = io_din[13] & io_din[2]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1683 = _T_1682 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1684 = _T_1683 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1685 = _T_1676 | _T_1684; // @[el2_ifu_compress_ctl.scala 186:52]
  wire  _T_1691 = io_din[14] & _T_4; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1692 = _T_1691 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1693 = _T_1685 | _T_1692; // @[el2_ifu_compress_ctl.scala 186:75]
  wire  _T_1702 = _T_703 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1703 = _T_1702 & io_din[0]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1704 = _T_1693 | _T_1703; // @[el2_ifu_compress_ctl.scala 186:98]
  wire  _T_1711 = _T_820 & io_din[12]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1712 = _T_1711 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1715 = _T_1712 & _T_147; // @[el2_ifu_compress_ctl.scala 187:54]
  wire  _T_1716 = _T_1704 | _T_1715; // @[el2_ifu_compress_ctl.scala 187:29]
  wire  _T_1725 = _T_642 & _T_487; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1726 = _T_1725 & io_din[1]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1729 = _T_1726 & _T_147; // @[el2_ifu_compress_ctl.scala 187:96]
  wire  _T_1730 = _T_1716 | _T_1729; // @[el2_ifu_compress_ctl.scala 187:69]
  wire  _T_1739 = _T_642 & io_din[12]; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1740 = _T_1739 & _T_830; // @[el2_ifu_compress_ctl.scala 29:110]
  wire  _T_1741 = _T_1730 | _T_1740; // @[el2_ifu_compress_ctl.scala 187:111]
  wire  _T_1748 = _T_1691 & _T_147; // @[el2_ifu_compress_ctl.scala 188:50]
  wire  legal = _T_1741 | _T_1748; // @[el2_ifu_compress_ctl.scala 188:30]
  wire [31:0] _T_1750 = legal ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [9:0] _T_1760 = {1'h0,out_30,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0,1'h0}; // @[Cat.scala 29:58]
  wire [18:0] _T_1769 = {_T_1760,1'h0,out_20,1'h0,1'h0,1'h0,1'h0,1'h0,out_14,out_13}; // @[Cat.scala 29:58]
  wire [27:0] _T_1778 = {_T_1769,out_12,1'h0,1'h0,1'h0,1'h0,1'h0,out_6,out_5,out_4}; // @[Cat.scala 29:58]
  wire [30:0] _T_1781 = {_T_1778,_T_228,out_2,1'h1}; // @[Cat.scala 29:58]
  assign io_dout = l3 & _T_1750; // @[el2_ifu_compress_ctl.scala 190:10]
  assign io_l1 = {_T_1234,_T_1232}; // @[el2_ifu_compress_ctl.scala 191:9]
  assign io_l2 = l2[31:0]; // @[el2_ifu_compress_ctl.scala 192:9]
  assign io_l3 = {_T_1401,_T_1400}; // @[el2_ifu_compress_ctl.scala 193:9]
  assign io_legal = _T_1741 | _T_1748; // @[el2_ifu_compress_ctl.scala 194:12]
  assign io_o = {_T_1781,1'h1}; // @[el2_ifu_compress_ctl.scala 195:8]
  assign io_sluimmd = {_T_1281,rs2d}; // @[el2_ifu_compress_ctl.scala 150:14]
  assign io_uimm5d = {io_din[12],rs2d}; // @[el2_ifu_compress_ctl.scala 205:13]
  assign io_ulwspimm7d = {_T_1258,io_din[6:4]}; // @[el2_ifu_compress_ctl.scala 206:17]
  assign io_ulwimm6d = {_T_1254,io_din[6]}; // @[el2_ifu_compress_ctl.scala 207:15]
  assign io_simm9d = {_T_1250,_T_1248}; // @[el2_ifu_compress_ctl.scala 208:13]
  assign io_uimm9d = {_T_1242,_T_1241}; // @[el2_ifu_compress_ctl.scala 209:13]
  assign io_simm5d = {io_din[12],rs2d}; // @[el2_ifu_compress_ctl.scala 210:13]
  assign io_sjald = {sjald_12,sjald_1}; // @[el2_ifu_compress_ctl.scala 204:12]
  assign io_l2_31 = l1[31:20] | _T_1328; // @[el2_ifu_compress_ctl.scala 152:12]
endmodule
