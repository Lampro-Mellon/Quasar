module rvecc_encode_64(
  input  [63:0] io_din,
  output [6:0]  io_ecc_out
);
  wire  w0_0 = io_din[0]; // @[el2_lib.scala 343:39]
  wire  w0_1 = io_din[1]; // @[el2_lib.scala 343:39]
  wire  w1_1 = io_din[2]; // @[el2_lib.scala 344:39]
  wire  w0_2 = io_din[3]; // @[el2_lib.scala 343:39]
  wire  w0_3 = io_din[4]; // @[el2_lib.scala 343:39]
  wire  w1_3 = io_din[5]; // @[el2_lib.scala 344:39]
  wire  w0_4 = io_din[6]; // @[el2_lib.scala 343:39]
  wire  w2_3 = io_din[7]; // @[el2_lib.scala 345:39]
  wire  w0_5 = io_din[8]; // @[el2_lib.scala 343:39]
  wire  w1_5 = io_din[9]; // @[el2_lib.scala 344:39]
  wire  w0_6 = io_din[10]; // @[el2_lib.scala 343:39]
  wire  w0_7 = io_din[11]; // @[el2_lib.scala 343:39]
  wire  w1_7 = io_din[12]; // @[el2_lib.scala 344:39]
  wire  w0_8 = io_din[13]; // @[el2_lib.scala 343:39]
  wire  w2_7 = io_din[14]; // @[el2_lib.scala 345:39]
  wire  w0_9 = io_din[15]; // @[el2_lib.scala 343:39]
  wire  w1_9 = io_din[16]; // @[el2_lib.scala 344:39]
  wire  w0_10 = io_din[17]; // @[el2_lib.scala 343:39]
  wire  w3_7 = io_din[18]; // @[el2_lib.scala 346:39]
  wire  w0_11 = io_din[19]; // @[el2_lib.scala 343:39]
  wire  w1_11 = io_din[20]; // @[el2_lib.scala 344:39]
  wire  w0_12 = io_din[21]; // @[el2_lib.scala 343:39]
  wire  w2_11 = io_din[22]; // @[el2_lib.scala 345:39]
  wire  w0_13 = io_din[23]; // @[el2_lib.scala 343:39]
  wire  w1_13 = io_din[24]; // @[el2_lib.scala 344:39]
  wire  w0_14 = io_din[25]; // @[el2_lib.scala 343:39]
  wire  w0_15 = io_din[26]; // @[el2_lib.scala 343:39]
  wire  w1_15 = io_din[27]; // @[el2_lib.scala 344:39]
  wire  w0_16 = io_din[28]; // @[el2_lib.scala 343:39]
  wire  w2_15 = io_din[29]; // @[el2_lib.scala 345:39]
  wire  w0_17 = io_din[30]; // @[el2_lib.scala 343:39]
  wire  w1_17 = io_din[31]; // @[el2_lib.scala 344:39]
  wire  w0_18 = io_din[32]; // @[el2_lib.scala 343:39]
  wire  w3_15 = io_din[33]; // @[el2_lib.scala 346:39]
  wire  w0_19 = io_din[34]; // @[el2_lib.scala 343:39]
  wire  w1_19 = io_din[35]; // @[el2_lib.scala 344:39]
  wire  w0_20 = io_din[36]; // @[el2_lib.scala 343:39]
  wire  w2_19 = io_din[37]; // @[el2_lib.scala 345:39]
  wire  w0_21 = io_din[38]; // @[el2_lib.scala 343:39]
  wire  w1_21 = io_din[39]; // @[el2_lib.scala 344:39]
  wire  w0_22 = io_din[40]; // @[el2_lib.scala 343:39]
  wire  w4_15 = io_din[41]; // @[el2_lib.scala 347:39]
  wire  w0_23 = io_din[42]; // @[el2_lib.scala 343:39]
  wire  w1_23 = io_din[43]; // @[el2_lib.scala 344:39]
  wire  w0_24 = io_din[44]; // @[el2_lib.scala 343:39]
  wire  w2_23 = io_din[45]; // @[el2_lib.scala 345:39]
  wire  w0_25 = io_din[46]; // @[el2_lib.scala 343:39]
  wire  w1_25 = io_din[47]; // @[el2_lib.scala 344:39]
  wire  w0_26 = io_din[48]; // @[el2_lib.scala 343:39]
  wire  w3_23 = io_din[49]; // @[el2_lib.scala 346:39]
  wire  w0_27 = io_din[50]; // @[el2_lib.scala 343:39]
  wire  w1_27 = io_din[51]; // @[el2_lib.scala 344:39]
  wire  w0_28 = io_din[52]; // @[el2_lib.scala 343:39]
  wire  w2_27 = io_din[53]; // @[el2_lib.scala 345:39]
  wire  w0_29 = io_din[54]; // @[el2_lib.scala 343:39]
  wire  w1_29 = io_din[55]; // @[el2_lib.scala 344:39]
  wire  w0_30 = io_din[56]; // @[el2_lib.scala 343:39]
  wire  w0_31 = io_din[57]; // @[el2_lib.scala 343:39]
  wire  w1_31 = io_din[58]; // @[el2_lib.scala 344:39]
  wire  w0_32 = io_din[59]; // @[el2_lib.scala 343:39]
  wire  w2_31 = io_din[60]; // @[el2_lib.scala 345:39]
  wire  w0_33 = io_din[61]; // @[el2_lib.scala 343:39]
  wire  w1_33 = io_din[62]; // @[el2_lib.scala 344:39]
  wire  w0_34 = io_din[63]; // @[el2_lib.scala 343:39]
  wire [6:0] _T_210 = {w0_34,w1_33,w0_33,w2_31,w0_32,w1_31,w0_31}; // @[el2_lib.scala 351:27]
  wire  _T_211 = ^_T_210; // @[el2_lib.scala 351:34]
  wire [6:0] _T_217 = {w0_18,w1_17,w0_17,w2_15,w0_16,w1_15,w0_15}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_224 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15}; // @[el2_lib.scala 351:44]
  wire [14:0] _T_225 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15,_T_217}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_232 = {w0_26,w1_25,w0_25,w2_23,w0_24,w1_23,w0_23,w4_15}; // @[el2_lib.scala 351:44]
  wire [30:0] _T_241 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_225}; // @[el2_lib.scala 351:44]
  wire  _T_242 = ^_T_241; // @[el2_lib.scala 351:51]
  wire [6:0] _T_248 = {w0_10,w1_9,w0_9,w2_7,w0_8,w1_7,w0_7}; // @[el2_lib.scala 351:61]
  wire [14:0] _T_256 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_248}; // @[el2_lib.scala 351:61]
  wire [30:0] _T_272 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_256}; // @[el2_lib.scala 351:61]
  wire  _T_273 = ^_T_272; // @[el2_lib.scala 351:68]
  wire [6:0] _T_279 = {w0_6,w1_5,w0_5,w2_3,w0_4,w1_3,w0_3}; // @[el2_lib.scala 351:78]
  wire [14:0] _T_287 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_279}; // @[el2_lib.scala 351:78]
  wire [30:0] _T_303 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_224,_T_287}; // @[el2_lib.scala 351:78]
  wire  _T_304 = ^_T_303; // @[el2_lib.scala 351:85]
  wire [7:0] _T_311 = {w2_7,w0_6,w1_5,w0_5,w2_3,w0_2,w1_1,w0_1}; // @[el2_lib.scala 351:95]
  wire [16:0] _T_320 = {w0_17,w2_15,w0_14,w1_13,w0_13,w2_11,w0_10,w1_9,w0_9,_T_311}; // @[el2_lib.scala 351:95]
  wire [8:0] _T_328 = {w1_25,w0_25,w2_23,w0_22,w1_21,w0_21,w2_19,w0_18,w1_17}; // @[el2_lib.scala 351:95]
  wire [17:0] _T_337 = {w0_34,w1_33,w0_33,w2_31,w0_30,w1_29,w0_29,w2_27,w0_26,_T_328}; // @[el2_lib.scala 351:95]
  wire [34:0] _T_338 = {_T_337,_T_320}; // @[el2_lib.scala 351:95]
  wire  _T_339 = ^_T_338; // @[el2_lib.scala 351:102]
  wire [7:0] _T_346 = {w1_7,w0_6,w1_5,w0_4,w1_3,w0_2,w1_1,w0_0}; // @[el2_lib.scala 351:112]
  wire [16:0] _T_355 = {w0_16,w1_15,w0_14,w1_13,w0_12,w1_11,w0_10,w1_9,w0_8,_T_346}; // @[el2_lib.scala 351:112]
  wire [8:0] _T_363 = {w1_25,w0_24,w1_23,w0_22,w1_21,w0_20,w1_19,w0_18,w1_17}; // @[el2_lib.scala 351:112]
  wire [17:0] _T_372 = {w0_34,w1_33,w0_32,w1_31,w0_30,w1_29,w0_28,w1_27,w0_26,_T_363}; // @[el2_lib.scala 351:112]
  wire [34:0] _T_373 = {_T_372,_T_355}; // @[el2_lib.scala 351:112]
  wire  _T_374 = ^_T_373; // @[el2_lib.scala 351:119]
  wire [7:0] _T_381 = {w0_7,w0_6,w0_5,w0_4,w0_3,w0_2,w0_1,w0_0}; // @[el2_lib.scala 351:129]
  wire [16:0] _T_390 = {w0_16,w0_15,w0_14,w0_13,w0_12,w0_11,w0_10,w0_9,w0_8,_T_381}; // @[el2_lib.scala 351:129]
  wire [8:0] _T_398 = {w0_25,w0_24,w0_23,w0_22,w0_21,w0_20,w0_19,w0_18,w0_17}; // @[el2_lib.scala 351:129]
  wire [17:0] _T_407 = {w0_34,w0_33,w0_32,w0_31,w0_30,w0_29,w0_28,w0_27,w0_26,_T_398}; // @[el2_lib.scala 351:129]
  wire [34:0] _T_408 = {_T_407,_T_390}; // @[el2_lib.scala 351:129]
  wire  _T_409 = ^_T_408; // @[el2_lib.scala 351:136]
  wire [2:0] _T_411 = {_T_339,_T_374,_T_409}; // @[Cat.scala 29:58]
  wire [3:0] _T_414 = {_T_211,_T_242,_T_273,_T_304}; // @[Cat.scala 29:58]
  assign io_ecc_out = {_T_414,_T_411}; // @[el2_lib.scala 351:16]
endmodule
module el2_ifu_mem_ctl(
  input          clock,
  input          reset,
  input          io_free_clk,
  input          io_active_clk,
  input          io_exu_flush_final,
  input          io_dec_tlu_flush_lower_wb,
  input          io_dec_tlu_flush_err_wb,
  input          io_dec_tlu_i0_commit_cmt,
  input          io_dec_tlu_force_halt,
  input  [30:0]  io_ifc_fetch_addr_bf,
  input          io_ifc_fetch_uncacheable_bf,
  input          io_ifc_fetch_req_bf,
  input          io_ifc_fetch_req_bf_raw,
  input          io_ifc_iccm_access_bf,
  input          io_ifc_region_acc_fault_bf,
  input          io_ifc_dma_access_ok,
  input          io_dec_tlu_fence_i_wb,
  input          io_ifu_bp_hit_taken_f,
  input          io_ifu_bp_inst_mask_f,
  input          io_ifu_axi_arready,
  input          io_ifu_axi_rvalid,
  input  [2:0]   io_ifu_axi_rid,
  input  [63:0]  io_ifu_axi_rdata,
  input  [1:0]   io_ifu_axi_rresp,
  input          io_ifu_bus_clk_en,
  input          io_dma_iccm_req,
  input  [31:0]  io_dma_mem_addr,
  input  [2:0]   io_dma_mem_sz,
  input          io_dma_mem_write,
  input  [63:0]  io_dma_mem_wdata,
  input  [2:0]   io_dma_mem_tag,
  input  [63:0]  io_ic_rd_data,
  input  [70:0]  io_ic_debug_rd_data,
  input  [25:0]  io_ictag_debug_rd_data,
  input  [1:0]   io_ic_eccerr,
  input  [1:0]   io_ic_parerr,
  input  [1:0]   io_ic_rd_hit,
  input          io_ic_tag_perr,
  input  [63:0]  io_iccm_rd_data,
  input  [77:0]  io_iccm_rd_data_ecc,
  input  [1:0]   io_ifu_fetch_val,
  input  [70:0]  io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0]  io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input          io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input          io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output         io_ifu_miss_state_idle,
  output         io_ifu_ic_mb_empty,
  output         io_ic_dma_active,
  output         io_ic_write_stall,
  output         io_ifu_pmu_ic_miss,
  output         io_ifu_pmu_ic_hit,
  output         io_ifu_pmu_bus_error,
  output         io_ifu_pmu_bus_busy,
  output         io_ifu_pmu_bus_trxn,
  output         io_ifu_axi_awvalid,
  output [2:0]   io_ifu_axi_awid,
  output [31:0]  io_ifu_axi_awaddr,
  output [3:0]   io_ifu_axi_awregion,
  output [7:0]   io_ifu_axi_awlen,
  output [2:0]   io_ifu_axi_awsize,
  output [1:0]   io_ifu_axi_awburst,
  output         io_ifu_axi_awlock,
  output [3:0]   io_ifu_axi_awcache,
  output [2:0]   io_ifu_axi_awprot,
  output [3:0]   io_ifu_axi_awqos,
  output         io_ifu_axi_wvalid,
  output [63:0]  io_ifu_axi_wdata,
  output [7:0]   io_ifu_axi_wstrb,
  output         io_ifu_axi_wlast,
  output         io_ifu_axi_bready,
  output         io_ifu_axi_arvalid,
  output [2:0]   io_ifu_axi_arid,
  output [31:0]  io_ifu_axi_araddr,
  output [3:0]   io_ifu_axi_arregion,
  output [7:0]   io_ifu_axi_arlen,
  output [2:0]   io_ifu_axi_arsize,
  output [1:0]   io_ifu_axi_arburst,
  output         io_ifu_axi_arlock,
  output [3:0]   io_ifu_axi_arcache,
  output [2:0]   io_ifu_axi_arprot,
  output [3:0]   io_ifu_axi_arqos,
  output         io_ifu_axi_rready,
  output         io_iccm_dma_ecc_error,
  output         io_iccm_dma_rvalid,
  output [63:0]  io_iccm_dma_rdata,
  output [2:0]   io_iccm_dma_rtag,
  output         io_iccm_ready,
  output [30:0]  io_ic_rw_addr,
  output [1:0]   io_ic_wr_en,
  output         io_ic_rd_en,
  output [70:0]  io_ic_wr_data_0,
  output [70:0]  io_ic_wr_data_1,
  output [70:0]  io_ic_debug_wr_data,
  output [70:0]  io_ifu_ic_debug_rd_data,
  output [9:0]   io_ic_debug_addr,
  output         io_ic_debug_rd_en,
  output         io_ic_debug_wr_en,
  output         io_ic_debug_tag_array,
  output [1:0]   io_ic_debug_way,
  output [1:0]   io_ic_tag_valid,
  output [14:0]  io_iccm_rw_addr,
  output         io_iccm_wren,
  output         io_iccm_rden,
  output [77:0]  io_iccm_wr_data,
  output [2:0]   io_iccm_wr_size,
  output         io_ic_hit_f,
  output         io_ic_access_fault_f,
  output [1:0]   io_ic_access_fault_type_f,
  output         io_iccm_rd_ecc_single_err,
  output         io_iccm_rd_ecc_double_err,
  output         io_ic_error_start,
  output         io_ifu_async_error_start,
  output         io_iccm_dma_sb_error,
  output [1:0]   io_ic_fetch_val_f,
  output [31:0]  io_ic_data_f,
  output [63:0]  io_ic_premux_data,
  output         io_ic_sel_premux_data,
  input          io_dec_tlu_core_ecc_disable,
  output         io_ifu_ic_debug_rd_data_valid,
  output         io_iccm_buf_correct_ecc,
  output         io_iccm_correction_state,
  input          io_scan_mode,
  output [141:0] io_data,
  output [6:0]   io_ic_wr_ecc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] m1_io_din; // @[el2_ifu_mem_ctl.scala 343:18]
  wire [6:0] m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 343:18]
  wire [63:0] m2_io_din; // @[el2_ifu_mem_ctl.scala 344:18]
  wire [6:0] m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 344:18]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 185:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 321:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 322:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 322:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 254:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 556:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 558:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 187:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 309:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 673:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 673:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 676:91]
  wire [1:0] _T_2240 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 676:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 323:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 276:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 676:113]
  wire [1:0] _T_2241 = _T_2240 & _GEN_465; // @[el2_ifu_mem_ctl.scala 676:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 662:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 676:130]
  wire [1:0] _T_2242 = _T_2241 | _GEN_466; // @[el2_ifu_mem_ctl.scala 676:130]
  wire  _T_2243 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 676:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_2243}; // @[el2_ifu_mem_ctl.scala 676:152]
  wire [1:0] _T_2244 = _T_2242 & _GEN_467; // @[el2_ifu_mem_ctl.scala 676:152]
  wire [1:0] _T_2233 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 676:91]
  wire [1:0] _T_2234 = _T_2233 & _GEN_465; // @[el2_ifu_mem_ctl.scala 676:113]
  wire [1:0] _T_2235 = _T_2234 | _GEN_466; // @[el2_ifu_mem_ctl.scala 676:130]
  wire [1:0] _T_2237 = _T_2235 & _GEN_467; // @[el2_ifu_mem_ctl.scala 676:152]
  wire [3:0] iccm_ecc_word_enable = {_T_2244,_T_2237}; // @[Cat.scala 29:58]
  wire  _T_2344 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_2345 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_2346 = _T_2344 ^ _T_2345; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2354 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_2355 = ^_T_2354; // @[el2_lib.scala 301:83]
  wire  _T_2356 = io_iccm_rd_data_ecc[37] ^ _T_2355; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2363 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2371 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2363}; // @[el2_lib.scala 301:103]
  wire  _T_2372 = ^_T_2371; // @[el2_lib.scala 301:110]
  wire  _T_2373 = io_iccm_rd_data_ecc[36] ^ _T_2372; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2380 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2388 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2380}; // @[el2_lib.scala 301:130]
  wire  _T_2389 = ^_T_2388; // @[el2_lib.scala 301:137]
  wire  _T_2390 = io_iccm_rd_data_ecc[35] ^ _T_2389; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2399 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2408 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2399}; // @[el2_lib.scala 301:157]
  wire  _T_2409 = ^_T_2408; // @[el2_lib.scala 301:164]
  wire  _T_2410 = io_iccm_rd_data_ecc[34] ^ _T_2409; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2419 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2428 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2419}; // @[el2_lib.scala 301:184]
  wire  _T_2429 = ^_T_2428; // @[el2_lib.scala 301:191]
  wire  _T_2430 = io_iccm_rd_data_ecc[33] ^ _T_2429; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2439 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2448 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_2439}; // @[el2_lib.scala 301:211]
  wire  _T_2449 = ^_T_2448; // @[el2_lib.scala 301:218]
  wire  _T_2450 = io_iccm_rd_data_ecc[32] ^ _T_2449; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2456 = {_T_2346,_T_2356,_T_2373,_T_2390,_T_2410,_T_2430,_T_2450}; // @[Cat.scala 29:58]
  wire  _T_2457 = _T_2456 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2458 = iccm_ecc_word_enable[0] & _T_2457; // @[el2_lib.scala 302:32]
  wire  _T_2460 = _T_2458 & _T_2456[6]; // @[el2_lib.scala 302:53]
  wire  _T_2729 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_2730 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_2731 = _T_2729 ^ _T_2730; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2739 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_2740 = ^_T_2739; // @[el2_lib.scala 301:83]
  wire  _T_2741 = io_iccm_rd_data_ecc[76] ^ _T_2740; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2748 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2756 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2748}; // @[el2_lib.scala 301:103]
  wire  _T_2757 = ^_T_2756; // @[el2_lib.scala 301:110]
  wire  _T_2758 = io_iccm_rd_data_ecc[75] ^ _T_2757; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2765 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2773 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2765}; // @[el2_lib.scala 301:130]
  wire  _T_2774 = ^_T_2773; // @[el2_lib.scala 301:137]
  wire  _T_2775 = io_iccm_rd_data_ecc[74] ^ _T_2774; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2784 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2793 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2784}; // @[el2_lib.scala 301:157]
  wire  _T_2794 = ^_T_2793; // @[el2_lib.scala 301:164]
  wire  _T_2795 = io_iccm_rd_data_ecc[73] ^ _T_2794; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2804 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2813 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2804}; // @[el2_lib.scala 301:184]
  wire  _T_2814 = ^_T_2813; // @[el2_lib.scala 301:191]
  wire  _T_2815 = io_iccm_rd_data_ecc[72] ^ _T_2814; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2824 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2833 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_2824}; // @[el2_lib.scala 301:211]
  wire  _T_2834 = ^_T_2833; // @[el2_lib.scala 301:218]
  wire  _T_2835 = io_iccm_rd_data_ecc[71] ^ _T_2834; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2841 = {_T_2731,_T_2741,_T_2758,_T_2775,_T_2795,_T_2815,_T_2835}; // @[Cat.scala 29:58]
  wire  _T_2842 = _T_2841 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2843 = iccm_ecc_word_enable[1] & _T_2842; // @[el2_lib.scala 302:32]
  wire  _T_2845 = _T_2843 & _T_2841[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_2460,_T_2845}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 190:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 640:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 192:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 485:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 192:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 192:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 192:72]
  wire  _T_1609 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1614 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1634 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 535:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 401:42]
  wire  _T_1636 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 535:79]
  wire  _T_1637 = _T_1634 | _T_1636; // @[el2_ifu_mem_ctl.scala 535:56]
  wire  _T_1638 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 535:122]
  wire  _T_1639 = ~_T_1638; // @[el2_ifu_mem_ctl.scala 535:101]
  wire  _T_1640 = _T_1637 & _T_1639; // @[el2_ifu_mem_ctl.scala 535:99]
  wire  _T_1641 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1655 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 542:45]
  wire  _T_1656 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 542:69]
  wire  _T_1657 = _T_1655 & _T_1656; // @[el2_ifu_mem_ctl.scala 542:67]
  wire  _T_1658 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_1641 ? _T_1657 : _T_1658; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_1614 ? _T_1640 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_1609 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 192:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 194:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 194:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 284:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 284:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 708:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 275:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 325:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 275:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 275:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 284:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 284:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 284:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 284:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 555:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 597:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 624:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 311:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 605:56]
  wire  _T_1760 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 622:69]
  wire  _T_1761 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 622:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_1760 : _T_1761; // @[el2_ifu_mem_ctl.scala 622:28]
  wire  _T_1707 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 601:68]
  wire  _T_1708 = ic_act_miss_f | _T_1707; // @[el2_ifu_mem_ctl.scala 601:48]
  wire  bus_reset_data_beat_cnt = _T_1708 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 601:91]
  wire  _T_1704 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 600:50]
  wire  _T_1705 = bus_ifu_wr_en_ff & _T_1704; // @[el2_ifu_mem_ctl.scala 600:48]
  wire  _T_1706 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 600:72]
  wire  bus_inc_data_beat_cnt = _T_1705 & _T_1706; // @[el2_ifu_mem_ctl.scala 600:70]
  wire [2:0] _T_1712 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 604:115]
  wire [2:0] _T_1714 = bus_inc_data_beat_cnt ? _T_1712 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_1709 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 602:32]
  wire  _T_1710 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 602:57]
  wire  bus_hold_data_beat_cnt = _T_1709 & _T_1710; // @[el2_ifu_mem_ctl.scala 602:55]
  wire [2:0] _T_1715 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_1714 | _T_1715; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 194:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 195:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 194:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 195:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 201:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 437:45]
  wire  _T_1279 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 458:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 414:60]
  wire  _T_1310 = _T_1279 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1283 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1311 = _T_1283 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1318 = _T_1310 | _T_1311; // @[Mux.scala 27:72]
  wire  _T_1287 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1312 = _T_1287 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1319 = _T_1318 | _T_1312; // @[Mux.scala 27:72]
  wire  _T_1291 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1313 = _T_1291 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1320 = _T_1319 | _T_1313; // @[Mux.scala 27:72]
  wire  _T_1295 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1314 = _T_1295 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1321 = _T_1320 | _T_1314; // @[Mux.scala 27:72]
  wire  _T_1299 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1315 = _T_1299 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1322 = _T_1321 | _T_1315; // @[Mux.scala 27:72]
  wire  _T_1303 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1316 = _T_1303 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1323 = _T_1322 | _T_1316; // @[Mux.scala 27:72]
  wire  _T_1307 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 458:127]
  wire  _T_1317 = _T_1307 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_1323 | _T_1317; // @[Mux.scala 27:72]
  wire  _T_1365 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 460:69]
  wire  _T_1366 = ic_miss_buff_data_valid_bypass_index & _T_1365; // @[el2_ifu_mem_ctl.scala 460:67]
  wire  _T_1368 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 460:91]
  wire  _T_1369 = _T_1366 & _T_1368; // @[el2_ifu_mem_ctl.scala 460:89]
  wire  _T_1374 = _T_1366 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 461:65]
  wire  _T_1375 = _T_1369 | _T_1374; // @[el2_ifu_mem_ctl.scala 460:112]
  wire  _T_1377 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 462:43]
  wire  _T_1380 = _T_1377 & _T_1368; // @[el2_ifu_mem_ctl.scala 462:65]
  wire  _T_1381 = _T_1375 | _T_1380; // @[el2_ifu_mem_ctl.scala 461:88]
  wire  _T_1385 = _T_1377 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 463:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 440:75]
  wire  _T_1325 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1349 = _T_1325 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1328 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1350 = _T_1328 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1357 = _T_1349 | _T_1350; // @[Mux.scala 27:72]
  wire  _T_1331 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1351 = _T_1331 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1358 = _T_1357 | _T_1351; // @[Mux.scala 27:72]
  wire  _T_1334 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1352 = _T_1334 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1359 = _T_1358 | _T_1352; // @[Mux.scala 27:72]
  wire  _T_1337 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1353 = _T_1337 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1360 = _T_1359 | _T_1353; // @[Mux.scala 27:72]
  wire  _T_1340 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1354 = _T_1340 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1361 = _T_1360 | _T_1354; // @[Mux.scala 27:72]
  wire  _T_1343 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1355 = _T_1343 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1362 = _T_1361 | _T_1355; // @[Mux.scala 27:72]
  wire  _T_1346 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 459:110]
  wire  _T_1356 = _T_1346 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_1362 | _T_1356; // @[Mux.scala 27:72]
  wire  _T_1386 = _T_1385 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 463:87]
  wire  _T_1387 = _T_1381 | _T_1386; // @[el2_ifu_mem_ctl.scala 462:88]
  wire  _T_1391 = ic_miss_buff_data_valid_bypass_index & _T_1307; // @[el2_ifu_mem_ctl.scala 464:43]
  wire  miss_buff_hit_unq_f = _T_1387 | _T_1391; // @[el2_ifu_mem_ctl.scala 463:131]
  wire  _T_1407 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 469:55]
  wire  _T_1408 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 469:87]
  wire  _T_1409 = _T_1407 | _T_1408; // @[el2_ifu_mem_ctl.scala 469:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_1409; // @[el2_ifu_mem_ctl.scala 469:41]
  wire  _T_1392 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 466:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 312:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 457:51]
  wire  _T_1393 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 466:68]
  wire  _T_1394 = miss_buff_hit_unq_f & _T_1393; // @[el2_ifu_mem_ctl.scala 466:66]
  wire  stream_hit_f = _T_1392 & _T_1394; // @[el2_ifu_mem_ctl.scala 466:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 279:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 279:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 279:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 607:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 634:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 205:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 205:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 205:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 205:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 207:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 208:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 209:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 209:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 209:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 197:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 209:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 209:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 210:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 210:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 210:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 210:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 211:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 212:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 209:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 208:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 207:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 206:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_1404 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 468:60]
  wire  _T_1405 = _T_1404 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 468:92]
  wire  stream_eol_f = _T_1405 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 468:110]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 220:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 220:87]
  wire  _T_113 = _T_111 & _T_1706; // @[el2_ifu_mem_ctl.scala 220:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 220:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 224:48]
  wire  _T_126 = _T_124 & _T_1706; // @[el2_ifu_mem_ctl.scala 224:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 285:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 285:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 285:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 285:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 285:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 285:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 286:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 339:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 286:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 286:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 286:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:50]
  wire  _T_137 = _T_135 & _T_1706; // @[el2_ifu_mem_ctl.scala 228:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 287:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 288:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 288:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 287:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:35]
  wire  _T_143 = _T_141 & _T_1706; // @[el2_ifu_mem_ctl.scala 229:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 234:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 233:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 238:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 238:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 195:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 195:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 195:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 195:91]
  wire  _T_30 = ic_act_miss_f & _T_1706; // @[el2_ifu_mem_ctl.scala 202:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 213:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 213:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 213:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 213:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 217:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 217:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 221:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 225:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 230:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 235:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 235:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 255:95]
  wire  _T_175 = _T_1407 & _T_174; // @[el2_ifu_mem_ctl.scala 255:93]
  wire  crit_wd_byp_ok_ff = _T_1408 | _T_175; // @[el2_ifu_mem_ctl.scala 255:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 256:36]
  wire  _T_180 = _T_1407 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 256:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 256:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 256:70]
  wire  _T_184 = _T_1407 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 257:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 257:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 256:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 257:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 258:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 258:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 257:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 260:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:35]
  reg [6:0] _T_4285; // @[el2_ifu_mem_ctl.scala 736:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_4285[5:0]; // @[el2_ifu_mem_ctl.scala 735:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 732:121]
  wire  _T_4150 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4152 = _T_4150 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3641; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_3641[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4153 = _T_4152 & _GEN_473; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4146 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4148 = _T_4146 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3637; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_3637[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4149 = _T_4148 & _GEN_475; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4142 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4144 = _T_4142 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3633; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_3633[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4145 = _T_4144 & _GEN_477; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4138 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4140 = _T_4138 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3629; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_3629[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4141 = _T_4140 & _GEN_479; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4134 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4136 = _T_4134 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3625; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_3625[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4137 = _T_4136 & _GEN_481; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4130 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4132 = _T_4130 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3621; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_3621[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4133 = _T_4132 & _GEN_483; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4126 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4128 = _T_4126 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3617; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_3617[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4129 = _T_4128 & _GEN_485; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4122 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4124 = _T_4122 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3613; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_3613[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4125 = _T_4124 & _GEN_487; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4118 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4120 = _T_4118 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3609; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_3609[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4121 = _T_4120 & _GEN_489; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4114 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4116 = _T_4114 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3605; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_3605[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4117 = _T_4116 & _GEN_491; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [59:0] _T_4162 = {_T_4153,_T_4149,_T_4145,_T_4141,_T_4137,_T_4133,_T_4129,_T_4125,_T_4121,_T_4117}; // @[Cat.scala 29:58]
  wire  _T_4110 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4112 = _T_4110 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3601; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_3601[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4113 = _T_4112 & _GEN_493; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4106 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4108 = _T_4106 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3597; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_3597[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4109 = _T_4108 & _GEN_495; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4102 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4104 = _T_4102 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3593; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_3593[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4105 = _T_4104 & _GEN_497; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4098 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4100 = _T_4098 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3589; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_3589[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4101 = _T_4100 & _GEN_499; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4094 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4096 = _T_4094 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3585; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_3585[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4097 = _T_4096 & _GEN_501; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4090 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4092 = _T_4090 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3581; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_3581[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4093 = _T_4092 & _GEN_503; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4086 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4088 = _T_4086 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3577; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_3577[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4089 = _T_4088 & _GEN_505; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4082 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4084 = _T_4082 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3573; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_3573[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4085 = _T_4084 & _GEN_507; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4078 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4080 = _T_4078 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3569; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_3569[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4081 = _T_4080 & _GEN_509; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [113:0] _T_4171 = {_T_4162,_T_4113,_T_4109,_T_4105,_T_4101,_T_4097,_T_4093,_T_4089,_T_4085,_T_4081}; // @[Cat.scala 29:58]
  wire  _T_4074 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4076 = _T_4074 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3565; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_3565[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4077 = _T_4076 & _GEN_511; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4070 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4072 = _T_4070 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3561; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_3561[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4073 = _T_4072 & _GEN_513; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4066 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4068 = _T_4066 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3557; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_3557[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4069 = _T_4068 & _GEN_515; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4062 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4064 = _T_4062 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3553; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_3553[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4065 = _T_4064 & _GEN_517; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4058 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4060 = _T_4058 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3549; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_3549[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4061 = _T_4060 & _GEN_519; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4054 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4056 = _T_4054 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3545; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_3545[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4057 = _T_4056 & _GEN_521; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4050 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4052 = _T_4050 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3541; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_3541[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4053 = _T_4052 & _GEN_523; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4046 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4048 = _T_4046 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3537; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_3537[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4049 = _T_4048 & _GEN_525; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4042 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4044 = _T_4042 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3533; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_3533[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4045 = _T_4044 & _GEN_527; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [167:0] _T_4180 = {_T_4171,_T_4077,_T_4073,_T_4069,_T_4065,_T_4061,_T_4057,_T_4053,_T_4049,_T_4045}; // @[Cat.scala 29:58]
  wire  _T_4038 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4040 = _T_4038 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3529; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_3529[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4041 = _T_4040 & _GEN_529; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4034 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4036 = _T_4034 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3525; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_3525[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4037 = _T_4036 & _GEN_531; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4030 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4032 = _T_4030 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3521; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_3521[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4033 = _T_4032 & _GEN_533; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4026 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4028 = _T_4026 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3517; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_3517[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4029 = _T_4028 & _GEN_535; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4022 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4024 = _T_4022 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3513; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_3513[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4025 = _T_4024 & _GEN_537; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4018 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4020 = _T_4018 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3509; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_3509[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4021 = _T_4020 & _GEN_539; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4014 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4016 = _T_4014 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3505; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_3505[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4017 = _T_4016 & _GEN_541; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4010 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4012 = _T_4010 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3501; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_3501[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4013 = _T_4012 & _GEN_543; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_4006 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4008 = _T_4006 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3497; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_3497[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4009 = _T_4008 & _GEN_545; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [221:0] _T_4189 = {_T_4180,_T_4041,_T_4037,_T_4033,_T_4029,_T_4025,_T_4021,_T_4017,_T_4013,_T_4009}; // @[Cat.scala 29:58]
  wire  _T_4002 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4004 = _T_4002 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3493; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_3493[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4005 = _T_4004 & _GEN_547; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3998 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_4000 = _T_3998 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3489; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_3489[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_4001 = _T_4000 & _GEN_549; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3994 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3996 = _T_3994 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3485; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_3485[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3997 = _T_3996 & _GEN_551; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3990 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3992 = _T_3990 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3481; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_3481[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3993 = _T_3992 & _GEN_553; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3986 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3988 = _T_3986 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3477; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_3477[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3989 = _T_3988 & _GEN_555; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3982 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3984 = _T_3982 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3473; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_3473[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3985 = _T_3984 & _GEN_557; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3978 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3980 = _T_3978 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3469; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_3469[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3981 = _T_3980 & _GEN_559; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3974 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3976 = _T_3974 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3465; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_3465[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3977 = _T_3976 & _GEN_561; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3970 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3972 = _T_3970 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3461; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_3461[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3973 = _T_3972 & _GEN_563; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [275:0] _T_4198 = {_T_4189,_T_4005,_T_4001,_T_3997,_T_3993,_T_3989,_T_3985,_T_3981,_T_3977,_T_3973}; // @[Cat.scala 29:58]
  wire  _T_3966 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3968 = _T_3966 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3457; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_3457[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3969 = _T_3968 & _GEN_565; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3962 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3964 = _T_3962 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3453; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_3453[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3965 = _T_3964 & _GEN_567; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3958 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3960 = _T_3958 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3449; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_3449[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3961 = _T_3960 & _GEN_569; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3954 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3956 = _T_3954 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3445; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_3445[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3957 = _T_3956 & _GEN_571; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3950 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3952 = _T_3950 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3441; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_3441[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3953 = _T_3952 & _GEN_573; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3946 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3948 = _T_3946 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3437; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_3437[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3949 = _T_3948 & _GEN_575; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3942 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3944 = _T_3942 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3433; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_3433[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3945 = _T_3944 & _GEN_577; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3938 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3940 = _T_3938 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3429; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_3429[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3941 = _T_3940 & _GEN_579; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3934 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3936 = _T_3934 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3425; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_3425[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3937 = _T_3936 & _GEN_581; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [329:0] _T_4207 = {_T_4198,_T_3969,_T_3965,_T_3961,_T_3957,_T_3953,_T_3949,_T_3945,_T_3941,_T_3937}; // @[Cat.scala 29:58]
  wire  _T_3930 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3932 = _T_3930 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3421; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_3421[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3933 = _T_3932 & _GEN_583; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3926 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3928 = _T_3926 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3417; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_3417[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3929 = _T_3928 & _GEN_585; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3922 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3924 = _T_3922 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3413; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_3413[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3925 = _T_3924 & _GEN_587; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3918 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3920 = _T_3918 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3409; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_3409[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3921 = _T_3920 & _GEN_589; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3914 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3916 = _T_3914 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3405; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_3405[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3917 = _T_3916 & _GEN_591; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3910 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3912 = _T_3910 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3401; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_3401[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3913 = _T_3912 & _GEN_593; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3906 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3908 = _T_3906 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3397; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_3397[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3909 = _T_3908 & _GEN_595; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3902 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3904 = _T_3902 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3393; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_3393[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3905 = _T_3904 & _GEN_597; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3898 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3900 = _T_3898 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3389; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_3389[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3901 = _T_3900 & _GEN_599; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [383:0] _T_4216 = {_T_4207,_T_3933,_T_3929,_T_3925,_T_3921,_T_3917,_T_3913,_T_3909,_T_3905,_T_3901}; // @[Cat.scala 29:58]
  wire  _T_3894 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3896 = _T_3894 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3385; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_3385[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3897 = _T_3896 & _GEN_600; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3890 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3892 = _T_3890 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3381; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_3381[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3893 = _T_3892 & _GEN_601; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3886 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3888 = _T_3886 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3377; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_3377[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3889 = _T_3888 & _GEN_602; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3882 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3884 = _T_3882 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3373; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_3373[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3885 = _T_3884 & _GEN_603; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3878 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3880 = _T_3878 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3369; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_3369[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3881 = _T_3880 & _GEN_604; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3874 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3876 = _T_3874 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3365; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_3365[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3877 = _T_3876 & _GEN_605; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3870 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3872 = _T_3870 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3361; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_3361[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3873 = _T_3872 & _GEN_606; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3866 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3868 = _T_3866 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3357; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_3357[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3869 = _T_3868 & _GEN_607; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3862 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3864 = _T_3862 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3353; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_3353[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3865 = _T_3864 & _GEN_608; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [437:0] _T_4225 = {_T_4216,_T_3897,_T_3893,_T_3889,_T_3885,_T_3881,_T_3877,_T_3873,_T_3869,_T_3865}; // @[Cat.scala 29:58]
  wire  _T_3858 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3860 = _T_3858 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3349; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_3349[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3861 = _T_3860 & _GEN_609; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3854 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3856 = _T_3854 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3345; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_3345[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3857 = _T_3856 & _GEN_610; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3850 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3852 = _T_3850 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3341; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_3341[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3853 = _T_3852 & _GEN_611; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3846 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3848 = _T_3846 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3337; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_3337[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3849 = _T_3848 & _GEN_612; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3842 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3844 = _T_3842 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3333; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_3333[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3845 = _T_3844 & _GEN_613; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3838 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3840 = _T_3838 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3329; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_3329[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3841 = _T_3840 & _GEN_614; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3834 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3836 = _T_3834 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3325; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_3325[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3837 = _T_3836 & _GEN_615; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3830 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3832 = _T_3830 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3321; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_3321[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3833 = _T_3832 & _GEN_616; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3826 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3828 = _T_3826 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3317; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_3317[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3829 = _T_3828 & _GEN_617; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [491:0] _T_4234 = {_T_4225,_T_3861,_T_3857,_T_3853,_T_3849,_T_3845,_T_3841,_T_3837,_T_3833,_T_3829}; // @[Cat.scala 29:58]
  wire  _T_3822 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3824 = _T_3822 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3313; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_3313[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3825 = _T_3824 & _GEN_618; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3818 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3820 = _T_3818 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3309; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_3309[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3821 = _T_3820 & _GEN_619; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3814 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3816 = _T_3814 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3305; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_3305[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3817 = _T_3816 & _GEN_620; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3810 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3812 = _T_3810 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3301; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_3301[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3813 = _T_3812 & _GEN_621; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3806 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3808 = _T_3806 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3297; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_3297[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3809 = _T_3808 & _GEN_622; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3802 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3804 = _T_3802 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3293; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_3293[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3805 = _T_3804 & _GEN_623; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3798 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3800 = _T_3798 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3289; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_3289[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3801 = _T_3800 & _GEN_624; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3794 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3796 = _T_3794 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3285; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_3285[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3797 = _T_3796 & _GEN_625; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3790 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3792 = _T_3790 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3281; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_3281[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3793 = _T_3792 & _GEN_626; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [545:0] _T_4243 = {_T_4234,_T_3825,_T_3821,_T_3817,_T_3813,_T_3809,_T_3805,_T_3801,_T_3797,_T_3793}; // @[Cat.scala 29:58]
  wire  _T_3786 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3788 = _T_3786 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3277; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_3277[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3789 = _T_3788 & _GEN_627; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3782 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3784 = _T_3782 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3273; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_3273[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3785 = _T_3784 & _GEN_628; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3778 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3780 = _T_3778 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3269; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_3269[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3781 = _T_3780 & _GEN_629; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3774 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3776 = _T_3774 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3265; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_3265[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3777 = _T_3776 & _GEN_630; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3770 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3772 = _T_3770 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3261; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_3261[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3773 = _T_3772 & _GEN_631; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3766 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3768 = _T_3766 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3257; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_3257[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3769 = _T_3768 & _GEN_632; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3762 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3764 = _T_3762 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3253; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_3253[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3765 = _T_3764 & _GEN_633; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3758 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3760 = _T_3758 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3249; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_3249[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3761 = _T_3760 & _GEN_634; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3754 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3756 = _T_3754 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3245; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_3245[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3757 = _T_3756 & _GEN_635; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [599:0] _T_4252 = {_T_4243,_T_3789,_T_3785,_T_3781,_T_3777,_T_3773,_T_3769,_T_3765,_T_3761,_T_3757}; // @[Cat.scala 29:58]
  wire  _T_3750 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3752 = _T_3750 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3241; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_3241[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3753 = _T_3752 & _GEN_636; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3746 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3748 = _T_3746 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3237; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_3237[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3749 = _T_3748 & _GEN_637; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3742 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3744 = _T_3742 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3233; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_3233[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3745 = _T_3744 & _GEN_638; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3738 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3740 = _T_3738 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3229; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_3229[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3741 = _T_3740 & _GEN_639; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3734 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3736 = _T_3734 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3225; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_3225[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3737 = _T_3736 & _GEN_640; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3730 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3732 = _T_3730 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3221; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_3221[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3733 = _T_3732 & _GEN_641; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3726 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3728 = _T_3726 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3217; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_3217[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3729 = _T_3728 & _GEN_642; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3722 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3724 = _T_3722 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3213; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_3213[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3725 = _T_3724 & _GEN_643; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3718 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3720 = _T_3718 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3209; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_3209[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3721 = _T_3720 & _GEN_644; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [653:0] _T_4261 = {_T_4252,_T_3753,_T_3749,_T_3745,_T_3741,_T_3737,_T_3733,_T_3729,_T_3725,_T_3721}; // @[Cat.scala 29:58]
  wire  _T_3714 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3716 = _T_3714 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3205; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_3205[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3717 = _T_3716 & _GEN_645; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3710 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3712 = _T_3710 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3201; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_3201[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3713 = _T_3712 & _GEN_646; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3706 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3708 = _T_3706 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3197; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_3197[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3709 = _T_3708 & _GEN_647; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3702 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3704 = _T_3702 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3193; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_3193[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3705 = _T_3704 & _GEN_648; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3698 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3700 = _T_3698 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3189; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_3189[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3701 = _T_3700 & _GEN_649; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3694 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3696 = _T_3694 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3185; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_3185[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3697 = _T_3696 & _GEN_650; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3690 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3692 = _T_3690 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3181; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_3181[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3693 = _T_3692 & _GEN_651; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3686 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3688 = _T_3686 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3177; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_3177[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3689 = _T_3688 & _GEN_652; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3682 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3684 = _T_3682 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3173; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_3173[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3685 = _T_3684 & _GEN_653; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [707:0] _T_4270 = {_T_4261,_T_3717,_T_3713,_T_3709,_T_3705,_T_3701,_T_3697,_T_3693,_T_3689,_T_3685}; // @[Cat.scala 29:58]
  wire  _T_3678 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3680 = _T_3678 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3169; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3169[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3681 = _T_3680 & _GEN_654; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3674 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3676 = _T_3674 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3165; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3165[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3677 = _T_3676 & _GEN_655; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3670 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3672 = _T_3670 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3161; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3161[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3673 = _T_3672 & _GEN_656; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3666 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3668 = _T_3666 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3157; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3157[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3669 = _T_3668 & _GEN_657; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3662 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3664 = _T_3662 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3153; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3153[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3665 = _T_3664 & _GEN_658; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3658 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3660 = _T_3658 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3149; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3149[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3661 = _T_3660 & _GEN_659; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3654 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3656 = _T_3654 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3145; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3145[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3657 = _T_3656 & _GEN_660; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3650 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3652 = _T_3650 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3141; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3141[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3653 = _T_3652 & _GEN_661; // @[el2_ifu_mem_ctl.scala 732:130]
  wire  _T_3646 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3648 = _T_3646 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3137; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3137[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3649 = _T_3648 & _GEN_662; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [761:0] _T_4279 = {_T_4270,_T_3681,_T_3677,_T_3673,_T_3669,_T_3665,_T_3661,_T_3657,_T_3653,_T_3649}; // @[Cat.scala 29:58]
  wire  _T_3642 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 732:121]
  wire [5:0] _T_3644 = _T_3642 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3133; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3133[0]; // @[el2_ifu_mem_ctl.scala 729:30 el2_ifu_mem_ctl.scala 731:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [5:0] _T_3645 = _T_3644 & _GEN_663; // @[el2_ifu_mem_ctl.scala 732:130]
  wire [767:0] _T_4280 = {_T_4279,_T_3645}; // @[Cat.scala 29:58]
  wire  way_status = _T_4280[0]; // @[el2_ifu_mem_ctl.scala 732:16]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 263:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 265:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 272:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 277:59]
  wire  _T_214 = _T_212 | _T_1392; // @[el2_ifu_mem_ctl.scala 277:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 277:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 283:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 283:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 283:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 290:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 290:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 290:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 291:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 291:32]
  wire  _T_274 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 294:75]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 294:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_1781 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 630:48]
  wire  _T_1782 = _T_1781 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 630:52]
  wire  bus_ifu_wr_data_error_ff = _T_1782 & miss_pending; // @[el2_ifu_mem_ctl.scala 630:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 376:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 375:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 294:145]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 294:143]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 297:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 298:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 317:30]
  wire  _T_9230 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 785:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 318:24]
  wire  _T_9232 = _T_9230 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 785:51]
  wire  _T_9234 = _T_9232 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 785:67]
  wire  _T_9236 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 785:86]
  wire  replace_way_mb_any_0 = _T_9234 | _T_9236; // @[el2_ifu_mem_ctl.scala 785:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9239 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:50]
  wire  _T_9241 = _T_9239 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:66]
  wire  _T_9243 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:85]
  wire  _T_9245 = _T_9243 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:100]
  wire  replace_way_mb_any_1 = _T_9241 | _T_9245; // @[el2_ifu_mem_ctl.scala 786:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 302:110]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 306:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 306:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 307:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 306:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 308:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 316:23]
  wire  _T_313 = _T_1407 & flush_final_f; // @[el2_ifu_mem_ctl.scala 320:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 320:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 320:53]
  wire  _T_1399 = ~_T_1394; // @[el2_ifu_mem_ctl.scala 467:46]
  wire  _T_1400 = _T_1392 & _T_1399; // @[el2_ifu_mem_ctl.scala 467:44]
  wire  stream_miss_f = _T_1400 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 467:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 320:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 320:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 326:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_1392; // @[el2_ifu_mem_ctl.scala 328:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 328:82]
  wire  _T_1413 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 472:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_1413}; // @[Cat.scala 29:58]
  wire  _T_1414 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1438 = _T_1414 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1417 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1439 = _T_1417 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1438 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1420 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1440 = _T_1420 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1423 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1441 = _T_1423 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1426 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1442 = _T_1426 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1429 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1443 = _T_1429 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1450 = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1432 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1444 = _T_1432 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1451 = _T_1450 | _T_1444; // @[Mux.scala 27:72]
  wire  _T_1435 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 473:81]
  wire  _T_1445 = _T_1435 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_1451 | _T_1445; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 474:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 332:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 332:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 627:61]
  wire  _T_1775 = ic_act_miss_f_delayed & _T_1408; // @[el2_ifu_mem_ctl.scala 628:53]
  wire  reset_tag_valid_for_miss = _T_1775 & _T_17; // @[el2_ifu_mem_ctl.scala 628:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 332:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 334:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 336:84]
  wire  _T_1769 = ~_T_1781; // @[el2_ifu_mem_ctl.scala 625:84]
  wire  _T_1770 = _T_100 & _T_1769; // @[el2_ifu_mem_ctl.scala 625:82]
  wire  bus_ifu_wr_en_ff_q = _T_1770 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 625:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 336:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 337:31]
  wire [6:0] ic_wr_ecc = m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 346:13]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] ic_miss_buff_ecc = m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 350:20]
  wire [3:0] _T_1454 = {ifu_bus_rid_ff[2:1],_T_1413,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1455 = _T_1454 == 4'h0; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_1502 = _T_1455 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1458 = _T_1454 == 4'h1; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_1503 = _T_1458 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1518 = _T_1502 | _T_1503; // @[Mux.scala 27:72]
  wire  _T_1461 = _T_1454 == 4'h2; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_1504 = _T_1461 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1519 = _T_1518 | _T_1504; // @[Mux.scala 27:72]
  wire  _T_1464 = _T_1454 == 4'h3; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_1505 = _T_1464 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1520 = _T_1519 | _T_1505; // @[Mux.scala 27:72]
  wire  _T_1467 = _T_1454 == 4'h4; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_1506 = _T_1467 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1521 = _T_1520 | _T_1506; // @[Mux.scala 27:72]
  wire  _T_1470 = _T_1454 == 4'h5; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_1507 = _T_1470 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1522 = _T_1521 | _T_1507; // @[Mux.scala 27:72]
  wire  _T_1473 = _T_1454 == 4'h6; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_1508 = _T_1473 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1523 = _T_1522 | _T_1508; // @[Mux.scala 27:72]
  wire  _T_1476 = _T_1454 == 4'h7; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_1509 = _T_1476 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1524 = _T_1523 | _T_1509; // @[Mux.scala 27:72]
  wire  _T_1479 = _T_1454 == 4'h8; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_1510 = _T_1479 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1525 = _T_1524 | _T_1510; // @[Mux.scala 27:72]
  wire  _T_1482 = _T_1454 == 4'h9; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_1511 = _T_1482 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1526 = _T_1525 | _T_1511; // @[Mux.scala 27:72]
  wire  _T_1485 = _T_1454 == 4'ha; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_1512 = _T_1485 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1527 = _T_1526 | _T_1512; // @[Mux.scala 27:72]
  wire  _T_1488 = _T_1454 == 4'hb; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_1513 = _T_1488 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1528 = _T_1527 | _T_1513; // @[Mux.scala 27:72]
  wire  _T_1491 = _T_1454 == 4'hc; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_1514 = _T_1491 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1529 = _T_1528 | _T_1514; // @[Mux.scala 27:72]
  wire  _T_1494 = _T_1454 == 4'hd; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_1515 = _T_1494 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1530 = _T_1529 | _T_1515; // @[Mux.scala 27:72]
  wire  _T_1497 = _T_1454 == 4'he; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_1516 = _T_1497 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1531 = _T_1530 | _T_1516; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1454 == 4'hf; // @[el2_ifu_mem_ctl.scala 475:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_1517 = _T_1500 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1532 = _T_1531 | _T_1517; // @[Mux.scala 27:72]
  wire [3:0] _T_1534 = {ifu_bus_rid_ff[2:1],_T_1413,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1535 = _T_1534 == 4'h0; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1558 = _T_1535 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1538 = _T_1534 == 4'h1; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1559 = _T_1538 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1566 = _T_1558 | _T_1559; // @[Mux.scala 27:72]
  wire  _T_1541 = _T_1534 == 4'h2; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1560 = _T_1541 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1567 = _T_1566 | _T_1560; // @[Mux.scala 27:72]
  wire  _T_1544 = _T_1534 == 4'h3; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1561 = _T_1544 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1568 = _T_1567 | _T_1561; // @[Mux.scala 27:72]
  wire  _T_1547 = _T_1534 == 4'h4; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1562 = _T_1547 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1569 = _T_1568 | _T_1562; // @[Mux.scala 27:72]
  wire  _T_1550 = _T_1534 == 4'h5; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1563 = _T_1550 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1570 = _T_1569 | _T_1563; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1534 == 4'h6; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1564 = _T_1553 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1571 = _T_1570 | _T_1564; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1534 == 4'h7; // @[el2_ifu_mem_ctl.scala 476:64]
  wire [31:0] _T_1565 = _T_1556 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1572 = _T_1571 | _T_1565; // @[Mux.scala 27:72]
  wire [141:0] _T_393 = {ic_wr_ecc,ifu_bus_rdata_ff,ic_miss_buff_ecc,_T_1532,_T_1572}; // @[Cat.scala 29:58]
  wire [141:0] _T_396 = {ic_miss_buff_ecc,_T_1532,_T_1572,ic_wr_ecc,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_393 : _T_396; // @[el2_ifu_mem_ctl.scala 366:28]
  wire  _T_353 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 356:56]
  wire  _T_354 = _T_353 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 356:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 422:28]
  wire  _T_572 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 623:35]
  wire  _T_441 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_441; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_498 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 413:118]
  wire  _T_499 = ic_miss_buff_data_valid[0] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_499; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_595 = _T_572 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_575 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_442 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_442; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_502 = ic_miss_buff_data_valid[1] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_502; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_596 = _T_575 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_603 = _T_595 | _T_596; // @[Mux.scala 27:72]
  wire  _T_578 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_443 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_443; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_505 = ic_miss_buff_data_valid[2] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_505; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_597 = _T_578 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_604 = _T_603 | _T_597; // @[Mux.scala 27:72]
  wire  _T_581 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_444 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_444; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_508 = ic_miss_buff_data_valid[3] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_508; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_598 = _T_581 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_605 = _T_604 | _T_598; // @[Mux.scala 27:72]
  wire  _T_584 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_445 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_445; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_511 = ic_miss_buff_data_valid[4] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_511; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_599 = _T_584 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_606 = _T_605 | _T_599; // @[Mux.scala 27:72]
  wire  _T_587 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_446 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_446; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_514 = ic_miss_buff_data_valid[5] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_514; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_600 = _T_587 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_607 = _T_606 | _T_600; // @[Mux.scala 27:72]
  wire  _T_590 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_447 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_447; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_517 = ic_miss_buff_data_valid[6] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_517; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_601 = _T_590 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_608 = _T_607 | _T_601; // @[Mux.scala 27:72]
  wire  _T_593 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 424:114]
  wire  _T_448 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 407:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_448; // @[el2_ifu_mem_ctl.scala 407:73]
  wire  _T_520 = ic_miss_buff_data_valid[7] & _T_498; // @[el2_ifu_mem_ctl.scala 413:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_520; // @[el2_ifu_mem_ctl.scala 413:88]
  wire  _T_602 = _T_593 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_608 | _T_602; // @[Mux.scala 27:72]
  wire  _T_611 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 425:58]
  wire  _T_612 = bypass_valid_value_check & _T_611; // @[el2_ifu_mem_ctl.scala 425:56]
  wire  _T_614 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 425:77]
  wire  _T_615 = _T_612 & _T_614; // @[el2_ifu_mem_ctl.scala 425:75]
  wire  _T_620 = _T_612 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 426:75]
  wire  _T_621 = _T_615 | _T_620; // @[el2_ifu_mem_ctl.scala 425:95]
  wire  _T_623 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 427:56]
  wire  _T_626 = _T_623 & _T_614; // @[el2_ifu_mem_ctl.scala 427:74]
  wire  _T_627 = _T_621 | _T_626; // @[el2_ifu_mem_ctl.scala 426:94]
  wire  _T_631 = _T_623 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 428:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 423:70]
  wire  _T_632 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_648 = _T_632 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_634 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_649 = _T_634 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_656 = _T_648 | _T_649; // @[Mux.scala 27:72]
  wire  _T_636 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_650 = _T_636 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_657 = _T_656 | _T_650; // @[Mux.scala 27:72]
  wire  _T_638 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_651 = _T_638 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_658 = _T_657 | _T_651; // @[Mux.scala 27:72]
  wire  _T_640 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_652 = _T_640 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_659 = _T_658 | _T_652; // @[Mux.scala 27:72]
  wire  _T_642 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_653 = _T_642 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_660 = _T_659 | _T_653; // @[Mux.scala 27:72]
  wire  _T_644 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_654 = _T_644 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_661 = _T_660 | _T_654; // @[Mux.scala 27:72]
  wire  _T_646 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 428:132]
  wire  _T_655 = _T_646 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_662 = _T_661 | _T_655; // @[Mux.scala 27:72]
  wire  _T_664 = _T_631 & _T_662; // @[el2_ifu_mem_ctl.scala 428:69]
  wire  _T_665 = _T_627 | _T_664; // @[el2_ifu_mem_ctl.scala 427:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 429:95]
  wire  _T_668 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 429:95]
  wire  _T_669 = bypass_valid_value_check & _T_668; // @[el2_ifu_mem_ctl.scala 429:56]
  wire  bypass_data_ready_in = _T_665 | _T_669; // @[el2_ifu_mem_ctl.scala 428:181]
  wire  _T_670 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 433:53]
  wire  _T_671 = _T_670 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 433:73]
  wire  _T_673 = _T_671 & _T_317; // @[el2_ifu_mem_ctl.scala 433:96]
  wire  _T_675 = _T_673 & _T_58; // @[el2_ifu_mem_ctl.scala 433:118]
  wire  _T_677 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 434:73]
  wire  _T_679 = _T_677 & _T_317; // @[el2_ifu_mem_ctl.scala 434:96]
  wire  _T_681 = _T_679 & _T_58; // @[el2_ifu_mem_ctl.scala 434:118]
  wire  _T_682 = _T_675 | _T_681; // @[el2_ifu_mem_ctl.scala 433:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 436:58]
  wire  _T_683 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 435:54]
  wire  _T_684 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 435:76]
  wire  _T_685 = _T_683 & _T_684; // @[el2_ifu_mem_ctl.scala 435:74]
  wire  _T_687 = _T_685 & _T_317; // @[el2_ifu_mem_ctl.scala 435:96]
  wire  ic_crit_wd_rdy_new_in = _T_682 | _T_687; // @[el2_ifu_mem_ctl.scala 434:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 633:43]
  wire  _T_408 = ic_crit_wd_rdy | _T_1392; // @[el2_ifu_mem_ctl.scala 380:38]
  wire  _T_410 = _T_408 | _T_1408; // @[el2_ifu_mem_ctl.scala 380:64]
  wire  _T_411 = ~_T_410; // @[el2_ifu_mem_ctl.scala 380:21]
  wire  _T_412 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 380:98]
  wire  sel_ic_data = _T_411 & _T_412; // @[el2_ifu_mem_ctl.scala 380:96]
  wire  _T_1575 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 478:44]
  wire  _T_781 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 447:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 419:60]
  wire  _T_725 = _T_572 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_726 = _T_575 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_733 = _T_725 | _T_726; // @[Mux.scala 27:72]
  wire  _T_727 = _T_578 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_734 = _T_733 | _T_727; // @[Mux.scala 27:72]
  wire  _T_728 = _T_581 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_735 = _T_734 | _T_728; // @[Mux.scala 27:72]
  wire  _T_729 = _T_584 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_736 = _T_735 | _T_729; // @[Mux.scala 27:72]
  wire  _T_730 = _T_587 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_737 = _T_736 | _T_730; // @[Mux.scala 27:72]
  wire  _T_731 = _T_590 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_738 = _T_737 | _T_731; // @[Mux.scala 27:72]
  wire  _T_732 = _T_593 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_738 | _T_732; // @[Mux.scala 27:72]
  wire  _T_764 = _T_1325 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_765 = _T_1328 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_772 = _T_764 | _T_765; // @[Mux.scala 27:72]
  wire  _T_766 = _T_1331 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_773 = _T_772 | _T_766; // @[Mux.scala 27:72]
  wire  _T_767 = _T_1334 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_774 = _T_773 | _T_767; // @[Mux.scala 27:72]
  wire  _T_768 = _T_1337 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_775 = _T_774 | _T_768; // @[Mux.scala 27:72]
  wire  _T_769 = _T_1340 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_776 = _T_775 | _T_769; // @[Mux.scala 27:72]
  wire  _T_770 = _T_1343 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_777 = _T_776 | _T_770; // @[Mux.scala 27:72]
  wire  _T_771 = _T_1346 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_777 | _T_771; // @[Mux.scala 27:72]
  wire  _T_782 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 449:70]
  wire  ifu_byp_data_err_new = _T_781 ? ic_miss_buff_data_error_bypass : _T_782; // @[el2_ifu_mem_ctl.scala 447:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 391:42]
  wire  _T_1576 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 478:91]
  wire  _T_1577 = ~_T_1576; // @[el2_ifu_mem_ctl.scala 478:60]
  wire  ic_rd_parity_final_err = _T_1575 & _T_1577; // @[el2_ifu_mem_ctl.scala 478:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_8848 = _T_3642 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 760:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_8850 = _T_3646 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9103 = _T_8848 | _T_8850; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_8852 = _T_3650 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9104 = _T_9103 | _T_8852; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_8854 = _T_3654 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9105 = _T_9104 | _T_8854; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_8856 = _T_3658 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9106 = _T_9105 | _T_8856; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_8858 = _T_3662 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9107 = _T_9106 | _T_8858; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_8860 = _T_3666 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9108 = _T_9107 | _T_8860; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_8862 = _T_3670 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9109 = _T_9108 | _T_8862; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_8864 = _T_3674 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9110 = _T_9109 | _T_8864; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_8866 = _T_3678 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9111 = _T_9110 | _T_8866; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_8868 = _T_3682 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9112 = _T_9111 | _T_8868; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_8870 = _T_3686 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9113 = _T_9112 | _T_8870; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_8872 = _T_3690 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9114 = _T_9113 | _T_8872; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_8874 = _T_3694 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9115 = _T_9114 | _T_8874; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_8876 = _T_3698 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9116 = _T_9115 | _T_8876; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_8878 = _T_3702 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9117 = _T_9116 | _T_8878; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_8880 = _T_3706 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9118 = _T_9117 | _T_8880; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_8882 = _T_3710 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9119 = _T_9118 | _T_8882; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_8884 = _T_3714 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9120 = _T_9119 | _T_8884; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_8886 = _T_3718 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9121 = _T_9120 | _T_8886; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_8888 = _T_3722 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9122 = _T_9121 | _T_8888; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_8890 = _T_3726 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9123 = _T_9122 | _T_8890; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_8892 = _T_3730 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9124 = _T_9123 | _T_8892; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_8894 = _T_3734 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9125 = _T_9124 | _T_8894; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_8896 = _T_3738 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9126 = _T_9125 | _T_8896; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_8898 = _T_3742 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9127 = _T_9126 | _T_8898; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_8900 = _T_3746 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9128 = _T_9127 | _T_8900; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_8902 = _T_3750 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9129 = _T_9128 | _T_8902; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_8904 = _T_3754 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9130 = _T_9129 | _T_8904; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_8906 = _T_3758 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9131 = _T_9130 | _T_8906; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_8908 = _T_3762 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9132 = _T_9131 | _T_8908; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_8910 = _T_3766 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9133 = _T_9132 | _T_8910; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_8912 = _T_3770 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9134 = _T_9133 | _T_8912; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_8914 = _T_3774 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9135 = _T_9134 | _T_8914; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_8916 = _T_3778 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9136 = _T_9135 | _T_8916; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_8918 = _T_3782 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9137 = _T_9136 | _T_8918; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_8920 = _T_3786 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9138 = _T_9137 | _T_8920; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_8922 = _T_3790 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9139 = _T_9138 | _T_8922; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_8924 = _T_3794 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9140 = _T_9139 | _T_8924; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_8926 = _T_3798 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9141 = _T_9140 | _T_8926; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_8928 = _T_3802 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9142 = _T_9141 | _T_8928; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_8930 = _T_3806 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9143 = _T_9142 | _T_8930; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_8932 = _T_3810 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9144 = _T_9143 | _T_8932; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_8934 = _T_3814 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9145 = _T_9144 | _T_8934; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_8936 = _T_3818 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9146 = _T_9145 | _T_8936; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_8938 = _T_3822 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9147 = _T_9146 | _T_8938; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_8940 = _T_3826 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9148 = _T_9147 | _T_8940; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_8942 = _T_3830 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9149 = _T_9148 | _T_8942; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_8944 = _T_3834 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9150 = _T_9149 | _T_8944; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_8946 = _T_3838 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9151 = _T_9150 | _T_8946; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_8948 = _T_3842 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9152 = _T_9151 | _T_8948; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_8950 = _T_3846 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9153 = _T_9152 | _T_8950; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_8952 = _T_3850 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9154 = _T_9153 | _T_8952; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_8954 = _T_3854 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9155 = _T_9154 | _T_8954; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_8956 = _T_3858 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9156 = _T_9155 | _T_8956; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_8958 = _T_3862 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9157 = _T_9156 | _T_8958; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_8960 = _T_3866 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9158 = _T_9157 | _T_8960; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_8962 = _T_3870 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9159 = _T_9158 | _T_8962; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_8964 = _T_3874 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9160 = _T_9159 | _T_8964; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_8966 = _T_3878 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9161 = _T_9160 | _T_8966; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_8968 = _T_3882 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9162 = _T_9161 | _T_8968; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_8970 = _T_3886 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9163 = _T_9162 | _T_8970; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_8972 = _T_3890 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9164 = _T_9163 | _T_8972; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_8974 = _T_3894 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9165 = _T_9164 | _T_8974; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_8976 = _T_3898 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9166 = _T_9165 | _T_8976; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_8978 = _T_3902 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9167 = _T_9166 | _T_8978; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_8980 = _T_3906 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9168 = _T_9167 | _T_8980; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_8982 = _T_3910 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9169 = _T_9168 | _T_8982; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_8984 = _T_3914 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9170 = _T_9169 | _T_8984; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_8986 = _T_3918 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9171 = _T_9170 | _T_8986; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_8988 = _T_3922 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9172 = _T_9171 | _T_8988; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_8990 = _T_3926 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9173 = _T_9172 | _T_8990; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_8992 = _T_3930 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9174 = _T_9173 | _T_8992; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_8994 = _T_3934 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9175 = _T_9174 | _T_8994; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_8996 = _T_3938 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9176 = _T_9175 | _T_8996; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_8998 = _T_3942 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9177 = _T_9176 | _T_8998; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9000 = _T_3946 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9178 = _T_9177 | _T_9000; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9002 = _T_3950 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9179 = _T_9178 | _T_9002; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9004 = _T_3954 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9180 = _T_9179 | _T_9004; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9006 = _T_3958 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9181 = _T_9180 | _T_9006; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9008 = _T_3962 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9182 = _T_9181 | _T_9008; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9010 = _T_3966 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9183 = _T_9182 | _T_9010; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9012 = _T_3970 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9184 = _T_9183 | _T_9012; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9014 = _T_3974 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9185 = _T_9184 | _T_9014; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9016 = _T_3978 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9186 = _T_9185 | _T_9016; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9018 = _T_3982 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9187 = _T_9186 | _T_9018; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9020 = _T_3986 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9188 = _T_9187 | _T_9020; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9022 = _T_3990 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9189 = _T_9188 | _T_9022; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9024 = _T_3994 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9190 = _T_9189 | _T_9024; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9026 = _T_3998 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9191 = _T_9190 | _T_9026; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9028 = _T_4002 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9192 = _T_9191 | _T_9028; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9030 = _T_4006 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9193 = _T_9192 | _T_9030; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9032 = _T_4010 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9194 = _T_9193 | _T_9032; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9034 = _T_4014 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9195 = _T_9194 | _T_9034; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9036 = _T_4018 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9196 = _T_9195 | _T_9036; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9038 = _T_4022 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9197 = _T_9196 | _T_9038; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9040 = _T_4026 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9198 = _T_9197 | _T_9040; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9042 = _T_4030 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9199 = _T_9198 | _T_9042; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9044 = _T_4034 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9200 = _T_9199 | _T_9044; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9046 = _T_4038 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9201 = _T_9200 | _T_9046; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9048 = _T_4042 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9202 = _T_9201 | _T_9048; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9050 = _T_4046 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9203 = _T_9202 | _T_9050; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9052 = _T_4050 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9204 = _T_9203 | _T_9052; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9054 = _T_4054 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9205 = _T_9204 | _T_9054; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9056 = _T_4058 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9206 = _T_9205 | _T_9056; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9058 = _T_4062 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9207 = _T_9206 | _T_9058; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9060 = _T_4066 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9208 = _T_9207 | _T_9060; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9062 = _T_4070 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9209 = _T_9208 | _T_9062; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9064 = _T_4074 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9210 = _T_9209 | _T_9064; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9066 = _T_4078 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9211 = _T_9210 | _T_9066; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9068 = _T_4082 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9212 = _T_9211 | _T_9068; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9070 = _T_4086 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9213 = _T_9212 | _T_9070; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9072 = _T_4090 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9214 = _T_9213 | _T_9072; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9074 = _T_4094 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9215 = _T_9214 | _T_9074; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9076 = _T_4098 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9216 = _T_9215 | _T_9076; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9078 = _T_4102 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9217 = _T_9216 | _T_9078; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9080 = _T_4106 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9218 = _T_9217 | _T_9080; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9082 = _T_4110 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9219 = _T_9218 | _T_9082; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9084 = _T_4114 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9220 = _T_9219 | _T_9084; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9086 = _T_4118 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9221 = _T_9220 | _T_9086; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9088 = _T_4122 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9222 = _T_9221 | _T_9088; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9090 = _T_4126 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9223 = _T_9222 | _T_9090; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9092 = _T_4130 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9224 = _T_9223 | _T_9092; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9094 = _T_4134 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9225 = _T_9224 | _T_9094; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9096 = _T_4138 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9226 = _T_9225 | _T_9096; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9098 = _T_4142 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9227 = _T_9226 | _T_9098; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9100 = _T_4146 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9228 = _T_9227 | _T_9100; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9102 = _T_4150 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9229 = _T_9228 | _T_9102; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8465 = _T_3642 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 760:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8467 = _T_3646 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8720 = _T_8465 | _T_8467; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8469 = _T_3650 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8721 = _T_8720 | _T_8469; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8471 = _T_3654 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8722 = _T_8721 | _T_8471; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8473 = _T_3658 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8723 = _T_8722 | _T_8473; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8475 = _T_3662 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8724 = _T_8723 | _T_8475; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8477 = _T_3666 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8725 = _T_8724 | _T_8477; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8479 = _T_3670 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8726 = _T_8725 | _T_8479; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8481 = _T_3674 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8727 = _T_8726 | _T_8481; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8483 = _T_3678 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8728 = _T_8727 | _T_8483; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8485 = _T_3682 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8729 = _T_8728 | _T_8485; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8487 = _T_3686 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8730 = _T_8729 | _T_8487; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8489 = _T_3690 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8731 = _T_8730 | _T_8489; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8491 = _T_3694 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8732 = _T_8731 | _T_8491; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8493 = _T_3698 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8733 = _T_8732 | _T_8493; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8495 = _T_3702 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8734 = _T_8733 | _T_8495; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8497 = _T_3706 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8735 = _T_8734 | _T_8497; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8499 = _T_3710 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8736 = _T_8735 | _T_8499; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8501 = _T_3714 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8737 = _T_8736 | _T_8501; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8503 = _T_3718 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8738 = _T_8737 | _T_8503; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8505 = _T_3722 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8739 = _T_8738 | _T_8505; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8507 = _T_3726 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8740 = _T_8739 | _T_8507; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8509 = _T_3730 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8741 = _T_8740 | _T_8509; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8511 = _T_3734 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8742 = _T_8741 | _T_8511; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8513 = _T_3738 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8743 = _T_8742 | _T_8513; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8515 = _T_3742 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8744 = _T_8743 | _T_8515; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8517 = _T_3746 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8745 = _T_8744 | _T_8517; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8519 = _T_3750 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8746 = _T_8745 | _T_8519; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8521 = _T_3754 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8747 = _T_8746 | _T_8521; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8523 = _T_3758 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8748 = _T_8747 | _T_8523; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_8525 = _T_3762 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8749 = _T_8748 | _T_8525; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_8527 = _T_3766 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8750 = _T_8749 | _T_8527; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_8529 = _T_3770 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8751 = _T_8750 | _T_8529; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_8531 = _T_3774 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8752 = _T_8751 | _T_8531; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_8533 = _T_3778 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8753 = _T_8752 | _T_8533; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_8535 = _T_3782 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8754 = _T_8753 | _T_8535; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_8537 = _T_3786 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8755 = _T_8754 | _T_8537; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_8539 = _T_3790 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8756 = _T_8755 | _T_8539; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_8541 = _T_3794 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8757 = _T_8756 | _T_8541; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_8543 = _T_3798 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8758 = _T_8757 | _T_8543; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_8545 = _T_3802 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8759 = _T_8758 | _T_8545; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_8547 = _T_3806 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8760 = _T_8759 | _T_8547; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_8549 = _T_3810 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8761 = _T_8760 | _T_8549; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_8551 = _T_3814 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8762 = _T_8761 | _T_8551; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_8553 = _T_3818 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8763 = _T_8762 | _T_8553; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_8555 = _T_3822 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8764 = _T_8763 | _T_8555; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_8557 = _T_3826 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8765 = _T_8764 | _T_8557; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_8559 = _T_3830 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8766 = _T_8765 | _T_8559; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_8561 = _T_3834 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8767 = _T_8766 | _T_8561; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_8563 = _T_3838 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8768 = _T_8767 | _T_8563; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_8565 = _T_3842 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8769 = _T_8768 | _T_8565; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_8567 = _T_3846 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8770 = _T_8769 | _T_8567; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_8569 = _T_3850 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8771 = _T_8770 | _T_8569; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_8571 = _T_3854 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8772 = _T_8771 | _T_8571; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_8573 = _T_3858 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8773 = _T_8772 | _T_8573; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_8575 = _T_3862 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8774 = _T_8773 | _T_8575; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_8577 = _T_3866 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8775 = _T_8774 | _T_8577; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_8579 = _T_3870 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8776 = _T_8775 | _T_8579; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_8581 = _T_3874 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8777 = _T_8776 | _T_8581; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_8583 = _T_3878 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8778 = _T_8777 | _T_8583; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_8585 = _T_3882 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8779 = _T_8778 | _T_8585; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_8587 = _T_3886 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8780 = _T_8779 | _T_8587; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_8589 = _T_3890 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8781 = _T_8780 | _T_8589; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_8591 = _T_3894 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8782 = _T_8781 | _T_8591; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_8593 = _T_3898 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8783 = _T_8782 | _T_8593; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_8595 = _T_3902 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8784 = _T_8783 | _T_8595; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_8597 = _T_3906 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8785 = _T_8784 | _T_8597; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_8599 = _T_3910 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8786 = _T_8785 | _T_8599; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_8601 = _T_3914 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8787 = _T_8786 | _T_8601; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_8603 = _T_3918 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8788 = _T_8787 | _T_8603; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_8605 = _T_3922 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8789 = _T_8788 | _T_8605; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_8607 = _T_3926 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8790 = _T_8789 | _T_8607; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_8609 = _T_3930 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8791 = _T_8790 | _T_8609; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_8611 = _T_3934 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8792 = _T_8791 | _T_8611; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_8613 = _T_3938 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8793 = _T_8792 | _T_8613; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_8615 = _T_3942 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8794 = _T_8793 | _T_8615; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_8617 = _T_3946 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8795 = _T_8794 | _T_8617; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_8619 = _T_3950 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8796 = _T_8795 | _T_8619; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_8621 = _T_3954 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8797 = _T_8796 | _T_8621; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_8623 = _T_3958 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8798 = _T_8797 | _T_8623; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_8625 = _T_3962 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8799 = _T_8798 | _T_8625; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_8627 = _T_3966 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8800 = _T_8799 | _T_8627; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_8629 = _T_3970 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8801 = _T_8800 | _T_8629; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_8631 = _T_3974 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8802 = _T_8801 | _T_8631; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_8633 = _T_3978 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8803 = _T_8802 | _T_8633; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_8635 = _T_3982 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8804 = _T_8803 | _T_8635; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_8637 = _T_3986 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8805 = _T_8804 | _T_8637; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_8639 = _T_3990 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8806 = _T_8805 | _T_8639; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_8641 = _T_3994 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8807 = _T_8806 | _T_8641; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_8643 = _T_3998 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8808 = _T_8807 | _T_8643; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_8645 = _T_4002 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8809 = _T_8808 | _T_8645; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_8647 = _T_4006 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8810 = _T_8809 | _T_8647; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_8649 = _T_4010 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8811 = _T_8810 | _T_8649; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_8651 = _T_4014 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8812 = _T_8811 | _T_8651; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_8653 = _T_4018 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8813 = _T_8812 | _T_8653; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_8655 = _T_4022 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8814 = _T_8813 | _T_8655; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_8657 = _T_4026 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8815 = _T_8814 | _T_8657; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_8659 = _T_4030 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8816 = _T_8815 | _T_8659; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_8661 = _T_4034 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8817 = _T_8816 | _T_8661; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_8663 = _T_4038 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8818 = _T_8817 | _T_8663; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_8665 = _T_4042 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8819 = _T_8818 | _T_8665; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_8667 = _T_4046 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8820 = _T_8819 | _T_8667; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_8669 = _T_4050 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8821 = _T_8820 | _T_8669; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_8671 = _T_4054 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8822 = _T_8821 | _T_8671; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_8673 = _T_4058 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8823 = _T_8822 | _T_8673; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_8675 = _T_4062 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8824 = _T_8823 | _T_8675; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_8677 = _T_4066 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8825 = _T_8824 | _T_8677; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_8679 = _T_4070 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8826 = _T_8825 | _T_8679; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_8681 = _T_4074 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8827 = _T_8826 | _T_8681; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_8683 = _T_4078 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8828 = _T_8827 | _T_8683; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_8685 = _T_4082 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8829 = _T_8828 | _T_8685; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_8687 = _T_4086 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8830 = _T_8829 | _T_8687; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_8689 = _T_4090 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8831 = _T_8830 | _T_8689; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_8691 = _T_4094 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8832 = _T_8831 | _T_8691; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_8693 = _T_4098 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8833 = _T_8832 | _T_8693; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_8695 = _T_4102 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8834 = _T_8833 | _T_8695; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_8697 = _T_4106 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8835 = _T_8834 | _T_8697; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_8699 = _T_4110 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8836 = _T_8835 | _T_8699; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_8701 = _T_4114 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8837 = _T_8836 | _T_8701; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_8703 = _T_4118 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8838 = _T_8837 | _T_8703; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_8705 = _T_4122 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8839 = _T_8838 | _T_8705; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_8707 = _T_4126 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8840 = _T_8839 | _T_8707; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_8709 = _T_4130 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8841 = _T_8840 | _T_8709; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_8711 = _T_4134 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8842 = _T_8841 | _T_8711; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_8713 = _T_4138 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8843 = _T_8842 | _T_8713; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_8715 = _T_4142 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8844 = _T_8843 | _T_8715; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_8717 = _T_4146 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8845 = _T_8844 | _T_8717; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_8719 = _T_4150 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_8846 = _T_8845 | _T_8719; // @[el2_ifu_mem_ctl.scala 760:91]
  wire [1:0] ic_tag_valid_unq = {_T_9229,_T_8846}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 833:54]
  wire [1:0] _T_9268 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9269 = ic_debug_way_ff & _T_9268; // @[el2_ifu_mem_ctl.scala 814:67]
  wire [1:0] _T_9270 = ic_tag_valid_unq & _T_9269; // @[el2_ifu_mem_ctl.scala 814:48]
  wire  ic_debug_tag_val_rd_out = |_T_9270; // @[el2_ifu_mem_ctl.scala 814:115]
  wire [65:0] _T_365 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_366; // @[el2_ifu_mem_ctl.scala 362:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_1710; // @[el2_ifu_mem_ctl.scala 374:80]
  wire  _T_406 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 379:98]
  wire  sel_byp_data = _T_410 & _T_406; // @[el2_ifu_mem_ctl.scala 379:96]
  wire [63:0] _T_417 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_418 = _T_417 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 386:64]
  wire [63:0] _T_420 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_1272 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 455:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_786 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_834 = _T_786 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_789 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_835 = _T_789 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_850 = _T_834 | _T_835; // @[Mux.scala 27:72]
  wire  _T_792 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_836 = _T_792 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_851 = _T_850 | _T_836; // @[Mux.scala 27:72]
  wire  _T_795 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_837 = _T_795 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_852 = _T_851 | _T_837; // @[Mux.scala 27:72]
  wire  _T_798 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_838 = _T_798 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_853 = _T_852 | _T_838; // @[Mux.scala 27:72]
  wire  _T_801 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_839 = _T_801 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_854 = _T_853 | _T_839; // @[Mux.scala 27:72]
  wire  _T_804 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_840 = _T_804 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_855 = _T_854 | _T_840; // @[Mux.scala 27:72]
  wire  _T_807 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_841 = _T_807 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_856 = _T_855 | _T_841; // @[Mux.scala 27:72]
  wire  _T_810 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_842 = _T_810 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_857 = _T_856 | _T_842; // @[Mux.scala 27:72]
  wire  _T_813 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_843 = _T_813 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_858 = _T_857 | _T_843; // @[Mux.scala 27:72]
  wire  _T_816 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_844 = _T_816 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_859 = _T_858 | _T_844; // @[Mux.scala 27:72]
  wire  _T_819 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_845 = _T_819 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_860 = _T_859 | _T_845; // @[Mux.scala 27:72]
  wire  _T_822 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_846 = _T_822 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_861 = _T_860 | _T_846; // @[Mux.scala 27:72]
  wire  _T_825 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_847 = _T_825 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_862 = _T_861 | _T_847; // @[Mux.scala 27:72]
  wire  _T_828 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_848 = _T_828 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_863 = _T_862 | _T_848; // @[Mux.scala 27:72]
  wire  _T_831 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 452:73]
  wire [15:0] _T_849 = _T_831 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_864 = _T_863 | _T_849; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_866 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_914 = _T_866 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_869 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_915 = _T_869 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_930 = _T_914 | _T_915; // @[Mux.scala 27:72]
  wire  _T_872 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_916 = _T_872 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_931 = _T_930 | _T_916; // @[Mux.scala 27:72]
  wire  _T_875 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_917 = _T_875 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_932 = _T_931 | _T_917; // @[Mux.scala 27:72]
  wire  _T_878 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_918 = _T_878 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_933 = _T_932 | _T_918; // @[Mux.scala 27:72]
  wire  _T_881 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_919 = _T_881 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_934 = _T_933 | _T_919; // @[Mux.scala 27:72]
  wire  _T_884 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_920 = _T_884 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_935 = _T_934 | _T_920; // @[Mux.scala 27:72]
  wire  _T_887 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_921 = _T_887 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_936 = _T_935 | _T_921; // @[Mux.scala 27:72]
  wire  _T_890 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_922 = _T_890 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_937 = _T_936 | _T_922; // @[Mux.scala 27:72]
  wire  _T_893 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_923 = _T_893 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_938 = _T_937 | _T_923; // @[Mux.scala 27:72]
  wire  _T_896 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_924 = _T_896 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_939 = _T_938 | _T_924; // @[Mux.scala 27:72]
  wire  _T_899 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_925 = _T_899 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_940 = _T_939 | _T_925; // @[Mux.scala 27:72]
  wire  _T_902 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_926 = _T_902 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_941 = _T_940 | _T_926; // @[Mux.scala 27:72]
  wire  _T_905 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_927 = _T_905 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_942 = _T_941 | _T_927; // @[Mux.scala 27:72]
  wire  _T_908 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_928 = _T_908 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_943 = _T_942 | _T_928; // @[Mux.scala 27:72]
  wire  _T_911 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 452:179]
  wire [31:0] _T_929 = _T_911 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_944 = _T_943 | _T_929; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_946 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_994 = _T_946 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_949 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_995 = _T_949 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1010 = _T_994 | _T_995; // @[Mux.scala 27:72]
  wire  _T_952 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_996 = _T_952 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1011 = _T_1010 | _T_996; // @[Mux.scala 27:72]
  wire  _T_955 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_997 = _T_955 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1012 = _T_1011 | _T_997; // @[Mux.scala 27:72]
  wire  _T_958 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_998 = _T_958 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1013 = _T_1012 | _T_998; // @[Mux.scala 27:72]
  wire  _T_961 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_999 = _T_961 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1014 = _T_1013 | _T_999; // @[Mux.scala 27:72]
  wire  _T_964 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1000 = _T_964 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1015 = _T_1014 | _T_1000; // @[Mux.scala 27:72]
  wire  _T_967 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1001 = _T_967 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1016 = _T_1015 | _T_1001; // @[Mux.scala 27:72]
  wire  _T_970 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1002 = _T_970 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1017 = _T_1016 | _T_1002; // @[Mux.scala 27:72]
  wire  _T_973 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1003 = _T_973 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1018 = _T_1017 | _T_1003; // @[Mux.scala 27:72]
  wire  _T_976 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1004 = _T_976 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1019 = _T_1018 | _T_1004; // @[Mux.scala 27:72]
  wire  _T_979 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1005 = _T_979 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1020 = _T_1019 | _T_1005; // @[Mux.scala 27:72]
  wire  _T_982 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1006 = _T_982 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1021 = _T_1020 | _T_1006; // @[Mux.scala 27:72]
  wire  _T_985 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1007 = _T_985 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1022 = _T_1021 | _T_1007; // @[Mux.scala 27:72]
  wire  _T_988 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1008 = _T_988 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1023 = _T_1022 | _T_1008; // @[Mux.scala 27:72]
  wire  _T_991 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 452:285]
  wire [31:0] _T_1009 = _T_991 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1024 = _T_1023 | _T_1009; // @[Mux.scala 27:72]
  wire [79:0] _T_1027 = {_T_864,_T_944,_T_1024}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1028 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1076 = _T_1028 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1031 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1077 = _T_1031 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1092 = _T_1076 | _T_1077; // @[Mux.scala 27:72]
  wire  _T_1034 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1078 = _T_1034 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1093 = _T_1092 | _T_1078; // @[Mux.scala 27:72]
  wire  _T_1037 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1079 = _T_1037 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1094 = _T_1093 | _T_1079; // @[Mux.scala 27:72]
  wire  _T_1040 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1080 = _T_1040 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1095 = _T_1094 | _T_1080; // @[Mux.scala 27:72]
  wire  _T_1043 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1081 = _T_1043 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1096 = _T_1095 | _T_1081; // @[Mux.scala 27:72]
  wire  _T_1046 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1082 = _T_1046 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1097 = _T_1096 | _T_1082; // @[Mux.scala 27:72]
  wire  _T_1049 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1083 = _T_1049 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1098 = _T_1097 | _T_1083; // @[Mux.scala 27:72]
  wire  _T_1052 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1084 = _T_1052 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1099 = _T_1098 | _T_1084; // @[Mux.scala 27:72]
  wire  _T_1055 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1085 = _T_1055 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1100 = _T_1099 | _T_1085; // @[Mux.scala 27:72]
  wire  _T_1058 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1086 = _T_1058 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1101 = _T_1100 | _T_1086; // @[Mux.scala 27:72]
  wire  _T_1061 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1087 = _T_1061 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1102 = _T_1101 | _T_1087; // @[Mux.scala 27:72]
  wire  _T_1064 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1088 = _T_1064 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1103 = _T_1102 | _T_1088; // @[Mux.scala 27:72]
  wire  _T_1067 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1089 = _T_1067 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1104 = _T_1103 | _T_1089; // @[Mux.scala 27:72]
  wire  _T_1070 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1090 = _T_1070 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1105 = _T_1104 | _T_1090; // @[Mux.scala 27:72]
  wire  _T_1073 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 453:73]
  wire [15:0] _T_1091 = _T_1073 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1106 = _T_1105 | _T_1091; // @[Mux.scala 27:72]
  wire [31:0] _T_1156 = _T_786 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1157 = _T_789 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1172 = _T_1156 | _T_1157; // @[Mux.scala 27:72]
  wire [31:0] _T_1158 = _T_792 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1173 = _T_1172 | _T_1158; // @[Mux.scala 27:72]
  wire [31:0] _T_1159 = _T_795 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1174 = _T_1173 | _T_1159; // @[Mux.scala 27:72]
  wire [31:0] _T_1160 = _T_798 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1175 = _T_1174 | _T_1160; // @[Mux.scala 27:72]
  wire [31:0] _T_1161 = _T_801 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1176 = _T_1175 | _T_1161; // @[Mux.scala 27:72]
  wire [31:0] _T_1162 = _T_804 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1177 = _T_1176 | _T_1162; // @[Mux.scala 27:72]
  wire [31:0] _T_1163 = _T_807 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1178 = _T_1177 | _T_1163; // @[Mux.scala 27:72]
  wire [31:0] _T_1164 = _T_810 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1179 = _T_1178 | _T_1164; // @[Mux.scala 27:72]
  wire [31:0] _T_1165 = _T_813 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1180 = _T_1179 | _T_1165; // @[Mux.scala 27:72]
  wire [31:0] _T_1166 = _T_816 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1181 = _T_1180 | _T_1166; // @[Mux.scala 27:72]
  wire [31:0] _T_1167 = _T_819 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1182 = _T_1181 | _T_1167; // @[Mux.scala 27:72]
  wire [31:0] _T_1168 = _T_822 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1183 = _T_1182 | _T_1168; // @[Mux.scala 27:72]
  wire [31:0] _T_1169 = _T_825 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1184 = _T_1183 | _T_1169; // @[Mux.scala 27:72]
  wire [31:0] _T_1170 = _T_828 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1185 = _T_1184 | _T_1170; // @[Mux.scala 27:72]
  wire [31:0] _T_1171 = _T_831 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1186 = _T_1185 | _T_1171; // @[Mux.scala 27:72]
  wire [79:0] _T_1269 = {_T_1106,_T_1186,_T_944}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1272 ? _T_1027 : _T_1269; // @[el2_ifu_mem_ctl.scala 451:37]
  wire [79:0] _T_1274 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_1272 ? ic_byp_data_only_pre_new : _T_1274; // @[el2_ifu_mem_ctl.scala 455:30]
  wire [79:0] _GEN_793 = {{16'd0}, _T_420}; // @[el2_ifu_mem_ctl.scala 386:109]
  wire [79:0] _T_421 = _GEN_793 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 386:109]
  wire [79:0] _GEN_794 = {{16'd0}, _T_418}; // @[el2_ifu_mem_ctl.scala 386:83]
  wire [79:0] ic_premux_data = _GEN_794 | _T_421; // @[el2_ifu_mem_ctl.scala 386:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 393:38]
  wire [1:0] _T_430 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 397:8]
  wire [7:0] _T_527 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_532 = ic_miss_buff_data_error[0] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  _T_1778 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 629:47]
  wire  _T_1779 = _T_1778 & _T_13; // @[el2_ifu_mem_ctl.scala 629:50]
  wire  bus_ifu_wr_data_error = _T_1779 & miss_pending; // @[el2_ifu_mem_ctl.scala 629:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_532; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_536 = ic_miss_buff_data_error[1] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_536; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_540 = ic_miss_buff_data_error[2] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_540; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_544 = ic_miss_buff_data_error[3] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_544; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_548 = ic_miss_buff_data_error[4] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_548; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_552 = ic_miss_buff_data_error[5] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_552; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_556 = ic_miss_buff_data_error[6] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_556; // @[el2_ifu_mem_ctl.scala 417:72]
  wire  _T_560 = ic_miss_buff_data_error[7] & _T_498; // @[el2_ifu_mem_ctl.scala 418:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_560; // @[el2_ifu_mem_ctl.scala 417:72]
  wire [7:0] _T_567 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_1584 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1592 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 498:65]
  wire  _T_1593 = _T_1592 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 498:88]
  wire  _T_1595 = _T_1593 & _T_1706; // @[el2_ifu_mem_ctl.scala 498:112]
  wire  _T_1596 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1597 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 503:50]
  wire  _T_1599 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1605 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1607 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_1605 | _T_1607; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_1599 ? _T_1597 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_1596 ? _T_1597 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_1584 ? _T_1595 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_1584 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_1598 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 504:56]
  wire  _GEN_43 = _T_1596 & _T_1598; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_1584 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 489:58]
  wire  _T_1581 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 488:49]
  wire  _T_1586 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 497:87]
  wire  _T_1600 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 507:54]
  wire  _T_1601 = _T_1600 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 507:84]
  wire  _T_1610 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 528:66]
  wire  _T_1611 = io_dec_tlu_flush_err_wb & _T_1610; // @[el2_ifu_mem_ctl.scala 528:52]
  wire  _T_1613 = _T_1611 & _T_1706; // @[el2_ifu_mem_ctl.scala 528:81]
  wire  _T_1615 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 531:59]
  wire  _T_1616 = _T_1615 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 531:86]
  wire  _T_1630 = _T_1615 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 534:81]
  wire  _T_1631 = _T_1630 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 534:103]
  wire  _T_1632 = _T_1631 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 534:126]
  wire  _T_1652 = _T_1630 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 541:103]
  wire  _T_1659 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 546:62]
  wire  _T_1660 = io_dec_tlu_flush_lower_wb & _T_1659; // @[el2_ifu_mem_ctl.scala 546:60]
  wire  _T_1661 = _T_1660 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 546:88]
  wire  _T_1662 = _T_1661 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 546:115]
  wire  _GEN_50 = _T_1658 & _T_1616; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_1641 ? _T_1652 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_1641 | _T_1658; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_1614 ? _T_1632 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_1614 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_1609 ? _T_1613 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_1674 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 563:64]
  wire  _T_1676 = _T_1674 & _T_1706; // @[el2_ifu_mem_ctl.scala 563:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_1678 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 563:133]
  wire  _T_1679 = _T_1678 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 563:164]
  wire  _T_1680 = _T_1679 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 563:184]
  wire  _T_1681 = _T_1680 & miss_pending; // @[el2_ifu_mem_ctl.scala 563:204]
  wire  _T_1682 = ~_T_1681; // @[el2_ifu_mem_ctl.scala 563:112]
  wire  ifc_bus_ic_req_ff_in = _T_1676 & _T_1682; // @[el2_ifu_mem_ctl.scala 563:110]
  wire  _T_1683 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 564:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 595:45]
  wire  _T_1700 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 598:35]
  wire  _T_1701 = _T_1700 & miss_pending; // @[el2_ifu_mem_ctl.scala 598:53]
  wire  bus_cmd_sent = _T_1701 & _T_1706; // @[el2_ifu_mem_ctl.scala 598:68]
  wire [2:0] _T_1691 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1693 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1695 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 596:51]
  wire  _T_1721 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 606:73]
  wire  _T_1722 = _T_1707 & _T_1721; // @[el2_ifu_mem_ctl.scala 606:71]
  wire  _T_1724 = last_data_recieved_ff & _T_498; // @[el2_ifu_mem_ctl.scala 606:114]
  wire  last_data_recieved_in = _T_1722 | _T_1724; // @[el2_ifu_mem_ctl.scala 606:89]
  wire [2:0] _T_1730 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 611:45]
  wire  _T_1733 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 612:81]
  wire  _T_1734 = _T_1733 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 612:97]
  wire  _T_1736 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 614:48]
  wire  _T_1737 = _T_1736 & miss_pending; // @[el2_ifu_mem_ctl.scala 614:68]
  wire  bus_inc_cmd_beat_cnt = _T_1737 & _T_1706; // @[el2_ifu_mem_ctl.scala 614:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 616:57]
  wire  _T_1741 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 617:31]
  wire  _T_1742 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 617:71]
  wire  _T_1743 = _T_1742 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 617:87]
  wire  _T_1744 = ~_T_1743; // @[el2_ifu_mem_ctl.scala 617:55]
  wire  bus_hold_cmd_beat_cnt = _T_1741 & _T_1744; // @[el2_ifu_mem_ctl.scala 617:53]
  wire  _T_1745 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 618:46]
  wire  bus_cmd_beat_en = _T_1745 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 618:62]
  wire [2:0] _T_1748 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 620:46]
  wire [2:0] _T_1750 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1751 = bus_inc_cmd_beat_cnt ? _T_1748 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1752 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1754 = _T_1750 | _T_1751; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_1754 | _T_1752; // @[Mux.scala 27:72]
  wire  _T_1758 = _T_1734 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 621:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 632:62]
  wire  _T_1786 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 637:50]
  wire  _T_1787 = io_ifc_dma_access_ok & _T_1786; // @[el2_ifu_mem_ctl.scala 637:47]
  wire  _T_1788 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 637:70]
  wire  ifc_dma_access_ok_d = _T_1787 & _T_1788; // @[el2_ifu_mem_ctl.scala 637:68]
  wire  _T_1792 = _T_1787 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 638:72]
  wire  _T_1793 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 638:111]
  wire  _T_1794 = _T_1792 & _T_1793; // @[el2_ifu_mem_ctl.scala 638:97]
  wire  ifc_dma_access_q_ok = _T_1794 & _T_1788; // @[el2_ifu_mem_ctl.scala 638:127]
  wire  _T_1797 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 641:40]
  wire  _T_1798 = _T_1797 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 641:58]
  wire  _T_1801 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 642:60]
  wire  _T_1802 = _T_1797 & _T_1801; // @[el2_ifu_mem_ctl.scala 642:58]
  wire  _T_1803 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 642:104]
  wire [2:0] _T_1808 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_1914 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_1923 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_1914}; // @[el2_lib.scala 268:22]
  wire  _T_1924 = ^_T_1923; // @[el2_lib.scala 268:29]
  wire [8:0] _T_1932 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_1941 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_1932}; // @[el2_lib.scala 268:39]
  wire  _T_1942 = ^_T_1941; // @[el2_lib.scala 268:46]
  wire [8:0] _T_1950 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_1959 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_1950}; // @[el2_lib.scala 268:56]
  wire  _T_1960 = ^_T_1959; // @[el2_lib.scala 268:63]
  wire [6:0] _T_1966 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_1974 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_1966}; // @[el2_lib.scala 268:73]
  wire  _T_1975 = ^_T_1974; // @[el2_lib.scala 268:80]
  wire [14:0] _T_1989 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_1966}; // @[el2_lib.scala 268:90]
  wire  _T_1990 = ^_T_1989; // @[el2_lib.scala 268:97]
  wire [5:0] _T_1995 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_1996 = ^_T_1995; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2001 = {_T_1924,_T_1942,_T_1960,_T_1975,_T_1990,_T_1996}; // @[Cat.scala 29:58]
  wire  _T_2002 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2003 = ^_T_2001; // @[el2_lib.scala 269:23]
  wire  _T_2004 = _T_2002 ^ _T_2003; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2110 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2119 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2110}; // @[el2_lib.scala 268:22]
  wire  _T_2120 = ^_T_2119; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2128 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2137 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2128}; // @[el2_lib.scala 268:39]
  wire  _T_2138 = ^_T_2137; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2146 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2155 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2146}; // @[el2_lib.scala 268:56]
  wire  _T_2156 = ^_T_2155; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2162 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2170 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2162}; // @[el2_lib.scala 268:73]
  wire  _T_2171 = ^_T_2170; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2185 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2162}; // @[el2_lib.scala 268:90]
  wire  _T_2186 = ^_T_2185; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2191 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_2192 = ^_T_2191; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2197 = {_T_2120,_T_2138,_T_2156,_T_2171,_T_2186,_T_2192}; // @[Cat.scala 29:58]
  wire  _T_2198 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_2199 = ^_T_2197; // @[el2_lib.scala 269:23]
  wire  _T_2200 = _T_2198 ^ _T_2199; // @[el2_lib.scala 269:18]
  wire [6:0] _T_2201 = {_T_2200,_T_2120,_T_2138,_T_2156,_T_2171,_T_2186,_T_2192}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2004,_T_1924,_T_1942,_T_1960,_T_1975,_T_1990,_T_1996,_T_2201}; // @[Cat.scala 29:58]
  wire  _T_2203 = ~_T_1797; // @[el2_ifu_mem_ctl.scala 647:45]
  wire  _T_2204 = iccm_correct_ecc & _T_2203; // @[el2_ifu_mem_ctl.scala 647:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_2205 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_2212 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 661:53]
  wire  _T_2544 = _T_2456[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2542 = _T_2456[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2540 = _T_2456[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2538 = _T_2456[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2536 = _T_2456[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2534 = _T_2456[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2532 = _T_2456[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2530 = _T_2456[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2528 = _T_2456[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2526 = _T_2456[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2602 = {_T_2544,_T_2542,_T_2540,_T_2538,_T_2536,_T_2534,_T_2532,_T_2530,_T_2528,_T_2526}; // @[el2_lib.scala 310:69]
  wire  _T_2524 = _T_2456[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2522 = _T_2456[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2520 = _T_2456[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2518 = _T_2456[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2516 = _T_2456[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2514 = _T_2456[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2512 = _T_2456[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2510 = _T_2456[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2508 = _T_2456[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2506 = _T_2456[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2593 = {_T_2524,_T_2522,_T_2520,_T_2518,_T_2516,_T_2514,_T_2512,_T_2510,_T_2508,_T_2506}; // @[el2_lib.scala 310:69]
  wire  _T_2504 = _T_2456[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2502 = _T_2456[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2500 = _T_2456[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2498 = _T_2456[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2496 = _T_2456[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2494 = _T_2456[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2492 = _T_2456[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2490 = _T_2456[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2488 = _T_2456[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2486 = _T_2456[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2583 = {_T_2504,_T_2502,_T_2500,_T_2498,_T_2496,_T_2494,_T_2492,_T_2490,_T_2488,_T_2486}; // @[el2_lib.scala 310:69]
  wire  _T_2484 = _T_2456[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2482 = _T_2456[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2480 = _T_2456[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2478 = _T_2456[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2476 = _T_2456[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2474 = _T_2456[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2472 = _T_2456[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2470 = _T_2456[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2468 = _T_2456[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_2584 = {_T_2583,_T_2484,_T_2482,_T_2480,_T_2478,_T_2476,_T_2474,_T_2472,_T_2470,_T_2468}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_2604 = {_T_2602,_T_2593,_T_2584}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2559 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2565 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_2559}; // @[Cat.scala 29:58]
  wire [38:0] _T_2605 = _T_2604 ^ _T_2565; // @[el2_lib.scala 310:76]
  wire [38:0] _T_2606 = _T_2460 ? _T_2605 : _T_2565; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_2606[37:32],_T_2606[30:16],_T_2606[14:8],_T_2606[6:4],_T_2606[2]}; // @[Cat.scala 29:58]
  wire  _T_2929 = _T_2841[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2927 = _T_2841[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2925 = _T_2841[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2923 = _T_2841[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2921 = _T_2841[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2919 = _T_2841[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2917 = _T_2841[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2915 = _T_2841[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2913 = _T_2841[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2911 = _T_2841[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2987 = {_T_2929,_T_2927,_T_2925,_T_2923,_T_2921,_T_2919,_T_2917,_T_2915,_T_2913,_T_2911}; // @[el2_lib.scala 310:69]
  wire  _T_2909 = _T_2841[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2907 = _T_2841[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2905 = _T_2841[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2903 = _T_2841[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2901 = _T_2841[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2899 = _T_2841[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2897 = _T_2841[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2895 = _T_2841[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2893 = _T_2841[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2891 = _T_2841[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2978 = {_T_2909,_T_2907,_T_2905,_T_2903,_T_2901,_T_2899,_T_2897,_T_2895,_T_2893,_T_2891}; // @[el2_lib.scala 310:69]
  wire  _T_2889 = _T_2841[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2887 = _T_2841[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2885 = _T_2841[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2883 = _T_2841[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2881 = _T_2841[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2879 = _T_2841[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2877 = _T_2841[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2875 = _T_2841[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2873 = _T_2841[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2871 = _T_2841[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2968 = {_T_2889,_T_2887,_T_2885,_T_2883,_T_2881,_T_2879,_T_2877,_T_2875,_T_2873,_T_2871}; // @[el2_lib.scala 310:69]
  wire  _T_2869 = _T_2841[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2867 = _T_2841[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2865 = _T_2841[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2863 = _T_2841[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2861 = _T_2841[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2859 = _T_2841[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2857 = _T_2841[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2855 = _T_2841[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2853 = _T_2841[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_2969 = {_T_2968,_T_2869,_T_2867,_T_2865,_T_2863,_T_2861,_T_2859,_T_2857,_T_2855,_T_2853}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_2989 = {_T_2987,_T_2978,_T_2969}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2944 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2950 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_2944}; // @[Cat.scala 29:58]
  wire [38:0] _T_2990 = _T_2989 ^ _T_2950; // @[el2_lib.scala 310:76]
  wire [38:0] _T_2991 = _T_2845 ? _T_2990 : _T_2950; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_2991[37:32],_T_2991[30:16],_T_2991[14:8],_T_2991[6:4],_T_2991[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 653:35]
  wire  _T_2464 = ~_T_2456[6]; // @[el2_lib.scala 303:55]
  wire  _T_2465 = _T_2458 & _T_2464; // @[el2_lib.scala 303:53]
  wire  _T_2849 = ~_T_2841[6]; // @[el2_lib.scala 303:55]
  wire  _T_2850 = _T_2843 & _T_2849; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_2465,_T_2850}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 655:53]
  wire [63:0] _T_2216 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_2217 = {iccm_dma_rdata_1_muxed,_T_2606[37:32],_T_2606[30:16],_T_2606[14:8],_T_2606[6:4],_T_2606[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 657:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 658:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 663:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 667:70]
  wire  _T_2222 = _T_1797 & _T_1786; // @[el2_ifu_mem_ctl.scala 670:65]
  wire  _T_2225 = _T_2203 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 671:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_2226 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_2228 = _T_2225 ? {{1'd0}, _T_2226} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 671:8]
  wire [31:0] _T_2229 = _T_2222 ? io_dma_mem_addr : {{16'd0}, _T_2228}; // @[el2_ifu_mem_ctl.scala 670:25]
  wire  _T_2618 = _T_2456 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_2619 = _T_2606[38] ^ _T_2618; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_2619,_T_2606[31],_T_2606[15],_T_2606[7],_T_2606[3],_T_2606[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3003 = _T_2841 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3004 = _T_2991[38] ^ _T_3003; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3004,_T_2991[31],_T_2991[15],_T_2991[7],_T_2991[3],_T_2991[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3020 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 683:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 685:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 686:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 694:62]
  wire  _T_3028 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 688:76]
  wire  _T_3029 = io_iccm_rd_ecc_single_err & _T_3028; // @[el2_ifu_mem_ctl.scala 688:74]
  wire  _T_3031 = _T_3029 & _T_317; // @[el2_ifu_mem_ctl.scala 688:104]
  wire  iccm_ecc_write_status = _T_3031 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 688:127]
  wire  _T_3032 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 689:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3032 & _T_317; // @[el2_ifu_mem_ctl.scala 689:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 693:51]
  wire [13:0] _T_3037 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 692:102]
  wire [38:0] _T_3041 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3046 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 697:41]
  wire  _T_3047 = io_ifc_fetch_req_bf & _T_3046; // @[el2_ifu_mem_ctl.scala 697:39]
  wire  _T_3048 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 697:72]
  wire  _T_3049 = _T_3047 & _T_3048; // @[el2_ifu_mem_ctl.scala 697:70]
  wire  _T_3051 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 698:34]
  wire  _T_3052 = _T_1392 & _T_3051; // @[el2_ifu_mem_ctl.scala 698:32]
  wire  _T_3055 = _T_1408 & _T_3051; // @[el2_ifu_mem_ctl.scala 699:37]
  wire  _T_3056 = _T_3052 | _T_3055; // @[el2_ifu_mem_ctl.scala 698:88]
  wire  _T_3057 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 700:19]
  wire  _T_3059 = _T_3057 & _T_3051; // @[el2_ifu_mem_ctl.scala 700:41]
  wire  _T_3060 = _T_3056 | _T_3059; // @[el2_ifu_mem_ctl.scala 699:88]
  wire  _T_3061 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 701:19]
  wire  _T_3063 = _T_3061 & _T_3051; // @[el2_ifu_mem_ctl.scala 701:35]
  wire  _T_3064 = _T_3060 | _T_3063; // @[el2_ifu_mem_ctl.scala 700:88]
  wire  _T_3067 = _T_1407 & _T_3051; // @[el2_ifu_mem_ctl.scala 702:38]
  wire  _T_3068 = _T_3064 | _T_3067; // @[el2_ifu_mem_ctl.scala 701:88]
  wire  _T_3070 = _T_1408 & miss_state_en; // @[el2_ifu_mem_ctl.scala 703:37]
  wire  _T_3071 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 703:71]
  wire  _T_3072 = _T_3070 & _T_3071; // @[el2_ifu_mem_ctl.scala 703:54]
  wire  _T_3073 = _T_3068 | _T_3072; // @[el2_ifu_mem_ctl.scala 702:57]
  wire  _T_3074 = ~_T_3073; // @[el2_ifu_mem_ctl.scala 698:5]
  wire  _T_3075 = _T_3049 & _T_3074; // @[el2_ifu_mem_ctl.scala 697:96]
  wire  _T_3076 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 704:28]
  wire  _T_3078 = _T_3076 & _T_3046; // @[el2_ifu_mem_ctl.scala 704:50]
  wire  _T_3080 = _T_3078 & _T_3048; // @[el2_ifu_mem_ctl.scala 704:81]
  wire  _T_3089 = ~_T_108; // @[el2_ifu_mem_ctl.scala 707:106]
  wire  _T_3090 = _T_1392 & _T_3089; // @[el2_ifu_mem_ctl.scala 707:104]
  wire  _T_3091 = _T_1408 | _T_3090; // @[el2_ifu_mem_ctl.scala 707:77]
  wire  _T_3095 = ~_T_51; // @[el2_ifu_mem_ctl.scala 707:172]
  wire  _T_3096 = _T_3091 & _T_3095; // @[el2_ifu_mem_ctl.scala 707:170]
  wire  _T_3097 = ~_T_3096; // @[el2_ifu_mem_ctl.scala 707:44]
  wire  _T_3101 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 710:64]
  wire  _T_3102 = ~_T_3101; // @[el2_ifu_mem_ctl.scala 710:50]
  wire  _T_3103 = _T_276 & _T_3102; // @[el2_ifu_mem_ctl.scala 710:48]
  wire  _T_3104 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 710:81]
  wire  ic_valid = _T_3103 & _T_3104; // @[el2_ifu_mem_ctl.scala 710:79]
  wire  _T_3106 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 711:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 714:14]
  wire  _T_3109 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 717:74]
  wire  _T_9251 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 791:45]
  wire  way_status_wr_en = _T_9251 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 791:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3109; // @[el2_ifu_mem_ctl.scala 717:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 719:14]
  wire [2:0] _T_3113 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 723:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 787:41]
  wire  way_status_new = _T_9251 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 790:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 725:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 727:132]
  wire  _T_3130 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3131 = _T_3130 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3132 = _T_3131 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3134 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3135 = _T_3134 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3136 = _T_3135 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3138 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3139 = _T_3138 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3140 = _T_3139 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3142 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3143 = _T_3142 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3144 = _T_3143 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3146 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3147 = _T_3146 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3148 = _T_3147 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3150 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3151 = _T_3150 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3152 = _T_3151 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3154 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3155 = _T_3154 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3156 = _T_3155 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3158 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 731:93]
  wire  _T_3159 = _T_3158 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 731:102]
  wire  _T_3160 = _T_3159 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3164 = _T_3131 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3168 = _T_3135 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3172 = _T_3139 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3176 = _T_3143 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3180 = _T_3147 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3184 = _T_3151 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3188 = _T_3155 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3192 = _T_3159 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3196 = _T_3131 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3200 = _T_3135 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3204 = _T_3139 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3208 = _T_3143 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3212 = _T_3147 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3216 = _T_3151 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3220 = _T_3155 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3224 = _T_3159 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3228 = _T_3131 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3232 = _T_3135 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3236 = _T_3139 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3240 = _T_3143 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3244 = _T_3147 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3248 = _T_3151 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3252 = _T_3155 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3256 = _T_3159 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3260 = _T_3131 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3264 = _T_3135 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3268 = _T_3139 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3272 = _T_3143 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3276 = _T_3147 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3280 = _T_3151 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3284 = _T_3155 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3288 = _T_3159 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3292 = _T_3131 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3296 = _T_3135 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3300 = _T_3139 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3304 = _T_3143 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3308 = _T_3147 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3312 = _T_3151 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3316 = _T_3155 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3320 = _T_3159 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3324 = _T_3131 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3328 = _T_3135 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3332 = _T_3139 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3336 = _T_3143 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3340 = _T_3147 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3344 = _T_3151 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3348 = _T_3155 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3352 = _T_3159 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3356 = _T_3131 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3360 = _T_3135 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3364 = _T_3139 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3368 = _T_3143 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3372 = _T_3147 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3376 = _T_3151 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3380 = _T_3155 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3384 = _T_3159 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3388 = _T_3131 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3392 = _T_3135 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3396 = _T_3139 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3400 = _T_3143 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3404 = _T_3147 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3408 = _T_3151 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3412 = _T_3155 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3416 = _T_3159 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3420 = _T_3131 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3424 = _T_3135 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3428 = _T_3139 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3432 = _T_3143 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3436 = _T_3147 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3440 = _T_3151 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3444 = _T_3155 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3448 = _T_3159 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3452 = _T_3131 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3456 = _T_3135 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3460 = _T_3139 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3464 = _T_3143 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3468 = _T_3147 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3472 = _T_3151 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3476 = _T_3155 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3480 = _T_3159 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3484 = _T_3131 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3488 = _T_3135 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3492 = _T_3139 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3496 = _T_3143 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3500 = _T_3147 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3504 = _T_3151 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3508 = _T_3155 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3512 = _T_3159 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3516 = _T_3131 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3520 = _T_3135 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3524 = _T_3139 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3528 = _T_3143 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3532 = _T_3147 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3536 = _T_3151 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3540 = _T_3155 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3544 = _T_3159 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3548 = _T_3131 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3552 = _T_3135 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3556 = _T_3139 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3560 = _T_3143 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3564 = _T_3147 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3568 = _T_3151 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3572 = _T_3155 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3576 = _T_3159 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3580 = _T_3131 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3584 = _T_3135 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3588 = _T_3139 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3592 = _T_3143 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3596 = _T_3147 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3600 = _T_3151 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3604 = _T_3155 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3608 = _T_3159 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3612 = _T_3131 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3616 = _T_3135 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3620 = _T_3139 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3624 = _T_3143 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3628 = _T_3147 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3632 = _T_3151 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3636 = _T_3155 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_3640 = _T_3159 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 731:124]
  wire  _T_9257 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 794:84]
  wire  _T_9258 = _T_9257 & miss_pending; // @[el2_ifu_mem_ctl.scala 794:108]
  wire  bus_wren_last_1 = _T_9258 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 794:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_9260 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 796:73]
  wire  _T_9255 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 794:84]
  wire  _T_9256 = _T_9255 & miss_pending; // @[el2_ifu_mem_ctl.scala 794:108]
  wire  bus_wren_last_0 = _T_9256 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 794:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_9259 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 796:73]
  wire [1:0] ifu_tag_wren = {_T_9260,_T_9259}; // @[Cat.scala 29:58]
  wire [1:0] _T_9294 = _T_3109 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9294 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 829:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 740:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 742:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 746:14]
  wire  _T_4289 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4291 = _T_4289 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4293 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4295 = _T_4293 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4296 = _T_4291 | _T_4295; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4297 = _T_4296 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4301 = _T_4289 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4305 = _T_4293 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4306 = _T_4301 | _T_4305; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4307 = _T_4306 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_0 = {_T_4297,_T_4307}; // @[Cat.scala 29:58]
  wire  _T_4309 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4311 = _T_4309 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4313 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4315 = _T_4313 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4316 = _T_4311 | _T_4315; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4317 = _T_4316 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4321 = _T_4309 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4325 = _T_4313 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4326 = _T_4321 | _T_4325; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4327 = _T_4326 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_1 = {_T_4317,_T_4327}; // @[Cat.scala 29:58]
  wire  _T_4329 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4331 = _T_4329 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4333 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4335 = _T_4333 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4336 = _T_4331 | _T_4335; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4337 = _T_4336 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4341 = _T_4329 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4345 = _T_4333 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4346 = _T_4341 | _T_4345; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4347 = _T_4346 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_2 = {_T_4337,_T_4347}; // @[Cat.scala 29:58]
  wire  _T_4349 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 750:82]
  wire  _T_4351 = _T_4349 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4353 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 751:74]
  wire  _T_4355 = _T_4353 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4356 = _T_4351 | _T_4355; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4357 = _T_4356 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire  _T_4361 = _T_4349 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 750:91]
  wire  _T_4365 = _T_4353 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 751:83]
  wire  _T_4366 = _T_4361 | _T_4365; // @[el2_ifu_mem_ctl.scala 750:113]
  wire  _T_4367 = _T_4366 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 751:106]
  wire [1:0] tag_valid_clken_3 = {_T_4357,_T_4367}; // @[Cat.scala 29:58]
  wire  _T_4370 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 756:64]
  wire  _T_4371 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 756:91]
  wire  _T_4372 = _T_4370 & _T_4371; // @[el2_ifu_mem_ctl.scala 756:89]
  wire  _T_4375 = _T_3642 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4376 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4378 = _T_4376 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4380 = _T_4378 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4381 = _T_4375 | _T_4380; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4391 = _T_3646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4392 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4394 = _T_4392 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4396 = _T_4394 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4397 = _T_4391 | _T_4396; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4407 = _T_3650 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4408 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4410 = _T_4408 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4412 = _T_4410 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4413 = _T_4407 | _T_4412; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4423 = _T_3654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4424 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4426 = _T_4424 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4428 = _T_4426 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4429 = _T_4423 | _T_4428; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4439 = _T_3658 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4440 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4442 = _T_4440 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4444 = _T_4442 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4445 = _T_4439 | _T_4444; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4455 = _T_3662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4456 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4458 = _T_4456 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4460 = _T_4458 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4461 = _T_4455 | _T_4460; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4471 = _T_3666 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4472 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4474 = _T_4472 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4476 = _T_4474 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4477 = _T_4471 | _T_4476; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4487 = _T_3670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4488 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4490 = _T_4488 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4492 = _T_4490 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4493 = _T_4487 | _T_4492; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4503 = _T_3674 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4504 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4506 = _T_4504 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4508 = _T_4506 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4509 = _T_4503 | _T_4508; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4519 = _T_3678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4520 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4522 = _T_4520 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4524 = _T_4522 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4525 = _T_4519 | _T_4524; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4535 = _T_3682 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4536 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4538 = _T_4536 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4540 = _T_4538 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4541 = _T_4535 | _T_4540; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4551 = _T_3686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4552 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4554 = _T_4552 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4556 = _T_4554 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4557 = _T_4551 | _T_4556; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4567 = _T_3690 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4568 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4570 = _T_4568 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4572 = _T_4570 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4573 = _T_4567 | _T_4572; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4583 = _T_3694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4584 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4586 = _T_4584 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4588 = _T_4586 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4589 = _T_4583 | _T_4588; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4599 = _T_3698 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4600 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4602 = _T_4600 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4604 = _T_4602 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4605 = _T_4599 | _T_4604; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4615 = _T_3702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4616 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4618 = _T_4616 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4620 = _T_4618 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4621 = _T_4615 | _T_4620; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4631 = _T_3706 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4632 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4634 = _T_4632 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4636 = _T_4634 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4637 = _T_4631 | _T_4636; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4647 = _T_3710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4648 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4650 = _T_4648 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4652 = _T_4650 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4653 = _T_4647 | _T_4652; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4663 = _T_3714 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4664 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4666 = _T_4664 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4668 = _T_4666 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4669 = _T_4663 | _T_4668; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4679 = _T_3718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4680 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4682 = _T_4680 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4684 = _T_4682 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4685 = _T_4679 | _T_4684; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4695 = _T_3722 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4696 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4698 = _T_4696 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4700 = _T_4698 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4701 = _T_4695 | _T_4700; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4711 = _T_3726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4712 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4714 = _T_4712 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4716 = _T_4714 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4717 = _T_4711 | _T_4716; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4727 = _T_3730 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4728 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4730 = _T_4728 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4732 = _T_4730 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4733 = _T_4727 | _T_4732; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4743 = _T_3734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4744 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4746 = _T_4744 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4748 = _T_4746 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4749 = _T_4743 | _T_4748; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4759 = _T_3738 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4760 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4762 = _T_4760 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4764 = _T_4762 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4765 = _T_4759 | _T_4764; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4775 = _T_3742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4776 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4778 = _T_4776 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4780 = _T_4778 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4781 = _T_4775 | _T_4780; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4791 = _T_3746 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4792 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4794 = _T_4792 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4796 = _T_4794 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4797 = _T_4791 | _T_4796; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4807 = _T_3750 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4808 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4810 = _T_4808 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4812 = _T_4810 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4813 = _T_4807 | _T_4812; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4823 = _T_3754 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4824 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4826 = _T_4824 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4828 = _T_4826 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4829 = _T_4823 | _T_4828; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4839 = _T_3758 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4840 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4842 = _T_4840 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4844 = _T_4842 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4845 = _T_4839 | _T_4844; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4855 = _T_3762 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4856 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4858 = _T_4856 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4860 = _T_4858 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4861 = _T_4855 | _T_4860; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4871 = _T_3766 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4872 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_4874 = _T_4872 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4876 = _T_4874 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4877 = _T_4871 | _T_4876; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4887 = _T_3642 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4890 = _T_4376 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4892 = _T_4890 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4893 = _T_4887 | _T_4892; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4903 = _T_3646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4906 = _T_4392 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4908 = _T_4906 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4909 = _T_4903 | _T_4908; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4919 = _T_3650 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4922 = _T_4408 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4924 = _T_4922 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4925 = _T_4919 | _T_4924; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4935 = _T_3654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4938 = _T_4424 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4940 = _T_4938 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4941 = _T_4935 | _T_4940; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4951 = _T_3658 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4954 = _T_4440 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4956 = _T_4954 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4957 = _T_4951 | _T_4956; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4967 = _T_3662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4970 = _T_4456 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4972 = _T_4970 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4973 = _T_4967 | _T_4972; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4983 = _T_3666 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_4986 = _T_4472 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_4988 = _T_4986 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_4989 = _T_4983 | _T_4988; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_4999 = _T_3670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5002 = _T_4488 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5004 = _T_5002 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5005 = _T_4999 | _T_5004; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5015 = _T_3674 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5018 = _T_4504 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5020 = _T_5018 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5021 = _T_5015 | _T_5020; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5031 = _T_3678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5034 = _T_4520 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5036 = _T_5034 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5037 = _T_5031 | _T_5036; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5047 = _T_3682 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5050 = _T_4536 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5052 = _T_5050 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5053 = _T_5047 | _T_5052; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5063 = _T_3686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5066 = _T_4552 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5068 = _T_5066 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5069 = _T_5063 | _T_5068; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5079 = _T_3690 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5082 = _T_4568 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5084 = _T_5082 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5085 = _T_5079 | _T_5084; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5095 = _T_3694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5098 = _T_4584 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5100 = _T_5098 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5101 = _T_5095 | _T_5100; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5111 = _T_3698 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5114 = _T_4600 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5116 = _T_5114 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5117 = _T_5111 | _T_5116; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5127 = _T_3702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5130 = _T_4616 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5132 = _T_5130 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5133 = _T_5127 | _T_5132; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5143 = _T_3706 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5146 = _T_4632 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5148 = _T_5146 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5149 = _T_5143 | _T_5148; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5159 = _T_3710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5162 = _T_4648 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5164 = _T_5162 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5165 = _T_5159 | _T_5164; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5175 = _T_3714 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5178 = _T_4664 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5180 = _T_5178 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5181 = _T_5175 | _T_5180; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5191 = _T_3718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5194 = _T_4680 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5196 = _T_5194 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5197 = _T_5191 | _T_5196; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5207 = _T_3722 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5210 = _T_4696 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5212 = _T_5210 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5213 = _T_5207 | _T_5212; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5223 = _T_3726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5226 = _T_4712 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5228 = _T_5226 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5229 = _T_5223 | _T_5228; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5239 = _T_3730 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5242 = _T_4728 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5244 = _T_5242 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5245 = _T_5239 | _T_5244; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5255 = _T_3734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5258 = _T_4744 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5260 = _T_5258 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5261 = _T_5255 | _T_5260; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5271 = _T_3738 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5274 = _T_4760 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5276 = _T_5274 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5277 = _T_5271 | _T_5276; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5287 = _T_3742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5290 = _T_4776 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5292 = _T_5290 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5293 = _T_5287 | _T_5292; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5303 = _T_3746 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5306 = _T_4792 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5308 = _T_5306 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5309 = _T_5303 | _T_5308; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5319 = _T_3750 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5322 = _T_4808 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5324 = _T_5322 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5325 = _T_5319 | _T_5324; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5335 = _T_3754 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5338 = _T_4824 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5340 = _T_5338 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5341 = _T_5335 | _T_5340; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5351 = _T_3758 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5354 = _T_4840 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5356 = _T_5354 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5357 = _T_5351 | _T_5356; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5367 = _T_3762 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5370 = _T_4856 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5372 = _T_5370 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5373 = _T_5367 | _T_5372; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5383 = _T_3766 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5386 = _T_4872 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5388 = _T_5386 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5389 = _T_5383 | _T_5388; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5399 = _T_3770 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5400 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5402 = _T_5400 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5404 = _T_5402 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5405 = _T_5399 | _T_5404; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5415 = _T_3774 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5416 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5418 = _T_5416 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5420 = _T_5418 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5421 = _T_5415 | _T_5420; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5431 = _T_3778 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5432 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5434 = _T_5432 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5436 = _T_5434 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5437 = _T_5431 | _T_5436; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5447 = _T_3782 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5448 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5450 = _T_5448 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5452 = _T_5450 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5453 = _T_5447 | _T_5452; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5463 = _T_3786 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5464 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5466 = _T_5464 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5468 = _T_5466 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5469 = _T_5463 | _T_5468; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5479 = _T_3790 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5480 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5482 = _T_5480 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5484 = _T_5482 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5485 = _T_5479 | _T_5484; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5495 = _T_3794 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5496 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5498 = _T_5496 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5500 = _T_5498 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5501 = _T_5495 | _T_5500; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5511 = _T_3798 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5512 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5514 = _T_5512 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5516 = _T_5514 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5517 = _T_5511 | _T_5516; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5527 = _T_3802 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5528 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5530 = _T_5528 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5532 = _T_5530 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5533 = _T_5527 | _T_5532; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5543 = _T_3806 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5544 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5546 = _T_5544 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5548 = _T_5546 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5549 = _T_5543 | _T_5548; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5559 = _T_3810 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5560 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5562 = _T_5560 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5564 = _T_5562 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5565 = _T_5559 | _T_5564; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5575 = _T_3814 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5576 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5578 = _T_5576 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5580 = _T_5578 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5581 = _T_5575 | _T_5580; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5591 = _T_3818 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5592 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5594 = _T_5592 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5596 = _T_5594 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5597 = _T_5591 | _T_5596; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5607 = _T_3822 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5608 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5610 = _T_5608 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5612 = _T_5610 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5613 = _T_5607 | _T_5612; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5623 = _T_3826 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5624 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5626 = _T_5624 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5628 = _T_5626 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5629 = _T_5623 | _T_5628; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5639 = _T_3830 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5640 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5642 = _T_5640 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5644 = _T_5642 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5645 = _T_5639 | _T_5644; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5655 = _T_3834 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5656 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5658 = _T_5656 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5660 = _T_5658 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5661 = _T_5655 | _T_5660; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5671 = _T_3838 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5672 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5674 = _T_5672 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5676 = _T_5674 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5677 = _T_5671 | _T_5676; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5687 = _T_3842 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5688 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5690 = _T_5688 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5692 = _T_5690 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5693 = _T_5687 | _T_5692; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5703 = _T_3846 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5704 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5706 = _T_5704 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5708 = _T_5706 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5709 = _T_5703 | _T_5708; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5719 = _T_3850 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5720 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5722 = _T_5720 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5724 = _T_5722 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5725 = _T_5719 | _T_5724; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5735 = _T_3854 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5736 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5738 = _T_5736 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5740 = _T_5738 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5741 = _T_5735 | _T_5740; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5751 = _T_3858 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5752 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5754 = _T_5752 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5756 = _T_5754 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5757 = _T_5751 | _T_5756; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5767 = _T_3862 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5768 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5770 = _T_5768 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5772 = _T_5770 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5773 = _T_5767 | _T_5772; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5783 = _T_3866 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5784 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5786 = _T_5784 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5788 = _T_5786 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5789 = _T_5783 | _T_5788; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5799 = _T_3870 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5800 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5802 = _T_5800 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5804 = _T_5802 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5805 = _T_5799 | _T_5804; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5815 = _T_3874 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5816 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5818 = _T_5816 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5820 = _T_5818 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5821 = _T_5815 | _T_5820; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5831 = _T_3878 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5832 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5834 = _T_5832 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5836 = _T_5834 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5837 = _T_5831 | _T_5836; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5847 = _T_3882 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5848 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5850 = _T_5848 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5852 = _T_5850 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5853 = _T_5847 | _T_5852; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5863 = _T_3886 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5864 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5866 = _T_5864 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5868 = _T_5866 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5869 = _T_5863 | _T_5868; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5879 = _T_3890 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5880 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5882 = _T_5880 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5884 = _T_5882 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5885 = _T_5879 | _T_5884; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5895 = _T_3894 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5896 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_5898 = _T_5896 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5900 = _T_5898 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5901 = _T_5895 | _T_5900; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5911 = _T_3770 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5914 = _T_5400 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5916 = _T_5914 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5917 = _T_5911 | _T_5916; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5927 = _T_3774 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5930 = _T_5416 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5932 = _T_5930 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5933 = _T_5927 | _T_5932; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5943 = _T_3778 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5946 = _T_5432 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5948 = _T_5946 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5949 = _T_5943 | _T_5948; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5959 = _T_3782 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5962 = _T_5448 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5964 = _T_5962 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5965 = _T_5959 | _T_5964; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5975 = _T_3786 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5978 = _T_5464 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5980 = _T_5978 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5981 = _T_5975 | _T_5980; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_5991 = _T_3790 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_5994 = _T_5480 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_5996 = _T_5994 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_5997 = _T_5991 | _T_5996; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6007 = _T_3794 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6010 = _T_5496 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6012 = _T_6010 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6013 = _T_6007 | _T_6012; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6023 = _T_3798 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6026 = _T_5512 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6028 = _T_6026 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6029 = _T_6023 | _T_6028; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6039 = _T_3802 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6042 = _T_5528 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6044 = _T_6042 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6045 = _T_6039 | _T_6044; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6055 = _T_3806 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6058 = _T_5544 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6060 = _T_6058 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6061 = _T_6055 | _T_6060; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6071 = _T_3810 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6074 = _T_5560 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6076 = _T_6074 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6077 = _T_6071 | _T_6076; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6087 = _T_3814 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6090 = _T_5576 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6092 = _T_6090 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6093 = _T_6087 | _T_6092; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6103 = _T_3818 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6106 = _T_5592 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6108 = _T_6106 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6109 = _T_6103 | _T_6108; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6119 = _T_3822 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6122 = _T_5608 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6124 = _T_6122 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6125 = _T_6119 | _T_6124; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6135 = _T_3826 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6138 = _T_5624 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6140 = _T_6138 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6141 = _T_6135 | _T_6140; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6151 = _T_3830 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6154 = _T_5640 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6156 = _T_6154 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6157 = _T_6151 | _T_6156; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6167 = _T_3834 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6170 = _T_5656 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6172 = _T_6170 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6173 = _T_6167 | _T_6172; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6183 = _T_3838 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6186 = _T_5672 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6188 = _T_6186 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6189 = _T_6183 | _T_6188; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6199 = _T_3842 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6202 = _T_5688 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6204 = _T_6202 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6205 = _T_6199 | _T_6204; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6215 = _T_3846 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6218 = _T_5704 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6220 = _T_6218 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6221 = _T_6215 | _T_6220; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6231 = _T_3850 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6234 = _T_5720 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6236 = _T_6234 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6237 = _T_6231 | _T_6236; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6247 = _T_3854 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6250 = _T_5736 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6252 = _T_6250 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6253 = _T_6247 | _T_6252; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6263 = _T_3858 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6266 = _T_5752 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6268 = _T_6266 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6269 = _T_6263 | _T_6268; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6279 = _T_3862 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6282 = _T_5768 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6284 = _T_6282 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6285 = _T_6279 | _T_6284; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6295 = _T_3866 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6298 = _T_5784 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6300 = _T_6298 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6301 = _T_6295 | _T_6300; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6311 = _T_3870 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6314 = _T_5800 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6316 = _T_6314 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6317 = _T_6311 | _T_6316; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6327 = _T_3874 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6330 = _T_5816 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6332 = _T_6330 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6333 = _T_6327 | _T_6332; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6343 = _T_3878 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6346 = _T_5832 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6348 = _T_6346 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6349 = _T_6343 | _T_6348; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6359 = _T_3882 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6362 = _T_5848 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6364 = _T_6362 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6365 = _T_6359 | _T_6364; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6375 = _T_3886 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6378 = _T_5864 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6380 = _T_6378 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6381 = _T_6375 | _T_6380; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6391 = _T_3890 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6394 = _T_5880 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6396 = _T_6394 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6397 = _T_6391 | _T_6396; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6407 = _T_3894 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6410 = _T_5896 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6412 = _T_6410 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6413 = _T_6407 | _T_6412; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6423 = _T_3898 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6424 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6426 = _T_6424 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6428 = _T_6426 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6429 = _T_6423 | _T_6428; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6439 = _T_3902 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6440 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6442 = _T_6440 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6444 = _T_6442 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6445 = _T_6439 | _T_6444; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6455 = _T_3906 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6456 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6458 = _T_6456 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6460 = _T_6458 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6461 = _T_6455 | _T_6460; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6471 = _T_3910 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6472 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6474 = _T_6472 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6476 = _T_6474 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6477 = _T_6471 | _T_6476; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6487 = _T_3914 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6488 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6490 = _T_6488 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6492 = _T_6490 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6493 = _T_6487 | _T_6492; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6503 = _T_3918 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6504 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6506 = _T_6504 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6508 = _T_6506 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6509 = _T_6503 | _T_6508; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6519 = _T_3922 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6520 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6522 = _T_6520 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6524 = _T_6522 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6525 = _T_6519 | _T_6524; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6535 = _T_3926 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6536 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6538 = _T_6536 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6540 = _T_6538 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6541 = _T_6535 | _T_6540; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6551 = _T_3930 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6552 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6554 = _T_6552 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6556 = _T_6554 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6557 = _T_6551 | _T_6556; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6567 = _T_3934 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6568 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6570 = _T_6568 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6572 = _T_6570 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6573 = _T_6567 | _T_6572; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6583 = _T_3938 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6584 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6586 = _T_6584 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6588 = _T_6586 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6589 = _T_6583 | _T_6588; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6599 = _T_3942 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6600 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6602 = _T_6600 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6604 = _T_6602 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6605 = _T_6599 | _T_6604; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6615 = _T_3946 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6616 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6618 = _T_6616 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6620 = _T_6618 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6621 = _T_6615 | _T_6620; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6631 = _T_3950 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6632 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6634 = _T_6632 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6636 = _T_6634 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6637 = _T_6631 | _T_6636; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6647 = _T_3954 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6648 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6650 = _T_6648 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6652 = _T_6650 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6653 = _T_6647 | _T_6652; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6663 = _T_3958 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6664 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6666 = _T_6664 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6668 = _T_6666 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6669 = _T_6663 | _T_6668; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6679 = _T_3962 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6680 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6682 = _T_6680 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6684 = _T_6682 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6685 = _T_6679 | _T_6684; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6695 = _T_3966 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6696 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6698 = _T_6696 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6700 = _T_6698 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6701 = _T_6695 | _T_6700; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6711 = _T_3970 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6712 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6714 = _T_6712 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6716 = _T_6714 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6717 = _T_6711 | _T_6716; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6727 = _T_3974 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6728 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6730 = _T_6728 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6732 = _T_6730 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6733 = _T_6727 | _T_6732; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6743 = _T_3978 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6744 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6746 = _T_6744 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6748 = _T_6746 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6749 = _T_6743 | _T_6748; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6759 = _T_3982 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6760 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6762 = _T_6760 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6764 = _T_6762 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6765 = _T_6759 | _T_6764; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6775 = _T_3986 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6776 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6778 = _T_6776 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6780 = _T_6778 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6781 = _T_6775 | _T_6780; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6791 = _T_3990 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6792 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6794 = _T_6792 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6796 = _T_6794 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6797 = _T_6791 | _T_6796; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6807 = _T_3994 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6808 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6810 = _T_6808 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6812 = _T_6810 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6813 = _T_6807 | _T_6812; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6823 = _T_3998 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6824 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6826 = _T_6824 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6828 = _T_6826 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6829 = _T_6823 | _T_6828; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6839 = _T_4002 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6840 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6842 = _T_6840 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6844 = _T_6842 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6845 = _T_6839 | _T_6844; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6855 = _T_4006 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6856 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6858 = _T_6856 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6860 = _T_6858 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6861 = _T_6855 | _T_6860; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6871 = _T_4010 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6872 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6874 = _T_6872 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6876 = _T_6874 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6877 = _T_6871 | _T_6876; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6887 = _T_4014 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6888 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6890 = _T_6888 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6892 = _T_6890 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6893 = _T_6887 | _T_6892; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6903 = _T_4018 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6904 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6906 = _T_6904 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6908 = _T_6906 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6909 = _T_6903 | _T_6908; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6919 = _T_4022 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6920 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_6922 = _T_6920 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6924 = _T_6922 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6925 = _T_6919 | _T_6924; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6935 = _T_3898 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6938 = _T_6424 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6940 = _T_6938 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6941 = _T_6935 | _T_6940; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6951 = _T_3902 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6954 = _T_6440 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6956 = _T_6954 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6957 = _T_6951 | _T_6956; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6967 = _T_3906 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6970 = _T_6456 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6972 = _T_6970 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6973 = _T_6967 | _T_6972; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6983 = _T_3910 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_6986 = _T_6472 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_6988 = _T_6986 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_6989 = _T_6983 | _T_6988; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_6999 = _T_3914 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7002 = _T_6488 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7004 = _T_7002 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7005 = _T_6999 | _T_7004; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7015 = _T_3918 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7018 = _T_6504 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7020 = _T_7018 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7021 = _T_7015 | _T_7020; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7031 = _T_3922 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7034 = _T_6520 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7036 = _T_7034 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7037 = _T_7031 | _T_7036; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7047 = _T_3926 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7050 = _T_6536 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7052 = _T_7050 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7053 = _T_7047 | _T_7052; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7063 = _T_3930 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7066 = _T_6552 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7068 = _T_7066 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7069 = _T_7063 | _T_7068; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7079 = _T_3934 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7082 = _T_6568 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7084 = _T_7082 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7085 = _T_7079 | _T_7084; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7095 = _T_3938 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7098 = _T_6584 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7100 = _T_7098 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7101 = _T_7095 | _T_7100; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7111 = _T_3942 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7114 = _T_6600 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7116 = _T_7114 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7117 = _T_7111 | _T_7116; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7127 = _T_3946 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7130 = _T_6616 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7132 = _T_7130 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7133 = _T_7127 | _T_7132; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7143 = _T_3950 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7146 = _T_6632 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7148 = _T_7146 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7149 = _T_7143 | _T_7148; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7159 = _T_3954 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7162 = _T_6648 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7164 = _T_7162 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7165 = _T_7159 | _T_7164; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7175 = _T_3958 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7178 = _T_6664 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7180 = _T_7178 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7181 = _T_7175 | _T_7180; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7191 = _T_3962 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7194 = _T_6680 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7196 = _T_7194 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7197 = _T_7191 | _T_7196; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7207 = _T_3966 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7210 = _T_6696 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7212 = _T_7210 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7213 = _T_7207 | _T_7212; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7223 = _T_3970 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7226 = _T_6712 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7228 = _T_7226 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7229 = _T_7223 | _T_7228; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7239 = _T_3974 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7242 = _T_6728 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7244 = _T_7242 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7245 = _T_7239 | _T_7244; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7255 = _T_3978 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7258 = _T_6744 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7260 = _T_7258 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7261 = _T_7255 | _T_7260; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7271 = _T_3982 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7274 = _T_6760 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7276 = _T_7274 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7277 = _T_7271 | _T_7276; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7287 = _T_3986 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7290 = _T_6776 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7292 = _T_7290 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7293 = _T_7287 | _T_7292; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7303 = _T_3990 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7306 = _T_6792 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7308 = _T_7306 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7309 = _T_7303 | _T_7308; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7319 = _T_3994 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7322 = _T_6808 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7324 = _T_7322 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7325 = _T_7319 | _T_7324; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7335 = _T_3998 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7338 = _T_6824 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7340 = _T_7338 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7341 = _T_7335 | _T_7340; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7351 = _T_4002 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7354 = _T_6840 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7356 = _T_7354 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7357 = _T_7351 | _T_7356; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7367 = _T_4006 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7370 = _T_6856 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7372 = _T_7370 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7373 = _T_7367 | _T_7372; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7383 = _T_4010 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7386 = _T_6872 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7388 = _T_7386 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7389 = _T_7383 | _T_7388; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7399 = _T_4014 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7402 = _T_6888 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7404 = _T_7402 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7405 = _T_7399 | _T_7404; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7415 = _T_4018 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7418 = _T_6904 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7420 = _T_7418 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7421 = _T_7415 | _T_7420; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7431 = _T_4022 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7434 = _T_6920 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7436 = _T_7434 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7437 = _T_7431 | _T_7436; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7447 = _T_4026 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7448 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7450 = _T_7448 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7452 = _T_7450 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7453 = _T_7447 | _T_7452; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7463 = _T_4030 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7464 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7466 = _T_7464 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7468 = _T_7466 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7469 = _T_7463 | _T_7468; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7479 = _T_4034 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7480 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7482 = _T_7480 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7484 = _T_7482 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7485 = _T_7479 | _T_7484; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7495 = _T_4038 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7496 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7498 = _T_7496 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7500 = _T_7498 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7501 = _T_7495 | _T_7500; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7511 = _T_4042 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7512 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7514 = _T_7512 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7516 = _T_7514 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7517 = _T_7511 | _T_7516; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7527 = _T_4046 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7528 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7530 = _T_7528 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7532 = _T_7530 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7533 = _T_7527 | _T_7532; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7543 = _T_4050 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7544 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7546 = _T_7544 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7548 = _T_7546 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7549 = _T_7543 | _T_7548; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7559 = _T_4054 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7560 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7562 = _T_7560 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7564 = _T_7562 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7565 = _T_7559 | _T_7564; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7575 = _T_4058 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7576 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7578 = _T_7576 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7580 = _T_7578 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7581 = _T_7575 | _T_7580; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7591 = _T_4062 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7592 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7594 = _T_7592 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7596 = _T_7594 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7597 = _T_7591 | _T_7596; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7607 = _T_4066 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7608 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7610 = _T_7608 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7612 = _T_7610 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7613 = _T_7607 | _T_7612; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7623 = _T_4070 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7624 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7626 = _T_7624 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7628 = _T_7626 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7629 = _T_7623 | _T_7628; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7639 = _T_4074 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7640 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7642 = _T_7640 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7644 = _T_7642 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7645 = _T_7639 | _T_7644; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7655 = _T_4078 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7656 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7658 = _T_7656 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7660 = _T_7658 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7661 = _T_7655 | _T_7660; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7671 = _T_4082 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7672 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7674 = _T_7672 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7676 = _T_7674 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7677 = _T_7671 | _T_7676; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7687 = _T_4086 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7688 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7690 = _T_7688 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7692 = _T_7690 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7693 = _T_7687 | _T_7692; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7703 = _T_4090 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7704 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7706 = _T_7704 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7708 = _T_7706 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7709 = _T_7703 | _T_7708; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7719 = _T_4094 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7720 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7722 = _T_7720 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7724 = _T_7722 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7725 = _T_7719 | _T_7724; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7735 = _T_4098 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7736 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7738 = _T_7736 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7740 = _T_7738 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7741 = _T_7735 | _T_7740; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7751 = _T_4102 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7752 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7754 = _T_7752 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7756 = _T_7754 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7757 = _T_7751 | _T_7756; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7767 = _T_4106 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7768 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7770 = _T_7768 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7772 = _T_7770 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7773 = _T_7767 | _T_7772; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7783 = _T_4110 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7784 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7786 = _T_7784 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7788 = _T_7786 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7789 = _T_7783 | _T_7788; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7799 = _T_4114 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7800 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7802 = _T_7800 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7804 = _T_7802 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7805 = _T_7799 | _T_7804; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7815 = _T_4118 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7816 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7818 = _T_7816 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7820 = _T_7818 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7821 = _T_7815 | _T_7820; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7831 = _T_4122 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7832 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7834 = _T_7832 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7836 = _T_7834 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7837 = _T_7831 | _T_7836; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7847 = _T_4126 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7848 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7850 = _T_7848 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7852 = _T_7850 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7853 = _T_7847 | _T_7852; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7863 = _T_4130 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7864 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7866 = _T_7864 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7868 = _T_7866 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7869 = _T_7863 | _T_7868; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7879 = _T_4134 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7880 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7882 = _T_7880 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7884 = _T_7882 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7885 = _T_7879 | _T_7884; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7895 = _T_4138 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7896 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7898 = _T_7896 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7900 = _T_7898 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7901 = _T_7895 | _T_7900; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7911 = _T_4142 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7912 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7914 = _T_7912 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7916 = _T_7914 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7917 = _T_7911 | _T_7916; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7927 = _T_4146 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7928 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7930 = _T_7928 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7932 = _T_7930 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7933 = _T_7927 | _T_7932; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7943 = _T_4150 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7944 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 757:101]
  wire  _T_7946 = _T_7944 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7948 = _T_7946 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7949 = _T_7943 | _T_7948; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7959 = _T_4026 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7962 = _T_7448 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7964 = _T_7962 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7965 = _T_7959 | _T_7964; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7975 = _T_4030 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7978 = _T_7464 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7980 = _T_7978 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7981 = _T_7975 | _T_7980; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_7991 = _T_4034 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_7994 = _T_7480 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_7996 = _T_7994 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_7997 = _T_7991 | _T_7996; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8007 = _T_4038 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8010 = _T_7496 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8012 = _T_8010 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8013 = _T_8007 | _T_8012; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8023 = _T_4042 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8026 = _T_7512 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8028 = _T_8026 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8029 = _T_8023 | _T_8028; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8039 = _T_4046 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8042 = _T_7528 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8044 = _T_8042 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8045 = _T_8039 | _T_8044; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8055 = _T_4050 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8058 = _T_7544 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8060 = _T_8058 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8061 = _T_8055 | _T_8060; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8071 = _T_4054 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8074 = _T_7560 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8076 = _T_8074 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8077 = _T_8071 | _T_8076; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8087 = _T_4058 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8090 = _T_7576 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8092 = _T_8090 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8093 = _T_8087 | _T_8092; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8103 = _T_4062 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8106 = _T_7592 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8108 = _T_8106 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8109 = _T_8103 | _T_8108; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8119 = _T_4066 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8122 = _T_7608 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8124 = _T_8122 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8125 = _T_8119 | _T_8124; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8135 = _T_4070 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8138 = _T_7624 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8140 = _T_8138 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8141 = _T_8135 | _T_8140; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8151 = _T_4074 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8154 = _T_7640 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8156 = _T_8154 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8157 = _T_8151 | _T_8156; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8167 = _T_4078 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8170 = _T_7656 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8172 = _T_8170 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8173 = _T_8167 | _T_8172; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8183 = _T_4082 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8186 = _T_7672 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8188 = _T_8186 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8189 = _T_8183 | _T_8188; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8199 = _T_4086 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8202 = _T_7688 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8204 = _T_8202 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8205 = _T_8199 | _T_8204; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8215 = _T_4090 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8218 = _T_7704 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8220 = _T_8218 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8221 = _T_8215 | _T_8220; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8231 = _T_4094 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8234 = _T_7720 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8236 = _T_8234 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8237 = _T_8231 | _T_8236; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8247 = _T_4098 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8250 = _T_7736 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8252 = _T_8250 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8253 = _T_8247 | _T_8252; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8263 = _T_4102 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8266 = _T_7752 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8268 = _T_8266 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8269 = _T_8263 | _T_8268; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8279 = _T_4106 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8282 = _T_7768 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8284 = _T_8282 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8285 = _T_8279 | _T_8284; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8295 = _T_4110 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8298 = _T_7784 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8300 = _T_8298 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8301 = _T_8295 | _T_8300; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8311 = _T_4114 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8314 = _T_7800 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8316 = _T_8314 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8317 = _T_8311 | _T_8316; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8327 = _T_4118 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8330 = _T_7816 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8332 = _T_8330 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8333 = _T_8327 | _T_8332; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8343 = _T_4122 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8346 = _T_7832 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8348 = _T_8346 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8349 = _T_8343 | _T_8348; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8359 = _T_4126 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8362 = _T_7848 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8364 = _T_8362 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8365 = _T_8359 | _T_8364; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8375 = _T_4130 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8378 = _T_7864 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8380 = _T_8378 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8381 = _T_8375 | _T_8380; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8391 = _T_4134 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8394 = _T_7880 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8396 = _T_8394 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8397 = _T_8391 | _T_8396; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8407 = _T_4138 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8410 = _T_7896 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8412 = _T_8410 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8413 = _T_8407 | _T_8412; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8423 = _T_4142 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8426 = _T_7912 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8428 = _T_8426 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8429 = _T_8423 | _T_8428; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8439 = _T_4146 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8442 = _T_7928 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8444 = _T_8442 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8445 = _T_8439 | _T_8444; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_8455 = _T_4150 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:58]
  wire  _T_8458 = _T_7944 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:123]
  wire  _T_8460 = _T_8458 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:144]
  wire  _T_8461 = _T_8455 | _T_8460; // @[el2_ifu_mem_ctl.scala 757:80]
  wire  _T_9262 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 811:63]
  wire  _T_9263 = _T_9262 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 811:85]
  wire [1:0] _T_9265 = _T_9263 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9272; // @[el2_ifu_mem_ctl.scala 816:57]
  reg  _T_9273; // @[el2_ifu_mem_ctl.scala 817:56]
  reg  _T_9274; // @[el2_ifu_mem_ctl.scala 818:59]
  wire  _T_9275 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 819:80]
  wire  _T_9276 = ifu_bus_arvalid_ff & _T_9275; // @[el2_ifu_mem_ctl.scala 819:78]
  wire  _T_9277 = _T_9276 & miss_pending; // @[el2_ifu_mem_ctl.scala 819:100]
  reg  _T_9278; // @[el2_ifu_mem_ctl.scala 819:58]
  reg  _T_9279; // @[el2_ifu_mem_ctl.scala 820:58]
  wire  _T_9282 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 827:71]
  wire  _T_9284 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 827:124]
  wire  _T_9286 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 828:50]
  wire  _T_9288 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 828:103]
  wire [3:0] _T_9291 = {_T_9282,_T_9284,_T_9286,_T_9288}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 830:53]
  reg  _T_9302; // @[Reg.scala 27:20]
  rvecc_encode_64 m1 ( // @[el2_ifu_mem_ctl.scala 343:18]
    .io_din(m1_io_din),
    .io_ecc_out(m1_io_ecc_out)
  );
  rvecc_encode_64 m2 ( // @[el2_ifu_mem_ctl.scala 344:18]
    .io_din(m2_io_din),
    .io_ecc_out(m2_io_ecc_out)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 329:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 328:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 192:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3097; // @[el2_ifu_mem_ctl.scala 707:21]
  assign io_ifu_pmu_ic_miss = _T_9272; // @[el2_ifu_mem_ctl.scala 816:22]
  assign io_ifu_pmu_ic_hit = _T_9273; // @[el2_ifu_mem_ctl.scala 817:21]
  assign io_ifu_pmu_bus_error = _T_9274; // @[el2_ifu_mem_ctl.scala 818:24]
  assign io_ifu_pmu_bus_busy = _T_9278; // @[el2_ifu_mem_ctl.scala 819:23]
  assign io_ifu_pmu_bus_trxn = _T_9279; // @[el2_ifu_mem_ctl.scala 820:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 143:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 142:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 141:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 152:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 145:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 138:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 136:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 134:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 135:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 144:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 153:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 148:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 569:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_1691; // @[el2_ifu_mem_ctl.scala 570:19]
  assign io_ifu_axi_araddr = _T_1693 & _T_1695; // @[el2_ifu_mem_ctl.scala 571:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 574:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 149:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 572:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 575:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 573:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 151:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 146:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 576:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 666:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 664:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 668:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 659:20]
  assign io_iccm_ready = _T_1794 & _T_1788; // @[el2_ifu_mem_ctl.scala 639:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 338:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 706:15]
  assign io_ic_rd_en = _T_3075 | _T_3080; // @[el2_ifu_mem_ctl.scala 697:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 353:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 353:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 354:23]
  assign io_ifu_ic_debug_rd_data = _T_366; // @[el2_ifu_mem_ctl.scala 362:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 823:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 825:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 826:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 824:25]
  assign io_ic_debug_way = _T_9291[1:0]; // @[el2_ifu_mem_ctl.scala 827:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9265; // @[el2_ifu_mem_ctl.scala 811:19]
  assign io_iccm_rw_addr = _T_2229[14:0]; // @[el2_ifu_mem_ctl.scala 670:19]
  assign io_iccm_wren = _T_1798 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 641:16]
  assign io_iccm_rden = _T_1802 | _T_1803; // @[el2_ifu_mem_ctl.scala 642:16]
  assign io_iccm_wr_data = _T_2204 ? _T_2205 : _T_2212; // @[el2_ifu_mem_ctl.scala 647:19]
  assign io_iccm_wr_size = _T_1808 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 644:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 290:15]
  assign io_ic_access_fault_f = _T_1576 & _T_317; // @[el2_ifu_mem_ctl.scala 395:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_430; // @[el2_ifu_mem_ctl.scala 396:29]
  assign io_iccm_rd_ecc_single_err = _T_3020 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 683:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 684:29]
  assign io_ic_error_start = _T_354 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 356:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 190:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 400:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 392:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 389:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 390:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9302; // @[el2_ifu_mem_ctl.scala 834:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_1581; // @[el2_ifu_mem_ctl.scala 488:27]
  assign io_iccm_correction_state = _T_1609 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 523:28 el2_ifu_mem_ctl.scala 536:32 el2_ifu_mem_ctl.scala 543:32 el2_ifu_mem_ctl.scala 550:32]
  assign io_data = {io_ic_wr_data_1,io_ic_wr_data_0}; // @[el2_ifu_mem_ctl.scala 351:11]
  assign io_ic_wr_ecc = m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 347:16]
  assign m1_io_din = ifu_bus_rdata_ff; // @[el2_ifu_mem_ctl.scala 345:13]
  assign m2_io_din = {_T_1532,_T_1572}; // @[el2_ifu_mem_ctl.scala 349:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4285 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_3641 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_3637 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_3633 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_3629 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_3625 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_3621 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_3617 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_3613 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_3609 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_3605 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_3601 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_3597 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_3593 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_3589 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_3585 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_3581 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_3577 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_3573 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_3569 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_3565 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_3561 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_3557 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_3553 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_3549 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_3545 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_3541 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_3537 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_3533 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_3529 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_3525 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_3521 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_3517 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_3513 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_3509 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_3505 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_3501 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_3497 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_3493 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_3489 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_3485 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_3481 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_3477 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_3473 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_3469 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_3465 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_3461 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_3457 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_3453 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_3449 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_3445 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_3441 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_3437 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_3433 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_3429 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_3425 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_3421 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_3417 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_3413 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_3409 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_3405 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_3401 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_3397 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_3393 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_3389 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_3385 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_3381 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_3377 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_3373 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_3369 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_3365 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_3361 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_3357 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_3353 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_3349 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_3345 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_3341 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_3337 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_3333 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_3329 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_3325 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_3321 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_3317 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_3313 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_3309 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_3305 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_3301 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_3297 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_3293 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_3289 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_3285 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_3281 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_3277 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_3273 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_3269 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_3265 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_3261 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_3257 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_3253 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_3249 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_3245 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_3241 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_3237 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_3233 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_3229 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_3225 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_3221 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_3217 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_3213 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_3209 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_3205 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_3201 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_3197 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_3193 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3189 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3185 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3181 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3177 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3173 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3169 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3165 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3161 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3157 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3153 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3149 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3145 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3141 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3137 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3133 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_366 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_9272 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_9273 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_9274 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_9278 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9279 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9302 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_3641 <= 3'h0;
    end else if (_T_3640) begin
      _T_3641 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3637 <= 3'h0;
    end else if (_T_3636) begin
      _T_3637 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3633 <= 3'h0;
    end else if (_T_3632) begin
      _T_3633 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3629 <= 3'h0;
    end else if (_T_3628) begin
      _T_3629 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3625 <= 3'h0;
    end else if (_T_3624) begin
      _T_3625 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3621 <= 3'h0;
    end else if (_T_3620) begin
      _T_3621 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3617 <= 3'h0;
    end else if (_T_3616) begin
      _T_3617 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3613 <= 3'h0;
    end else if (_T_3612) begin
      _T_3613 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3609 <= 3'h0;
    end else if (_T_3608) begin
      _T_3609 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3605 <= 3'h0;
    end else if (_T_3604) begin
      _T_3605 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3601 <= 3'h0;
    end else if (_T_3600) begin
      _T_3601 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3597 <= 3'h0;
    end else if (_T_3596) begin
      _T_3597 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3593 <= 3'h0;
    end else if (_T_3592) begin
      _T_3593 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3589 <= 3'h0;
    end else if (_T_3588) begin
      _T_3589 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3585 <= 3'h0;
    end else if (_T_3584) begin
      _T_3585 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3581 <= 3'h0;
    end else if (_T_3580) begin
      _T_3581 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3577 <= 3'h0;
    end else if (_T_3576) begin
      _T_3577 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3573 <= 3'h0;
    end else if (_T_3572) begin
      _T_3573 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3569 <= 3'h0;
    end else if (_T_3568) begin
      _T_3569 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3565 <= 3'h0;
    end else if (_T_3564) begin
      _T_3565 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3561 <= 3'h0;
    end else if (_T_3560) begin
      _T_3561 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3557 <= 3'h0;
    end else if (_T_3556) begin
      _T_3557 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3553 <= 3'h0;
    end else if (_T_3552) begin
      _T_3553 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3549 <= 3'h0;
    end else if (_T_3548) begin
      _T_3549 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3545 <= 3'h0;
    end else if (_T_3544) begin
      _T_3545 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3541 <= 3'h0;
    end else if (_T_3540) begin
      _T_3541 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3537 <= 3'h0;
    end else if (_T_3536) begin
      _T_3537 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3533 <= 3'h0;
    end else if (_T_3532) begin
      _T_3533 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3529 <= 3'h0;
    end else if (_T_3528) begin
      _T_3529 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3525 <= 3'h0;
    end else if (_T_3524) begin
      _T_3525 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3521 <= 3'h0;
    end else if (_T_3520) begin
      _T_3521 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3517 <= 3'h0;
    end else if (_T_3516) begin
      _T_3517 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3513 <= 3'h0;
    end else if (_T_3512) begin
      _T_3513 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3509 <= 3'h0;
    end else if (_T_3508) begin
      _T_3509 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3505 <= 3'h0;
    end else if (_T_3504) begin
      _T_3505 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3501 <= 3'h0;
    end else if (_T_3500) begin
      _T_3501 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3497 <= 3'h0;
    end else if (_T_3496) begin
      _T_3497 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3493 <= 3'h0;
    end else if (_T_3492) begin
      _T_3493 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3489 <= 3'h0;
    end else if (_T_3488) begin
      _T_3489 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3485 <= 3'h0;
    end else if (_T_3484) begin
      _T_3485 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3481 <= 3'h0;
    end else if (_T_3480) begin
      _T_3481 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3477 <= 3'h0;
    end else if (_T_3476) begin
      _T_3477 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3473 <= 3'h0;
    end else if (_T_3472) begin
      _T_3473 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3469 <= 3'h0;
    end else if (_T_3468) begin
      _T_3469 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3465 <= 3'h0;
    end else if (_T_3464) begin
      _T_3465 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3461 <= 3'h0;
    end else if (_T_3460) begin
      _T_3461 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3457 <= 3'h0;
    end else if (_T_3456) begin
      _T_3457 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3453 <= 3'h0;
    end else if (_T_3452) begin
      _T_3453 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3449 <= 3'h0;
    end else if (_T_3448) begin
      _T_3449 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3445 <= 3'h0;
    end else if (_T_3444) begin
      _T_3445 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3441 <= 3'h0;
    end else if (_T_3440) begin
      _T_3441 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3437 <= 3'h0;
    end else if (_T_3436) begin
      _T_3437 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3433 <= 3'h0;
    end else if (_T_3432) begin
      _T_3433 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3429 <= 3'h0;
    end else if (_T_3428) begin
      _T_3429 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3425 <= 3'h0;
    end else if (_T_3424) begin
      _T_3425 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3421 <= 3'h0;
    end else if (_T_3420) begin
      _T_3421 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3417 <= 3'h0;
    end else if (_T_3416) begin
      _T_3417 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3413 <= 3'h0;
    end else if (_T_3412) begin
      _T_3413 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3409 <= 3'h0;
    end else if (_T_3408) begin
      _T_3409 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3405 <= 3'h0;
    end else if (_T_3404) begin
      _T_3405 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3401 <= 3'h0;
    end else if (_T_3400) begin
      _T_3401 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3397 <= 3'h0;
    end else if (_T_3396) begin
      _T_3397 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3393 <= 3'h0;
    end else if (_T_3392) begin
      _T_3393 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3389 <= 3'h0;
    end else if (_T_3388) begin
      _T_3389 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3385 <= 3'h0;
    end else if (_T_3384) begin
      _T_3385 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3381 <= 3'h0;
    end else if (_T_3380) begin
      _T_3381 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3377 <= 3'h0;
    end else if (_T_3376) begin
      _T_3377 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3373 <= 3'h0;
    end else if (_T_3372) begin
      _T_3373 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3369 <= 3'h0;
    end else if (_T_3368) begin
      _T_3369 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3365 <= 3'h0;
    end else if (_T_3364) begin
      _T_3365 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3361 <= 3'h0;
    end else if (_T_3360) begin
      _T_3361 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3357 <= 3'h0;
    end else if (_T_3356) begin
      _T_3357 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3353 <= 3'h0;
    end else if (_T_3352) begin
      _T_3353 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3349 <= 3'h0;
    end else if (_T_3348) begin
      _T_3349 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3345 <= 3'h0;
    end else if (_T_3344) begin
      _T_3345 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3341 <= 3'h0;
    end else if (_T_3340) begin
      _T_3341 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3337 <= 3'h0;
    end else if (_T_3336) begin
      _T_3337 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3333 <= 3'h0;
    end else if (_T_3332) begin
      _T_3333 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3329 <= 3'h0;
    end else if (_T_3328) begin
      _T_3329 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3325 <= 3'h0;
    end else if (_T_3324) begin
      _T_3325 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3321 <= 3'h0;
    end else if (_T_3320) begin
      _T_3321 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3317 <= 3'h0;
    end else if (_T_3316) begin
      _T_3317 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3313 <= 3'h0;
    end else if (_T_3312) begin
      _T_3313 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3309 <= 3'h0;
    end else if (_T_3308) begin
      _T_3309 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3305 <= 3'h0;
    end else if (_T_3304) begin
      _T_3305 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3301 <= 3'h0;
    end else if (_T_3300) begin
      _T_3301 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3297 <= 3'h0;
    end else if (_T_3296) begin
      _T_3297 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3293 <= 3'h0;
    end else if (_T_3292) begin
      _T_3293 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3289 <= 3'h0;
    end else if (_T_3288) begin
      _T_3289 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3285 <= 3'h0;
    end else if (_T_3284) begin
      _T_3285 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3281 <= 3'h0;
    end else if (_T_3280) begin
      _T_3281 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3277 <= 3'h0;
    end else if (_T_3276) begin
      _T_3277 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3273 <= 3'h0;
    end else if (_T_3272) begin
      _T_3273 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3269 <= 3'h0;
    end else if (_T_3268) begin
      _T_3269 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3265 <= 3'h0;
    end else if (_T_3264) begin
      _T_3265 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3261 <= 3'h0;
    end else if (_T_3260) begin
      _T_3261 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3257 <= 3'h0;
    end else if (_T_3256) begin
      _T_3257 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3253 <= 3'h0;
    end else if (_T_3252) begin
      _T_3253 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3249 <= 3'h0;
    end else if (_T_3248) begin
      _T_3249 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3245 <= 3'h0;
    end else if (_T_3244) begin
      _T_3245 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3241 <= 3'h0;
    end else if (_T_3240) begin
      _T_3241 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3237 <= 3'h0;
    end else if (_T_3236) begin
      _T_3237 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3233 <= 3'h0;
    end else if (_T_3232) begin
      _T_3233 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3229 <= 3'h0;
    end else if (_T_3228) begin
      _T_3229 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3225 <= 3'h0;
    end else if (_T_3224) begin
      _T_3225 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3221 <= 3'h0;
    end else if (_T_3220) begin
      _T_3221 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3217 <= 3'h0;
    end else if (_T_3216) begin
      _T_3217 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3213 <= 3'h0;
    end else if (_T_3212) begin
      _T_3213 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3209 <= 3'h0;
    end else if (_T_3208) begin
      _T_3209 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3205 <= 3'h0;
    end else if (_T_3204) begin
      _T_3205 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3201 <= 3'h0;
    end else if (_T_3200) begin
      _T_3201 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3197 <= 3'h0;
    end else if (_T_3196) begin
      _T_3197 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3193 <= 3'h0;
    end else if (_T_3192) begin
      _T_3193 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3189 <= 3'h0;
    end else if (_T_3188) begin
      _T_3189 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3185 <= 3'h0;
    end else if (_T_3184) begin
      _T_3185 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3181 <= 3'h0;
    end else if (_T_3180) begin
      _T_3181 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3177 <= 3'h0;
    end else if (_T_3176) begin
      _T_3177 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3173 <= 3'h0;
    end else if (_T_3172) begin
      _T_3173 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3169 <= 3'h0;
    end else if (_T_3168) begin
      _T_3169 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3165 <= 3'h0;
    end else if (_T_3164) begin
      _T_3165 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3161 <= 3'h0;
    end else if (_T_3160) begin
      _T_3161 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3157 <= 3'h0;
    end else if (_T_3156) begin
      _T_3157 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3153 <= 3'h0;
    end else if (_T_3152) begin
      _T_3153 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3149 <= 3'h0;
    end else if (_T_3148) begin
      _T_3149 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3145 <= 3'h0;
    end else if (_T_3144) begin
      _T_3145 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3141 <= 3'h0;
    end else if (_T_3140) begin
      _T_3141 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3137 <= 3'h0;
    end else if (_T_3136) begin
      _T_3137 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3133 <= 3'h0;
    end else if (_T_3132) begin
      _T_3133 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_289;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_1734) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_1730;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_4893) begin
      ic_tag_valid_out_1_0 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_4909) begin
      ic_tag_valid_out_1_1 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_4925) begin
      ic_tag_valid_out_1_2 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_4941) begin
      ic_tag_valid_out_1_3 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_4957) begin
      ic_tag_valid_out_1_4 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_4973) begin
      ic_tag_valid_out_1_5 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_4989) begin
      ic_tag_valid_out_1_6 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5005) begin
      ic_tag_valid_out_1_7 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5021) begin
      ic_tag_valid_out_1_8 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5037) begin
      ic_tag_valid_out_1_9 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5053) begin
      ic_tag_valid_out_1_10 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5069) begin
      ic_tag_valid_out_1_11 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5085) begin
      ic_tag_valid_out_1_12 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5101) begin
      ic_tag_valid_out_1_13 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5117) begin
      ic_tag_valid_out_1_14 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5133) begin
      ic_tag_valid_out_1_15 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5149) begin
      ic_tag_valid_out_1_16 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5165) begin
      ic_tag_valid_out_1_17 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5181) begin
      ic_tag_valid_out_1_18 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5197) begin
      ic_tag_valid_out_1_19 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5213) begin
      ic_tag_valid_out_1_20 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5229) begin
      ic_tag_valid_out_1_21 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5245) begin
      ic_tag_valid_out_1_22 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5261) begin
      ic_tag_valid_out_1_23 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5277) begin
      ic_tag_valid_out_1_24 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5293) begin
      ic_tag_valid_out_1_25 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5309) begin
      ic_tag_valid_out_1_26 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5325) begin
      ic_tag_valid_out_1_27 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_5341) begin
      ic_tag_valid_out_1_28 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_5357) begin
      ic_tag_valid_out_1_29 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_5373) begin
      ic_tag_valid_out_1_30 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_5389) begin
      ic_tag_valid_out_1_31 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_5917) begin
      ic_tag_valid_out_1_32 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_5933) begin
      ic_tag_valid_out_1_33 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_5949) begin
      ic_tag_valid_out_1_34 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_5965) begin
      ic_tag_valid_out_1_35 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_5981) begin
      ic_tag_valid_out_1_36 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_5997) begin
      ic_tag_valid_out_1_37 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6013) begin
      ic_tag_valid_out_1_38 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6029) begin
      ic_tag_valid_out_1_39 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6045) begin
      ic_tag_valid_out_1_40 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6061) begin
      ic_tag_valid_out_1_41 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6077) begin
      ic_tag_valid_out_1_42 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6093) begin
      ic_tag_valid_out_1_43 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6109) begin
      ic_tag_valid_out_1_44 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6125) begin
      ic_tag_valid_out_1_45 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6141) begin
      ic_tag_valid_out_1_46 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6157) begin
      ic_tag_valid_out_1_47 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6173) begin
      ic_tag_valid_out_1_48 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6189) begin
      ic_tag_valid_out_1_49 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6205) begin
      ic_tag_valid_out_1_50 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6221) begin
      ic_tag_valid_out_1_51 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6237) begin
      ic_tag_valid_out_1_52 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6253) begin
      ic_tag_valid_out_1_53 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6269) begin
      ic_tag_valid_out_1_54 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6285) begin
      ic_tag_valid_out_1_55 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6301) begin
      ic_tag_valid_out_1_56 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6317) begin
      ic_tag_valid_out_1_57 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6333) begin
      ic_tag_valid_out_1_58 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6349) begin
      ic_tag_valid_out_1_59 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6365) begin
      ic_tag_valid_out_1_60 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6381) begin
      ic_tag_valid_out_1_61 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_6397) begin
      ic_tag_valid_out_1_62 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_6413) begin
      ic_tag_valid_out_1_63 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_6941) begin
      ic_tag_valid_out_1_64 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_6957) begin
      ic_tag_valid_out_1_65 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_6973) begin
      ic_tag_valid_out_1_66 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_6989) begin
      ic_tag_valid_out_1_67 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7005) begin
      ic_tag_valid_out_1_68 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7021) begin
      ic_tag_valid_out_1_69 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7037) begin
      ic_tag_valid_out_1_70 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7053) begin
      ic_tag_valid_out_1_71 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7069) begin
      ic_tag_valid_out_1_72 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7085) begin
      ic_tag_valid_out_1_73 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7101) begin
      ic_tag_valid_out_1_74 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7117) begin
      ic_tag_valid_out_1_75 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7133) begin
      ic_tag_valid_out_1_76 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7149) begin
      ic_tag_valid_out_1_77 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7165) begin
      ic_tag_valid_out_1_78 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7181) begin
      ic_tag_valid_out_1_79 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7197) begin
      ic_tag_valid_out_1_80 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7213) begin
      ic_tag_valid_out_1_81 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7229) begin
      ic_tag_valid_out_1_82 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7245) begin
      ic_tag_valid_out_1_83 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7261) begin
      ic_tag_valid_out_1_84 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7277) begin
      ic_tag_valid_out_1_85 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7293) begin
      ic_tag_valid_out_1_86 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7309) begin
      ic_tag_valid_out_1_87 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7325) begin
      ic_tag_valid_out_1_88 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7341) begin
      ic_tag_valid_out_1_89 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7357) begin
      ic_tag_valid_out_1_90 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7373) begin
      ic_tag_valid_out_1_91 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7389) begin
      ic_tag_valid_out_1_92 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7405) begin
      ic_tag_valid_out_1_93 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7421) begin
      ic_tag_valid_out_1_94 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7437) begin
      ic_tag_valid_out_1_95 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_7965) begin
      ic_tag_valid_out_1_96 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_7981) begin
      ic_tag_valid_out_1_97 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_7997) begin
      ic_tag_valid_out_1_98 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8013) begin
      ic_tag_valid_out_1_99 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8029) begin
      ic_tag_valid_out_1_100 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8045) begin
      ic_tag_valid_out_1_101 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8061) begin
      ic_tag_valid_out_1_102 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8077) begin
      ic_tag_valid_out_1_103 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8093) begin
      ic_tag_valid_out_1_104 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8109) begin
      ic_tag_valid_out_1_105 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8125) begin
      ic_tag_valid_out_1_106 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8141) begin
      ic_tag_valid_out_1_107 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8157) begin
      ic_tag_valid_out_1_108 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8173) begin
      ic_tag_valid_out_1_109 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8189) begin
      ic_tag_valid_out_1_110 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8205) begin
      ic_tag_valid_out_1_111 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8221) begin
      ic_tag_valid_out_1_112 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8237) begin
      ic_tag_valid_out_1_113 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8253) begin
      ic_tag_valid_out_1_114 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8269) begin
      ic_tag_valid_out_1_115 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8285) begin
      ic_tag_valid_out_1_116 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8301) begin
      ic_tag_valid_out_1_117 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8317) begin
      ic_tag_valid_out_1_118 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8333) begin
      ic_tag_valid_out_1_119 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8349) begin
      ic_tag_valid_out_1_120 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8365) begin
      ic_tag_valid_out_1_121 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8381) begin
      ic_tag_valid_out_1_122 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8397) begin
      ic_tag_valid_out_1_123 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8413) begin
      ic_tag_valid_out_1_124 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8429) begin
      ic_tag_valid_out_1_125 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8445) begin
      ic_tag_valid_out_1_126 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8461) begin
      ic_tag_valid_out_1_127 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_4381) begin
      ic_tag_valid_out_0_0 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_4397) begin
      ic_tag_valid_out_0_1 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_4413) begin
      ic_tag_valid_out_0_2 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_4429) begin
      ic_tag_valid_out_0_3 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_4445) begin
      ic_tag_valid_out_0_4 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_4461) begin
      ic_tag_valid_out_0_5 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_4477) begin
      ic_tag_valid_out_0_6 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_4493) begin
      ic_tag_valid_out_0_7 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_4509) begin
      ic_tag_valid_out_0_8 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_4525) begin
      ic_tag_valid_out_0_9 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_4541) begin
      ic_tag_valid_out_0_10 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_4557) begin
      ic_tag_valid_out_0_11 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_4573) begin
      ic_tag_valid_out_0_12 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_4589) begin
      ic_tag_valid_out_0_13 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_4605) begin
      ic_tag_valid_out_0_14 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_4621) begin
      ic_tag_valid_out_0_15 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_4637) begin
      ic_tag_valid_out_0_16 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_4653) begin
      ic_tag_valid_out_0_17 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_4669) begin
      ic_tag_valid_out_0_18 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_4685) begin
      ic_tag_valid_out_0_19 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_4701) begin
      ic_tag_valid_out_0_20 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_4717) begin
      ic_tag_valid_out_0_21 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_4733) begin
      ic_tag_valid_out_0_22 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_4749) begin
      ic_tag_valid_out_0_23 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_4765) begin
      ic_tag_valid_out_0_24 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_4781) begin
      ic_tag_valid_out_0_25 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_4797) begin
      ic_tag_valid_out_0_26 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_4813) begin
      ic_tag_valid_out_0_27 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_4829) begin
      ic_tag_valid_out_0_28 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_4845) begin
      ic_tag_valid_out_0_29 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_4861) begin
      ic_tag_valid_out_0_30 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_4877) begin
      ic_tag_valid_out_0_31 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_5405) begin
      ic_tag_valid_out_0_32 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_5421) begin
      ic_tag_valid_out_0_33 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_5437) begin
      ic_tag_valid_out_0_34 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_5453) begin
      ic_tag_valid_out_0_35 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_5469) begin
      ic_tag_valid_out_0_36 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_5485) begin
      ic_tag_valid_out_0_37 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_5501) begin
      ic_tag_valid_out_0_38 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_5517) begin
      ic_tag_valid_out_0_39 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_5533) begin
      ic_tag_valid_out_0_40 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_5549) begin
      ic_tag_valid_out_0_41 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_5565) begin
      ic_tag_valid_out_0_42 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_5581) begin
      ic_tag_valid_out_0_43 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_5597) begin
      ic_tag_valid_out_0_44 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_5613) begin
      ic_tag_valid_out_0_45 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_5629) begin
      ic_tag_valid_out_0_46 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_5645) begin
      ic_tag_valid_out_0_47 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_5661) begin
      ic_tag_valid_out_0_48 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_5677) begin
      ic_tag_valid_out_0_49 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_5693) begin
      ic_tag_valid_out_0_50 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_5709) begin
      ic_tag_valid_out_0_51 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_5725) begin
      ic_tag_valid_out_0_52 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_5741) begin
      ic_tag_valid_out_0_53 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_5757) begin
      ic_tag_valid_out_0_54 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_5773) begin
      ic_tag_valid_out_0_55 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_5789) begin
      ic_tag_valid_out_0_56 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_5805) begin
      ic_tag_valid_out_0_57 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_5821) begin
      ic_tag_valid_out_0_58 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_5837) begin
      ic_tag_valid_out_0_59 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_5853) begin
      ic_tag_valid_out_0_60 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_5869) begin
      ic_tag_valid_out_0_61 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_5885) begin
      ic_tag_valid_out_0_62 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_5901) begin
      ic_tag_valid_out_0_63 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_6429) begin
      ic_tag_valid_out_0_64 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_6445) begin
      ic_tag_valid_out_0_65 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_6461) begin
      ic_tag_valid_out_0_66 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_6477) begin
      ic_tag_valid_out_0_67 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_6493) begin
      ic_tag_valid_out_0_68 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_6509) begin
      ic_tag_valid_out_0_69 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_6525) begin
      ic_tag_valid_out_0_70 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_6541) begin
      ic_tag_valid_out_0_71 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_6557) begin
      ic_tag_valid_out_0_72 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_6573) begin
      ic_tag_valid_out_0_73 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_6589) begin
      ic_tag_valid_out_0_74 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_6605) begin
      ic_tag_valid_out_0_75 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_6621) begin
      ic_tag_valid_out_0_76 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_6637) begin
      ic_tag_valid_out_0_77 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_6653) begin
      ic_tag_valid_out_0_78 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_6669) begin
      ic_tag_valid_out_0_79 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_6685) begin
      ic_tag_valid_out_0_80 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_6701) begin
      ic_tag_valid_out_0_81 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_6717) begin
      ic_tag_valid_out_0_82 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_6733) begin
      ic_tag_valid_out_0_83 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_6749) begin
      ic_tag_valid_out_0_84 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_6765) begin
      ic_tag_valid_out_0_85 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_6781) begin
      ic_tag_valid_out_0_86 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_6797) begin
      ic_tag_valid_out_0_87 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_6813) begin
      ic_tag_valid_out_0_88 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_6829) begin
      ic_tag_valid_out_0_89 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_6845) begin
      ic_tag_valid_out_0_90 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_6861) begin
      ic_tag_valid_out_0_91 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_6877) begin
      ic_tag_valid_out_0_92 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_6893) begin
      ic_tag_valid_out_0_93 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_6909) begin
      ic_tag_valid_out_0_94 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_6925) begin
      ic_tag_valid_out_0_95 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7453) begin
      ic_tag_valid_out_0_96 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_7469) begin
      ic_tag_valid_out_0_97 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_7485) begin
      ic_tag_valid_out_0_98 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_7501) begin
      ic_tag_valid_out_0_99 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_7517) begin
      ic_tag_valid_out_0_100 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_7533) begin
      ic_tag_valid_out_0_101 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_7549) begin
      ic_tag_valid_out_0_102 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_7565) begin
      ic_tag_valid_out_0_103 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_7581) begin
      ic_tag_valid_out_0_104 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_7597) begin
      ic_tag_valid_out_0_105 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_7613) begin
      ic_tag_valid_out_0_106 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_7629) begin
      ic_tag_valid_out_0_107 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_7645) begin
      ic_tag_valid_out_0_108 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_7661) begin
      ic_tag_valid_out_0_109 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_7677) begin
      ic_tag_valid_out_0_110 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_7693) begin
      ic_tag_valid_out_0_111 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_7709) begin
      ic_tag_valid_out_0_112 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_7725) begin
      ic_tag_valid_out_0_113 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_7741) begin
      ic_tag_valid_out_0_114 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_7757) begin
      ic_tag_valid_out_0_115 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_7773) begin
      ic_tag_valid_out_0_116 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_7789) begin
      ic_tag_valid_out_0_117 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_7805) begin
      ic_tag_valid_out_0_118 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_7821) begin
      ic_tag_valid_out_0_119 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_7837) begin
      ic_tag_valid_out_0_120 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_7853) begin
      ic_tag_valid_out_0_121 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_7869) begin
      ic_tag_valid_out_0_122 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_7885) begin
      ic_tag_valid_out_0_123 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_7901) begin
      ic_tag_valid_out_0_124 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_7917) begin
      ic_tag_valid_out_0_125 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_7933) begin
      ic_tag_valid_out_0_126 <= _T_4372;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_7949) begin
      ic_tag_valid_out_0_127 <= _T_4372;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_366 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_366 <= {{5'd0}, _T_365};
    end else begin
      _T_366 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_1683) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_1758) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_1802;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_1584) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_1586) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_1596) begin
        perr_state <= 3'h0;
      end else if (_T_1599) begin
        if (_T_1601) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_1605) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_1609) begin
        err_stop_state <= 2'h1;
      end else if (_T_1614) begin
        if (_T_1616) begin
          err_stop_state <= 2'h0;
        end else if (_T_1637) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_1641) begin
        if (_T_1616) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_1658) begin
        if (_T_1662) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_527;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_4285 <= 7'h0;
    end else if (_T_3106) begin
      _T_4285 <= io_ic_debug_addr[9:3];
    end else begin
      _T_4285 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_567;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3041;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_2216;
    end else begin
      iccm_dma_rdata <= _T_2217;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3037;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3106) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3109) begin
      way_status_new_ff <= _T_3113;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3109) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_9302 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9302 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_9272 <= 1'h0;
    end else begin
      _T_9272 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_9273 <= 1'h0;
    end else begin
      _T_9273 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_9274 <= 1'h0;
    end else begin
      _T_9274 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_9278 <= 1'h0;
    end else begin
      _T_9278 <= _T_9277;
    end
    if (reset) begin
      _T_9279 <= 1'h0;
    end else begin
      _T_9279 <= bus_cmd_sent;
    end
  end
endmodule
