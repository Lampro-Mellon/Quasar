module rvclkhdr(
  input   io_clk,
  input   io_en
);
  wire  clkhdr_Q; // @[lib.scala 334:26]
  wire  clkhdr_CK; // @[lib.scala 334:26]
  wire  clkhdr_EN; // @[lib.scala 334:26]
  wire  clkhdr_SE; // @[lib.scala 334:26]
  gated_latch clkhdr ( // @[lib.scala 334:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign clkhdr_CK = io_clk; // @[lib.scala 336:18]
  assign clkhdr_EN = io_en; // @[lib.scala 337:18]
  assign clkhdr_SE = 1'h0; // @[lib.scala 338:18]
endmodule
module ifu_bp_ctl(
  input         clock,
  input         reset,
  input         io_active_clk,
  input         io_ic_hit_f,
  input         io_exu_flush_final,
  input  [30:0] io_ifc_fetch_addr_f,
  input         io_ifc_fetch_req_f,
  input         io_dec_bp_dec_tlu_br0_r_pkt_valid,
  input  [1:0]  io_dec_bp_dec_tlu_br0_r_pkt_bits_hist,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_way,
  input         io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,
  input         io_dec_bp_dec_tlu_flush_leak_one_wb,
  input         io_dec_bp_dec_tlu_bpred_disable,
  input         io_dec_tlu_flush_lower_wb,
  input  [7:0]  io_exu_bp_exu_i0_br_index_r,
  input  [7:0]  io_exu_bp_exu_i0_br_fghr_r,
  input         io_exu_bp_exu_i0_br_way_r,
  input         io_exu_bp_exu_mp_pkt_valid,
  input         io_exu_bp_exu_mp_pkt_bits_misp,
  input         io_exu_bp_exu_mp_pkt_bits_ataken,
  input         io_exu_bp_exu_mp_pkt_bits_boffset,
  input         io_exu_bp_exu_mp_pkt_bits_pc4,
  input  [1:0]  io_exu_bp_exu_mp_pkt_bits_hist,
  input  [11:0] io_exu_bp_exu_mp_pkt_bits_toffset,
  input         io_exu_bp_exu_mp_pkt_bits_br_error,
  input         io_exu_bp_exu_mp_pkt_bits_br_start_error,
  input         io_exu_bp_exu_mp_pkt_bits_pcall,
  input         io_exu_bp_exu_mp_pkt_bits_pja,
  input         io_exu_bp_exu_mp_pkt_bits_way,
  input         io_exu_bp_exu_mp_pkt_bits_pret,
  input  [30:0] io_exu_bp_exu_mp_pkt_bits_prett,
  input  [7:0]  io_exu_bp_exu_mp_eghr,
  input  [7:0]  io_exu_bp_exu_mp_fghr,
  input  [7:0]  io_exu_bp_exu_mp_index,
  input  [4:0]  io_exu_bp_exu_mp_btag,
  input  [8:0]  io_dec_fa_error_index,
  output        io_ifu_bp_hit_taken_f,
  output [30:0] io_ifu_bp_btb_target_f,
  output        io_ifu_bp_inst_mask_f,
  output [7:0]  io_ifu_bp_fghr_f,
  output [1:0]  io_ifu_bp_way_f,
  output [1:0]  io_ifu_bp_ret_f,
  output [1:0]  io_ifu_bp_hist1_f,
  output [1:0]  io_ifu_bp_hist0_f,
  output [1:0]  io_ifu_bp_pc4_f,
  output [1:0]  io_ifu_bp_valid_f,
  output [11:0] io_ifu_bp_poffset_f,
  output [8:0]  io_ifu_bp_fa_index_f_0,
  output [8:0]  io_ifu_bp_fa_index_f_1,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_638;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
  reg [31:0] _RAND_901;
  reg [31:0] _RAND_902;
  reg [31:0] _RAND_903;
  reg [31:0] _RAND_904;
  reg [31:0] _RAND_905;
  reg [31:0] _RAND_906;
  reg [31:0] _RAND_907;
  reg [31:0] _RAND_908;
  reg [31:0] _RAND_909;
  reg [31:0] _RAND_910;
  reg [31:0] _RAND_911;
  reg [31:0] _RAND_912;
  reg [31:0] _RAND_913;
  reg [31:0] _RAND_914;
  reg [31:0] _RAND_915;
  reg [31:0] _RAND_916;
  reg [31:0] _RAND_917;
  reg [31:0] _RAND_918;
  reg [31:0] _RAND_919;
  reg [31:0] _RAND_920;
  reg [31:0] _RAND_921;
  reg [31:0] _RAND_922;
  reg [31:0] _RAND_923;
  reg [31:0] _RAND_924;
  reg [31:0] _RAND_925;
  reg [31:0] _RAND_926;
  reg [31:0] _RAND_927;
  reg [31:0] _RAND_928;
  reg [31:0] _RAND_929;
  reg [31:0] _RAND_930;
  reg [31:0] _RAND_931;
  reg [31:0] _RAND_932;
  reg [31:0] _RAND_933;
  reg [31:0] _RAND_934;
  reg [31:0] _RAND_935;
  reg [31:0] _RAND_936;
  reg [31:0] _RAND_937;
  reg [31:0] _RAND_938;
  reg [31:0] _RAND_939;
  reg [31:0] _RAND_940;
  reg [31:0] _RAND_941;
  reg [31:0] _RAND_942;
  reg [31:0] _RAND_943;
  reg [31:0] _RAND_944;
  reg [31:0] _RAND_945;
  reg [31:0] _RAND_946;
  reg [31:0] _RAND_947;
  reg [31:0] _RAND_948;
  reg [31:0] _RAND_949;
  reg [31:0] _RAND_950;
  reg [31:0] _RAND_951;
  reg [31:0] _RAND_952;
  reg [31:0] _RAND_953;
  reg [31:0] _RAND_954;
  reg [31:0] _RAND_955;
  reg [31:0] _RAND_956;
  reg [31:0] _RAND_957;
  reg [31:0] _RAND_958;
  reg [31:0] _RAND_959;
  reg [31:0] _RAND_960;
  reg [31:0] _RAND_961;
  reg [31:0] _RAND_962;
  reg [31:0] _RAND_963;
  reg [31:0] _RAND_964;
  reg [31:0] _RAND_965;
  reg [31:0] _RAND_966;
  reg [31:0] _RAND_967;
  reg [31:0] _RAND_968;
  reg [31:0] _RAND_969;
  reg [31:0] _RAND_970;
  reg [31:0] _RAND_971;
  reg [31:0] _RAND_972;
  reg [31:0] _RAND_973;
  reg [31:0] _RAND_974;
  reg [31:0] _RAND_975;
  reg [31:0] _RAND_976;
  reg [31:0] _RAND_977;
  reg [31:0] _RAND_978;
  reg [31:0] _RAND_979;
  reg [31:0] _RAND_980;
  reg [31:0] _RAND_981;
  reg [31:0] _RAND_982;
  reg [31:0] _RAND_983;
  reg [31:0] _RAND_984;
  reg [31:0] _RAND_985;
  reg [31:0] _RAND_986;
  reg [31:0] _RAND_987;
  reg [31:0] _RAND_988;
  reg [31:0] _RAND_989;
  reg [31:0] _RAND_990;
  reg [31:0] _RAND_991;
  reg [31:0] _RAND_992;
  reg [31:0] _RAND_993;
  reg [31:0] _RAND_994;
  reg [31:0] _RAND_995;
  reg [31:0] _RAND_996;
  reg [31:0] _RAND_997;
  reg [31:0] _RAND_998;
  reg [31:0] _RAND_999;
  reg [31:0] _RAND_1000;
  reg [31:0] _RAND_1001;
  reg [31:0] _RAND_1002;
  reg [31:0] _RAND_1003;
  reg [31:0] _RAND_1004;
  reg [31:0] _RAND_1005;
  reg [31:0] _RAND_1006;
  reg [31:0] _RAND_1007;
  reg [31:0] _RAND_1008;
  reg [31:0] _RAND_1009;
  reg [31:0] _RAND_1010;
  reg [31:0] _RAND_1011;
  reg [31:0] _RAND_1012;
  reg [31:0] _RAND_1013;
  reg [31:0] _RAND_1014;
  reg [31:0] _RAND_1015;
  reg [31:0] _RAND_1016;
  reg [31:0] _RAND_1017;
  reg [31:0] _RAND_1018;
  reg [31:0] _RAND_1019;
  reg [31:0] _RAND_1020;
  reg [31:0] _RAND_1021;
  reg [31:0] _RAND_1022;
  reg [31:0] _RAND_1023;
  reg [31:0] _RAND_1024;
  reg [31:0] _RAND_1025;
  reg [31:0] _RAND_1026;
  reg [255:0] _RAND_1027;
  reg [31:0] _RAND_1028;
  reg [31:0] _RAND_1029;
  reg [31:0] _RAND_1030;
  reg [31:0] _RAND_1031;
  reg [31:0] _RAND_1032;
  reg [31:0] _RAND_1033;
  reg [31:0] _RAND_1034;
  reg [31:0] _RAND_1035;
  reg [31:0] _RAND_1036;
  reg [31:0] _RAND_1037;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_1_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_2_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_3_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_4_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_5_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_6_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_7_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_8_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_9_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_10_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_11_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_12_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_13_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_14_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_15_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_16_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_17_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_18_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_19_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_20_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_21_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_22_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_23_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_23_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_24_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_24_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_25_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_25_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_26_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_26_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_27_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_27_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_28_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_28_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_29_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_29_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_30_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_30_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_31_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_31_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_32_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_32_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_33_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_33_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_34_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_34_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_35_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_35_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_36_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_36_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_37_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_37_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_38_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_38_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_39_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_39_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_40_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_40_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_41_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_41_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_42_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_42_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_43_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_43_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_44_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_44_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_45_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_45_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_46_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_46_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_47_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_47_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_48_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_48_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_49_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_49_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_50_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_50_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_51_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_51_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_52_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_52_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_53_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_53_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_54_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_54_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_55_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_55_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_56_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_56_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_57_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_57_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_58_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_58_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_59_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_59_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_60_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_60_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_61_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_61_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_62_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_62_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_63_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_63_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_64_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_64_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_65_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_65_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_66_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_66_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_67_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_67_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_68_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_68_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_69_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_69_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_70_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_70_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_71_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_71_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_72_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_72_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_73_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_73_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_74_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_74_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_75_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_75_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_76_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_76_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_77_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_77_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_78_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_78_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_79_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_79_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_80_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_80_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_81_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_81_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_82_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_82_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_83_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_83_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_84_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_84_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_85_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_85_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_86_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_86_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_87_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_87_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_88_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_88_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_89_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_89_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_90_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_90_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_91_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_91_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_92_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_92_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_93_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_93_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_94_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_94_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_95_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_95_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_96_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_96_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_97_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_97_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_98_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_98_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_99_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_99_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_100_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_100_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_101_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_101_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_102_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_102_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_103_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_103_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_104_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_104_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_105_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_105_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_106_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_106_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_107_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_107_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_108_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_108_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_109_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_109_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_110_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_110_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_111_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_111_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_112_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_112_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_113_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_113_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_114_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_114_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_115_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_115_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_116_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_116_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_117_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_117_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_118_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_118_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_119_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_119_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_120_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_120_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_121_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_121_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_122_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_122_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_123_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_123_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_124_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_124_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_125_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_125_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_126_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_126_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_127_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_127_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_128_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_128_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_129_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_129_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_130_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_130_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_131_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_131_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_132_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_132_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_133_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_133_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_134_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_134_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_135_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_135_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_136_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_136_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_137_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_137_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_138_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_138_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_139_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_139_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_140_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_140_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_141_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_141_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_142_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_142_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_143_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_143_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_144_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_144_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_145_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_145_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_146_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_146_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_147_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_147_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_148_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_148_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_149_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_149_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_150_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_150_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_151_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_151_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_152_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_152_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_153_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_153_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_154_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_154_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_155_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_155_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_156_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_156_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_157_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_157_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_158_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_158_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_159_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_159_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_160_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_160_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_161_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_161_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_162_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_162_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_163_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_163_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_164_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_164_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_165_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_165_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_166_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_166_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_167_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_167_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_168_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_168_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_169_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_169_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_170_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_170_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_171_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_171_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_172_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_172_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_173_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_173_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_174_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_174_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_175_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_175_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_176_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_176_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_177_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_177_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_178_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_178_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_179_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_179_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_180_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_180_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_181_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_181_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_182_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_182_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_183_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_183_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_184_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_184_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_185_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_185_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_186_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_186_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_187_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_187_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_188_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_188_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_189_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_189_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_190_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_190_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_191_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_191_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_192_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_192_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_193_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_193_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_194_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_194_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_195_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_195_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_196_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_196_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_197_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_197_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_198_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_198_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_199_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_199_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_200_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_200_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_201_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_201_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_202_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_202_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_203_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_203_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_204_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_204_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_205_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_205_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_206_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_206_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_207_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_207_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_208_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_208_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_209_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_209_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_210_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_210_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_211_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_211_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_212_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_212_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_213_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_213_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_214_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_214_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_215_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_215_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_216_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_216_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_217_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_217_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_218_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_218_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_219_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_219_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_220_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_220_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_221_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_221_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_222_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_222_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_223_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_223_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_224_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_224_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_225_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_225_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_226_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_226_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_227_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_227_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_228_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_228_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_229_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_229_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_230_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_230_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_231_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_231_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_232_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_232_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_233_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_233_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_234_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_234_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_235_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_235_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_236_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_236_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_237_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_237_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_238_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_238_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_239_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_239_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_240_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_240_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_241_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_241_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_242_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_242_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_243_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_243_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_244_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_244_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_245_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_245_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_246_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_246_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_247_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_247_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_248_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_248_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_249_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_249_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_250_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_250_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_251_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_251_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_252_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_252_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_253_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_253_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_254_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_254_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_255_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_255_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_256_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_256_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_257_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_257_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_258_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_258_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_259_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_259_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_260_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_260_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_261_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_261_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_262_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_262_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_263_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_263_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_264_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_264_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_265_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_265_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_266_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_266_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_267_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_267_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_268_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_268_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_269_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_269_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_270_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_270_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_271_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_271_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_272_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_272_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_273_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_273_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_274_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_274_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_275_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_275_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_276_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_276_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_277_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_277_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_278_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_278_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_279_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_279_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_280_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_280_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_281_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_281_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_282_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_282_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_283_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_283_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_284_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_284_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_285_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_285_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_286_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_286_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_287_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_287_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_288_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_288_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_289_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_289_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_290_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_290_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_291_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_291_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_292_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_292_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_293_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_293_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_294_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_294_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_295_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_295_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_296_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_296_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_297_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_297_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_298_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_298_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_299_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_299_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_300_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_300_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_301_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_301_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_302_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_302_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_303_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_303_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_304_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_304_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_305_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_305_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_306_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_306_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_307_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_307_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_308_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_308_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_309_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_309_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_310_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_310_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_311_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_311_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_312_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_312_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_313_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_313_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_314_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_314_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_315_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_315_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_316_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_316_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_317_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_317_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_318_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_318_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_319_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_319_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_320_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_320_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_321_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_321_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_322_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_322_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_323_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_323_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_324_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_324_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_325_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_325_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_326_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_326_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_327_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_327_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_328_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_328_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_329_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_329_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_330_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_330_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_331_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_331_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_332_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_332_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_333_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_333_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_334_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_334_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_335_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_335_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_336_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_336_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_337_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_337_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_338_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_338_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_339_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_339_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_340_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_340_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_341_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_341_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_342_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_342_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_343_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_343_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_344_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_344_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_345_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_345_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_346_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_346_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_347_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_347_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_348_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_348_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_349_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_349_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_350_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_350_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_351_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_351_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_352_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_352_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_353_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_353_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_354_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_354_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_355_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_355_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_356_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_356_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_357_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_357_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_358_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_358_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_359_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_359_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_360_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_360_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_361_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_361_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_362_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_362_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_363_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_363_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_364_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_364_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_365_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_365_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_366_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_366_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_367_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_367_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_368_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_368_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_369_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_369_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_370_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_370_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_371_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_371_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_372_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_372_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_373_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_373_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_374_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_374_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_375_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_375_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_376_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_376_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_377_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_377_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_378_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_378_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_379_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_379_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_380_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_380_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_381_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_381_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_382_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_382_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_383_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_383_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_384_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_384_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_385_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_385_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_386_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_386_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_387_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_387_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_388_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_388_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_389_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_389_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_390_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_390_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_391_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_391_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_392_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_392_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_393_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_393_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_394_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_394_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_395_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_395_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_396_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_396_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_397_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_397_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_398_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_398_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_399_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_399_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_400_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_400_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_401_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_401_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_402_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_402_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_403_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_403_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_404_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_404_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_405_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_405_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_406_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_406_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_407_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_407_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_408_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_408_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_409_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_409_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_410_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_410_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_411_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_411_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_412_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_412_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_413_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_413_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_414_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_414_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_415_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_415_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_416_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_416_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_417_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_417_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_418_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_418_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_419_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_419_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_420_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_420_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_421_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_421_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_422_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_422_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_423_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_423_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_424_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_424_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_425_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_425_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_426_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_426_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_427_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_427_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_428_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_428_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_429_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_429_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_430_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_430_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_431_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_431_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_432_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_432_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_433_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_433_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_434_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_434_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_435_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_435_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_436_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_436_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_437_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_437_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_438_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_438_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_439_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_439_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_440_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_440_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_441_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_441_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_442_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_442_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_443_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_443_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_444_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_444_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_445_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_445_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_446_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_446_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_447_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_447_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_448_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_448_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_449_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_449_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_450_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_450_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_451_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_451_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_452_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_452_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_453_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_453_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_454_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_454_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_455_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_455_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_456_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_456_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_457_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_457_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_458_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_458_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_459_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_459_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_460_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_460_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_461_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_461_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_462_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_462_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_463_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_463_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_464_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_464_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_465_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_465_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_466_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_466_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_467_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_467_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_468_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_468_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_469_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_469_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_470_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_470_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_471_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_471_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_472_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_472_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_473_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_473_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_474_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_474_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_475_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_475_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_476_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_476_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_477_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_477_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_478_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_478_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_479_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_479_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_480_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_480_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_481_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_481_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_482_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_482_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_483_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_483_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_484_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_484_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_485_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_485_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_486_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_486_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_487_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_487_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_488_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_488_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_489_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_489_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_490_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_490_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_491_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_491_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_492_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_492_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_493_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_493_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_494_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_494_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_495_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_495_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_496_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_496_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_497_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_497_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_498_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_498_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_499_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_499_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_500_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_500_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_501_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_501_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_502_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_502_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_503_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_503_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_504_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_504_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_505_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_505_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_506_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_506_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_507_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_507_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_508_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_508_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_509_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_509_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_510_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_510_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_511_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_511_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_512_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_512_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_513_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_513_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_514_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_514_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_515_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_515_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_516_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_516_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_517_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_517_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_518_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_518_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_519_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_519_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_520_io_clk; // @[lib.scala 409:23]
  wire  rvclkhdr_520_io_en; // @[lib.scala 409:23]
  wire  rvclkhdr_521_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_521_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_522_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_523_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_524_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_525_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_526_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_527_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_528_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_529_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_530_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_531_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_532_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_533_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_534_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_535_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_536_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_537_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_538_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_539_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_540_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_541_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_542_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_543_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_544_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_545_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_546_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_547_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_548_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_549_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_550_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_551_io_en; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_clk; // @[lib.scala 343:22]
  wire  rvclkhdr_552_io_en; // @[lib.scala 343:22]
  wire  _T_21 = io_dec_bp_dec_tlu_flush_leak_one_wb & io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 135:54]
  reg  leak_one_f_d1; // @[Reg.scala 27:20]
  wire  _T_22 = ~io_dec_tlu_flush_lower_wb; // @[ifu_bp_ctl.scala 135:102]
  wire  _T_23 = leak_one_f_d1 & _T_22; // @[ifu_bp_ctl.scala 135:100]
  wire  leak_one_f = _T_21 | _T_23; // @[ifu_bp_ctl.scala 135:83]
  wire  _T = ~leak_one_f; // @[ifu_bp_ctl.scala 82:58]
  wire  exu_mp_valid = io_exu_bp_exu_mp_pkt_bits_misp & _T; // @[ifu_bp_ctl.scala 82:56]
  wire  dec_tlu_error_wb = io_dec_bp_dec_tlu_br0_r_pkt_bits_br_start_error | io_dec_bp_dec_tlu_br0_r_pkt_bits_br_error; // @[ifu_bp_ctl.scala 105:50]
  wire [7:0] _T_4 = io_ifc_fetch_addr_f[8:1] ^ io_ifc_fetch_addr_f[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_f = _T_4 ^ io_ifc_fetch_addr_f[24:17]; // @[lib.scala 51:85]
  wire [29:0] fetch_addr_p1_f = io_ifc_fetch_addr_f[30:1] + 30'h1; // @[ifu_bp_ctl.scala 113:51]
  wire [30:0] _T_8 = {fetch_addr_p1_f,1'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_11 = _T_8[8:1] ^ _T_8[16:9]; // @[lib.scala 51:47]
  wire [7:0] btb_rd_addr_p1_f = _T_11 ^ _T_8[24:17]; // @[lib.scala 51:85]
  wire  _T_147 = ~io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 191:37]
  wire  _T_2661 = btb_rd_addr_f == 8'h0; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_3173 = _T_2661 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_2663 = btb_rd_addr_f == 8'h1; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_3174 = _T_2663 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3429 = _T_3173 | _T_3174; // @[Mux.scala 27:72]
  wire  _T_2665 = btb_rd_addr_f == 8'h2; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_3175 = _T_2665 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3430 = _T_3429 | _T_3175; // @[Mux.scala 27:72]
  wire  _T_2667 = btb_rd_addr_f == 8'h3; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_3176 = _T_2667 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3431 = _T_3430 | _T_3176; // @[Mux.scala 27:72]
  wire  _T_2669 = btb_rd_addr_f == 8'h4; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_3177 = _T_2669 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3432 = _T_3431 | _T_3177; // @[Mux.scala 27:72]
  wire  _T_2671 = btb_rd_addr_f == 8'h5; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_3178 = _T_2671 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3433 = _T_3432 | _T_3178; // @[Mux.scala 27:72]
  wire  _T_2673 = btb_rd_addr_f == 8'h6; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_3179 = _T_2673 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3434 = _T_3433 | _T_3179; // @[Mux.scala 27:72]
  wire  _T_2675 = btb_rd_addr_f == 8'h7; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_3180 = _T_2675 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3435 = _T_3434 | _T_3180; // @[Mux.scala 27:72]
  wire  _T_2677 = btb_rd_addr_f == 8'h8; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_3181 = _T_2677 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3436 = _T_3435 | _T_3181; // @[Mux.scala 27:72]
  wire  _T_2679 = btb_rd_addr_f == 8'h9; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_3182 = _T_2679 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3437 = _T_3436 | _T_3182; // @[Mux.scala 27:72]
  wire  _T_2681 = btb_rd_addr_f == 8'ha; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_3183 = _T_2681 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3438 = _T_3437 | _T_3183; // @[Mux.scala 27:72]
  wire  _T_2683 = btb_rd_addr_f == 8'hb; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_3184 = _T_2683 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3439 = _T_3438 | _T_3184; // @[Mux.scala 27:72]
  wire  _T_2685 = btb_rd_addr_f == 8'hc; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_3185 = _T_2685 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3440 = _T_3439 | _T_3185; // @[Mux.scala 27:72]
  wire  _T_2687 = btb_rd_addr_f == 8'hd; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_3186 = _T_2687 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3441 = _T_3440 | _T_3186; // @[Mux.scala 27:72]
  wire  _T_2689 = btb_rd_addr_f == 8'he; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_3187 = _T_2689 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3442 = _T_3441 | _T_3187; // @[Mux.scala 27:72]
  wire  _T_2691 = btb_rd_addr_f == 8'hf; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_3188 = _T_2691 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3443 = _T_3442 | _T_3188; // @[Mux.scala 27:72]
  wire  _T_2693 = btb_rd_addr_f == 8'h10; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_3189 = _T_2693 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3444 = _T_3443 | _T_3189; // @[Mux.scala 27:72]
  wire  _T_2695 = btb_rd_addr_f == 8'h11; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_3190 = _T_2695 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3445 = _T_3444 | _T_3190; // @[Mux.scala 27:72]
  wire  _T_2697 = btb_rd_addr_f == 8'h12; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_3191 = _T_2697 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3446 = _T_3445 | _T_3191; // @[Mux.scala 27:72]
  wire  _T_2699 = btb_rd_addr_f == 8'h13; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_3192 = _T_2699 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3447 = _T_3446 | _T_3192; // @[Mux.scala 27:72]
  wire  _T_2701 = btb_rd_addr_f == 8'h14; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_3193 = _T_2701 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3448 = _T_3447 | _T_3193; // @[Mux.scala 27:72]
  wire  _T_2703 = btb_rd_addr_f == 8'h15; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_3194 = _T_2703 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3449 = _T_3448 | _T_3194; // @[Mux.scala 27:72]
  wire  _T_2705 = btb_rd_addr_f == 8'h16; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_3195 = _T_2705 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3450 = _T_3449 | _T_3195; // @[Mux.scala 27:72]
  wire  _T_2707 = btb_rd_addr_f == 8'h17; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_3196 = _T_2707 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3451 = _T_3450 | _T_3196; // @[Mux.scala 27:72]
  wire  _T_2709 = btb_rd_addr_f == 8'h18; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_3197 = _T_2709 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3452 = _T_3451 | _T_3197; // @[Mux.scala 27:72]
  wire  _T_2711 = btb_rd_addr_f == 8'h19; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_3198 = _T_2711 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3453 = _T_3452 | _T_3198; // @[Mux.scala 27:72]
  wire  _T_2713 = btb_rd_addr_f == 8'h1a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_3199 = _T_2713 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3454 = _T_3453 | _T_3199; // @[Mux.scala 27:72]
  wire  _T_2715 = btb_rd_addr_f == 8'h1b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_3200 = _T_2715 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3455 = _T_3454 | _T_3200; // @[Mux.scala 27:72]
  wire  _T_2717 = btb_rd_addr_f == 8'h1c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_3201 = _T_2717 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3456 = _T_3455 | _T_3201; // @[Mux.scala 27:72]
  wire  _T_2719 = btb_rd_addr_f == 8'h1d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_3202 = _T_2719 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3457 = _T_3456 | _T_3202; // @[Mux.scala 27:72]
  wire  _T_2721 = btb_rd_addr_f == 8'h1e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_3203 = _T_2721 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3458 = _T_3457 | _T_3203; // @[Mux.scala 27:72]
  wire  _T_2723 = btb_rd_addr_f == 8'h1f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_3204 = _T_2723 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3459 = _T_3458 | _T_3204; // @[Mux.scala 27:72]
  wire  _T_2725 = btb_rd_addr_f == 8'h20; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_3205 = _T_2725 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3460 = _T_3459 | _T_3205; // @[Mux.scala 27:72]
  wire  _T_2727 = btb_rd_addr_f == 8'h21; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_3206 = _T_2727 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3461 = _T_3460 | _T_3206; // @[Mux.scala 27:72]
  wire  _T_2729 = btb_rd_addr_f == 8'h22; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_3207 = _T_2729 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3462 = _T_3461 | _T_3207; // @[Mux.scala 27:72]
  wire  _T_2731 = btb_rd_addr_f == 8'h23; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_3208 = _T_2731 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3463 = _T_3462 | _T_3208; // @[Mux.scala 27:72]
  wire  _T_2733 = btb_rd_addr_f == 8'h24; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_3209 = _T_2733 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3464 = _T_3463 | _T_3209; // @[Mux.scala 27:72]
  wire  _T_2735 = btb_rd_addr_f == 8'h25; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_3210 = _T_2735 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3465 = _T_3464 | _T_3210; // @[Mux.scala 27:72]
  wire  _T_2737 = btb_rd_addr_f == 8'h26; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_3211 = _T_2737 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3466 = _T_3465 | _T_3211; // @[Mux.scala 27:72]
  wire  _T_2739 = btb_rd_addr_f == 8'h27; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_3212 = _T_2739 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3467 = _T_3466 | _T_3212; // @[Mux.scala 27:72]
  wire  _T_2741 = btb_rd_addr_f == 8'h28; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_3213 = _T_2741 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3468 = _T_3467 | _T_3213; // @[Mux.scala 27:72]
  wire  _T_2743 = btb_rd_addr_f == 8'h29; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_3214 = _T_2743 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3469 = _T_3468 | _T_3214; // @[Mux.scala 27:72]
  wire  _T_2745 = btb_rd_addr_f == 8'h2a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_3215 = _T_2745 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3470 = _T_3469 | _T_3215; // @[Mux.scala 27:72]
  wire  _T_2747 = btb_rd_addr_f == 8'h2b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_3216 = _T_2747 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3471 = _T_3470 | _T_3216; // @[Mux.scala 27:72]
  wire  _T_2749 = btb_rd_addr_f == 8'h2c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_3217 = _T_2749 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3472 = _T_3471 | _T_3217; // @[Mux.scala 27:72]
  wire  _T_2751 = btb_rd_addr_f == 8'h2d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_3218 = _T_2751 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3473 = _T_3472 | _T_3218; // @[Mux.scala 27:72]
  wire  _T_2753 = btb_rd_addr_f == 8'h2e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_3219 = _T_2753 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3474 = _T_3473 | _T_3219; // @[Mux.scala 27:72]
  wire  _T_2755 = btb_rd_addr_f == 8'h2f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_3220 = _T_2755 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3475 = _T_3474 | _T_3220; // @[Mux.scala 27:72]
  wire  _T_2757 = btb_rd_addr_f == 8'h30; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_3221 = _T_2757 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3476 = _T_3475 | _T_3221; // @[Mux.scala 27:72]
  wire  _T_2759 = btb_rd_addr_f == 8'h31; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_3222 = _T_2759 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3477 = _T_3476 | _T_3222; // @[Mux.scala 27:72]
  wire  _T_2761 = btb_rd_addr_f == 8'h32; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_3223 = _T_2761 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3478 = _T_3477 | _T_3223; // @[Mux.scala 27:72]
  wire  _T_2763 = btb_rd_addr_f == 8'h33; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_3224 = _T_2763 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3479 = _T_3478 | _T_3224; // @[Mux.scala 27:72]
  wire  _T_2765 = btb_rd_addr_f == 8'h34; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_3225 = _T_2765 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3480 = _T_3479 | _T_3225; // @[Mux.scala 27:72]
  wire  _T_2767 = btb_rd_addr_f == 8'h35; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_3226 = _T_2767 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3481 = _T_3480 | _T_3226; // @[Mux.scala 27:72]
  wire  _T_2769 = btb_rd_addr_f == 8'h36; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_3227 = _T_2769 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3482 = _T_3481 | _T_3227; // @[Mux.scala 27:72]
  wire  _T_2771 = btb_rd_addr_f == 8'h37; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_3228 = _T_2771 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3483 = _T_3482 | _T_3228; // @[Mux.scala 27:72]
  wire  _T_2773 = btb_rd_addr_f == 8'h38; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_3229 = _T_2773 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3484 = _T_3483 | _T_3229; // @[Mux.scala 27:72]
  wire  _T_2775 = btb_rd_addr_f == 8'h39; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_3230 = _T_2775 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3485 = _T_3484 | _T_3230; // @[Mux.scala 27:72]
  wire  _T_2777 = btb_rd_addr_f == 8'h3a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_3231 = _T_2777 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3486 = _T_3485 | _T_3231; // @[Mux.scala 27:72]
  wire  _T_2779 = btb_rd_addr_f == 8'h3b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_3232 = _T_2779 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3487 = _T_3486 | _T_3232; // @[Mux.scala 27:72]
  wire  _T_2781 = btb_rd_addr_f == 8'h3c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_3233 = _T_2781 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3488 = _T_3487 | _T_3233; // @[Mux.scala 27:72]
  wire  _T_2783 = btb_rd_addr_f == 8'h3d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_3234 = _T_2783 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3489 = _T_3488 | _T_3234; // @[Mux.scala 27:72]
  wire  _T_2785 = btb_rd_addr_f == 8'h3e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_3235 = _T_2785 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3490 = _T_3489 | _T_3235; // @[Mux.scala 27:72]
  wire  _T_2787 = btb_rd_addr_f == 8'h3f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_3236 = _T_2787 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3491 = _T_3490 | _T_3236; // @[Mux.scala 27:72]
  wire  _T_2789 = btb_rd_addr_f == 8'h40; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_3237 = _T_2789 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3492 = _T_3491 | _T_3237; // @[Mux.scala 27:72]
  wire  _T_2791 = btb_rd_addr_f == 8'h41; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_3238 = _T_2791 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3493 = _T_3492 | _T_3238; // @[Mux.scala 27:72]
  wire  _T_2793 = btb_rd_addr_f == 8'h42; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_3239 = _T_2793 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3494 = _T_3493 | _T_3239; // @[Mux.scala 27:72]
  wire  _T_2795 = btb_rd_addr_f == 8'h43; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_3240 = _T_2795 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3495 = _T_3494 | _T_3240; // @[Mux.scala 27:72]
  wire  _T_2797 = btb_rd_addr_f == 8'h44; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_3241 = _T_2797 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3496 = _T_3495 | _T_3241; // @[Mux.scala 27:72]
  wire  _T_2799 = btb_rd_addr_f == 8'h45; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_3242 = _T_2799 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3497 = _T_3496 | _T_3242; // @[Mux.scala 27:72]
  wire  _T_2801 = btb_rd_addr_f == 8'h46; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_3243 = _T_2801 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3498 = _T_3497 | _T_3243; // @[Mux.scala 27:72]
  wire  _T_2803 = btb_rd_addr_f == 8'h47; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_3244 = _T_2803 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3499 = _T_3498 | _T_3244; // @[Mux.scala 27:72]
  wire  _T_2805 = btb_rd_addr_f == 8'h48; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_3245 = _T_2805 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3500 = _T_3499 | _T_3245; // @[Mux.scala 27:72]
  wire  _T_2807 = btb_rd_addr_f == 8'h49; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_3246 = _T_2807 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3501 = _T_3500 | _T_3246; // @[Mux.scala 27:72]
  wire  _T_2809 = btb_rd_addr_f == 8'h4a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_3247 = _T_2809 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3502 = _T_3501 | _T_3247; // @[Mux.scala 27:72]
  wire  _T_2811 = btb_rd_addr_f == 8'h4b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_3248 = _T_2811 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3503 = _T_3502 | _T_3248; // @[Mux.scala 27:72]
  wire  _T_2813 = btb_rd_addr_f == 8'h4c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_3249 = _T_2813 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3504 = _T_3503 | _T_3249; // @[Mux.scala 27:72]
  wire  _T_2815 = btb_rd_addr_f == 8'h4d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_3250 = _T_2815 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3505 = _T_3504 | _T_3250; // @[Mux.scala 27:72]
  wire  _T_2817 = btb_rd_addr_f == 8'h4e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_3251 = _T_2817 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3506 = _T_3505 | _T_3251; // @[Mux.scala 27:72]
  wire  _T_2819 = btb_rd_addr_f == 8'h4f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_3252 = _T_2819 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3507 = _T_3506 | _T_3252; // @[Mux.scala 27:72]
  wire  _T_2821 = btb_rd_addr_f == 8'h50; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_3253 = _T_2821 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3508 = _T_3507 | _T_3253; // @[Mux.scala 27:72]
  wire  _T_2823 = btb_rd_addr_f == 8'h51; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_3254 = _T_2823 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3509 = _T_3508 | _T_3254; // @[Mux.scala 27:72]
  wire  _T_2825 = btb_rd_addr_f == 8'h52; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_3255 = _T_2825 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3510 = _T_3509 | _T_3255; // @[Mux.scala 27:72]
  wire  _T_2827 = btb_rd_addr_f == 8'h53; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_3256 = _T_2827 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3511 = _T_3510 | _T_3256; // @[Mux.scala 27:72]
  wire  _T_2829 = btb_rd_addr_f == 8'h54; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_3257 = _T_2829 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3512 = _T_3511 | _T_3257; // @[Mux.scala 27:72]
  wire  _T_2831 = btb_rd_addr_f == 8'h55; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_3258 = _T_2831 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3513 = _T_3512 | _T_3258; // @[Mux.scala 27:72]
  wire  _T_2833 = btb_rd_addr_f == 8'h56; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_3259 = _T_2833 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3514 = _T_3513 | _T_3259; // @[Mux.scala 27:72]
  wire  _T_2835 = btb_rd_addr_f == 8'h57; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_3260 = _T_2835 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3515 = _T_3514 | _T_3260; // @[Mux.scala 27:72]
  wire  _T_2837 = btb_rd_addr_f == 8'h58; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_3261 = _T_2837 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3516 = _T_3515 | _T_3261; // @[Mux.scala 27:72]
  wire  _T_2839 = btb_rd_addr_f == 8'h59; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_3262 = _T_2839 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3517 = _T_3516 | _T_3262; // @[Mux.scala 27:72]
  wire  _T_2841 = btb_rd_addr_f == 8'h5a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_3263 = _T_2841 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3518 = _T_3517 | _T_3263; // @[Mux.scala 27:72]
  wire  _T_2843 = btb_rd_addr_f == 8'h5b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_3264 = _T_2843 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3519 = _T_3518 | _T_3264; // @[Mux.scala 27:72]
  wire  _T_2845 = btb_rd_addr_f == 8'h5c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_3265 = _T_2845 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3520 = _T_3519 | _T_3265; // @[Mux.scala 27:72]
  wire  _T_2847 = btb_rd_addr_f == 8'h5d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_3266 = _T_2847 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3521 = _T_3520 | _T_3266; // @[Mux.scala 27:72]
  wire  _T_2849 = btb_rd_addr_f == 8'h5e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_3267 = _T_2849 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3522 = _T_3521 | _T_3267; // @[Mux.scala 27:72]
  wire  _T_2851 = btb_rd_addr_f == 8'h5f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_3268 = _T_2851 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3523 = _T_3522 | _T_3268; // @[Mux.scala 27:72]
  wire  _T_2853 = btb_rd_addr_f == 8'h60; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_3269 = _T_2853 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3524 = _T_3523 | _T_3269; // @[Mux.scala 27:72]
  wire  _T_2855 = btb_rd_addr_f == 8'h61; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_3270 = _T_2855 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3525 = _T_3524 | _T_3270; // @[Mux.scala 27:72]
  wire  _T_2857 = btb_rd_addr_f == 8'h62; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_3271 = _T_2857 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3526 = _T_3525 | _T_3271; // @[Mux.scala 27:72]
  wire  _T_2859 = btb_rd_addr_f == 8'h63; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_3272 = _T_2859 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3527 = _T_3526 | _T_3272; // @[Mux.scala 27:72]
  wire  _T_2861 = btb_rd_addr_f == 8'h64; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_3273 = _T_2861 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3528 = _T_3527 | _T_3273; // @[Mux.scala 27:72]
  wire  _T_2863 = btb_rd_addr_f == 8'h65; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_3274 = _T_2863 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3529 = _T_3528 | _T_3274; // @[Mux.scala 27:72]
  wire  _T_2865 = btb_rd_addr_f == 8'h66; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_3275 = _T_2865 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3530 = _T_3529 | _T_3275; // @[Mux.scala 27:72]
  wire  _T_2867 = btb_rd_addr_f == 8'h67; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_3276 = _T_2867 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3531 = _T_3530 | _T_3276; // @[Mux.scala 27:72]
  wire  _T_2869 = btb_rd_addr_f == 8'h68; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_3277 = _T_2869 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3532 = _T_3531 | _T_3277; // @[Mux.scala 27:72]
  wire  _T_2871 = btb_rd_addr_f == 8'h69; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_3278 = _T_2871 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3533 = _T_3532 | _T_3278; // @[Mux.scala 27:72]
  wire  _T_2873 = btb_rd_addr_f == 8'h6a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_3279 = _T_2873 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3534 = _T_3533 | _T_3279; // @[Mux.scala 27:72]
  wire  _T_2875 = btb_rd_addr_f == 8'h6b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_3280 = _T_2875 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3535 = _T_3534 | _T_3280; // @[Mux.scala 27:72]
  wire  _T_2877 = btb_rd_addr_f == 8'h6c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_3281 = _T_2877 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3536 = _T_3535 | _T_3281; // @[Mux.scala 27:72]
  wire  _T_2879 = btb_rd_addr_f == 8'h6d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_3282 = _T_2879 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3537 = _T_3536 | _T_3282; // @[Mux.scala 27:72]
  wire  _T_2881 = btb_rd_addr_f == 8'h6e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_3283 = _T_2881 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3538 = _T_3537 | _T_3283; // @[Mux.scala 27:72]
  wire  _T_2883 = btb_rd_addr_f == 8'h6f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_3284 = _T_2883 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3539 = _T_3538 | _T_3284; // @[Mux.scala 27:72]
  wire  _T_2885 = btb_rd_addr_f == 8'h70; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_3285 = _T_2885 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3540 = _T_3539 | _T_3285; // @[Mux.scala 27:72]
  wire  _T_2887 = btb_rd_addr_f == 8'h71; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_3286 = _T_2887 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3541 = _T_3540 | _T_3286; // @[Mux.scala 27:72]
  wire  _T_2889 = btb_rd_addr_f == 8'h72; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_3287 = _T_2889 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3542 = _T_3541 | _T_3287; // @[Mux.scala 27:72]
  wire  _T_2891 = btb_rd_addr_f == 8'h73; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_3288 = _T_2891 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3543 = _T_3542 | _T_3288; // @[Mux.scala 27:72]
  wire  _T_2893 = btb_rd_addr_f == 8'h74; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_3289 = _T_2893 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3544 = _T_3543 | _T_3289; // @[Mux.scala 27:72]
  wire  _T_2895 = btb_rd_addr_f == 8'h75; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_3290 = _T_2895 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3545 = _T_3544 | _T_3290; // @[Mux.scala 27:72]
  wire  _T_2897 = btb_rd_addr_f == 8'h76; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_3291 = _T_2897 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3546 = _T_3545 | _T_3291; // @[Mux.scala 27:72]
  wire  _T_2899 = btb_rd_addr_f == 8'h77; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_3292 = _T_2899 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3547 = _T_3546 | _T_3292; // @[Mux.scala 27:72]
  wire  _T_2901 = btb_rd_addr_f == 8'h78; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_3293 = _T_2901 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3548 = _T_3547 | _T_3293; // @[Mux.scala 27:72]
  wire  _T_2903 = btb_rd_addr_f == 8'h79; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_3294 = _T_2903 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3549 = _T_3548 | _T_3294; // @[Mux.scala 27:72]
  wire  _T_2905 = btb_rd_addr_f == 8'h7a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_3295 = _T_2905 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3550 = _T_3549 | _T_3295; // @[Mux.scala 27:72]
  wire  _T_2907 = btb_rd_addr_f == 8'h7b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_3296 = _T_2907 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3551 = _T_3550 | _T_3296; // @[Mux.scala 27:72]
  wire  _T_2909 = btb_rd_addr_f == 8'h7c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_3297 = _T_2909 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3552 = _T_3551 | _T_3297; // @[Mux.scala 27:72]
  wire  _T_2911 = btb_rd_addr_f == 8'h7d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_3298 = _T_2911 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3553 = _T_3552 | _T_3298; // @[Mux.scala 27:72]
  wire  _T_2913 = btb_rd_addr_f == 8'h7e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_3299 = _T_2913 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3554 = _T_3553 | _T_3299; // @[Mux.scala 27:72]
  wire  _T_2915 = btb_rd_addr_f == 8'h7f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_3300 = _T_2915 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3555 = _T_3554 | _T_3300; // @[Mux.scala 27:72]
  wire  _T_2917 = btb_rd_addr_f == 8'h80; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_3301 = _T_2917 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3556 = _T_3555 | _T_3301; // @[Mux.scala 27:72]
  wire  _T_2919 = btb_rd_addr_f == 8'h81; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_3302 = _T_2919 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3557 = _T_3556 | _T_3302; // @[Mux.scala 27:72]
  wire  _T_2921 = btb_rd_addr_f == 8'h82; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_3303 = _T_2921 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3558 = _T_3557 | _T_3303; // @[Mux.scala 27:72]
  wire  _T_2923 = btb_rd_addr_f == 8'h83; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_3304 = _T_2923 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3559 = _T_3558 | _T_3304; // @[Mux.scala 27:72]
  wire  _T_2925 = btb_rd_addr_f == 8'h84; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_3305 = _T_2925 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3560 = _T_3559 | _T_3305; // @[Mux.scala 27:72]
  wire  _T_2927 = btb_rd_addr_f == 8'h85; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_3306 = _T_2927 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3561 = _T_3560 | _T_3306; // @[Mux.scala 27:72]
  wire  _T_2929 = btb_rd_addr_f == 8'h86; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_3307 = _T_2929 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3562 = _T_3561 | _T_3307; // @[Mux.scala 27:72]
  wire  _T_2931 = btb_rd_addr_f == 8'h87; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_3308 = _T_2931 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3563 = _T_3562 | _T_3308; // @[Mux.scala 27:72]
  wire  _T_2933 = btb_rd_addr_f == 8'h88; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_3309 = _T_2933 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3564 = _T_3563 | _T_3309; // @[Mux.scala 27:72]
  wire  _T_2935 = btb_rd_addr_f == 8'h89; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_3310 = _T_2935 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3565 = _T_3564 | _T_3310; // @[Mux.scala 27:72]
  wire  _T_2937 = btb_rd_addr_f == 8'h8a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_3311 = _T_2937 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3566 = _T_3565 | _T_3311; // @[Mux.scala 27:72]
  wire  _T_2939 = btb_rd_addr_f == 8'h8b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_3312 = _T_2939 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3567 = _T_3566 | _T_3312; // @[Mux.scala 27:72]
  wire  _T_2941 = btb_rd_addr_f == 8'h8c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_3313 = _T_2941 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3568 = _T_3567 | _T_3313; // @[Mux.scala 27:72]
  wire  _T_2943 = btb_rd_addr_f == 8'h8d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_3314 = _T_2943 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3569 = _T_3568 | _T_3314; // @[Mux.scala 27:72]
  wire  _T_2945 = btb_rd_addr_f == 8'h8e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_3315 = _T_2945 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3570 = _T_3569 | _T_3315; // @[Mux.scala 27:72]
  wire  _T_2947 = btb_rd_addr_f == 8'h8f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_3316 = _T_2947 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3571 = _T_3570 | _T_3316; // @[Mux.scala 27:72]
  wire  _T_2949 = btb_rd_addr_f == 8'h90; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_3317 = _T_2949 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3572 = _T_3571 | _T_3317; // @[Mux.scala 27:72]
  wire  _T_2951 = btb_rd_addr_f == 8'h91; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_3318 = _T_2951 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3573 = _T_3572 | _T_3318; // @[Mux.scala 27:72]
  wire  _T_2953 = btb_rd_addr_f == 8'h92; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_3319 = _T_2953 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3574 = _T_3573 | _T_3319; // @[Mux.scala 27:72]
  wire  _T_2955 = btb_rd_addr_f == 8'h93; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_3320 = _T_2955 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3575 = _T_3574 | _T_3320; // @[Mux.scala 27:72]
  wire  _T_2957 = btb_rd_addr_f == 8'h94; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_3321 = _T_2957 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3576 = _T_3575 | _T_3321; // @[Mux.scala 27:72]
  wire  _T_2959 = btb_rd_addr_f == 8'h95; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_3322 = _T_2959 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3577 = _T_3576 | _T_3322; // @[Mux.scala 27:72]
  wire  _T_2961 = btb_rd_addr_f == 8'h96; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_3323 = _T_2961 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3578 = _T_3577 | _T_3323; // @[Mux.scala 27:72]
  wire  _T_2963 = btb_rd_addr_f == 8'h97; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_3324 = _T_2963 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3579 = _T_3578 | _T_3324; // @[Mux.scala 27:72]
  wire  _T_2965 = btb_rd_addr_f == 8'h98; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_3325 = _T_2965 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3580 = _T_3579 | _T_3325; // @[Mux.scala 27:72]
  wire  _T_2967 = btb_rd_addr_f == 8'h99; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_3326 = _T_2967 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3581 = _T_3580 | _T_3326; // @[Mux.scala 27:72]
  wire  _T_2969 = btb_rd_addr_f == 8'h9a; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_3327 = _T_2969 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3582 = _T_3581 | _T_3327; // @[Mux.scala 27:72]
  wire  _T_2971 = btb_rd_addr_f == 8'h9b; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_3328 = _T_2971 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3583 = _T_3582 | _T_3328; // @[Mux.scala 27:72]
  wire  _T_2973 = btb_rd_addr_f == 8'h9c; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_3329 = _T_2973 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3584 = _T_3583 | _T_3329; // @[Mux.scala 27:72]
  wire  _T_2975 = btb_rd_addr_f == 8'h9d; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_3330 = _T_2975 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3585 = _T_3584 | _T_3330; // @[Mux.scala 27:72]
  wire  _T_2977 = btb_rd_addr_f == 8'h9e; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_3331 = _T_2977 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3586 = _T_3585 | _T_3331; // @[Mux.scala 27:72]
  wire  _T_2979 = btb_rd_addr_f == 8'h9f; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_3332 = _T_2979 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3587 = _T_3586 | _T_3332; // @[Mux.scala 27:72]
  wire  _T_2981 = btb_rd_addr_f == 8'ha0; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_3333 = _T_2981 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3588 = _T_3587 | _T_3333; // @[Mux.scala 27:72]
  wire  _T_2983 = btb_rd_addr_f == 8'ha1; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_3334 = _T_2983 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3589 = _T_3588 | _T_3334; // @[Mux.scala 27:72]
  wire  _T_2985 = btb_rd_addr_f == 8'ha2; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_3335 = _T_2985 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3590 = _T_3589 | _T_3335; // @[Mux.scala 27:72]
  wire  _T_2987 = btb_rd_addr_f == 8'ha3; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_3336 = _T_2987 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3591 = _T_3590 | _T_3336; // @[Mux.scala 27:72]
  wire  _T_2989 = btb_rd_addr_f == 8'ha4; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_3337 = _T_2989 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3592 = _T_3591 | _T_3337; // @[Mux.scala 27:72]
  wire  _T_2991 = btb_rd_addr_f == 8'ha5; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_3338 = _T_2991 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3593 = _T_3592 | _T_3338; // @[Mux.scala 27:72]
  wire  _T_2993 = btb_rd_addr_f == 8'ha6; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_3339 = _T_2993 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3594 = _T_3593 | _T_3339; // @[Mux.scala 27:72]
  wire  _T_2995 = btb_rd_addr_f == 8'ha7; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_3340 = _T_2995 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3595 = _T_3594 | _T_3340; // @[Mux.scala 27:72]
  wire  _T_2997 = btb_rd_addr_f == 8'ha8; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_3341 = _T_2997 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3596 = _T_3595 | _T_3341; // @[Mux.scala 27:72]
  wire  _T_2999 = btb_rd_addr_f == 8'ha9; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_3342 = _T_2999 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3597 = _T_3596 | _T_3342; // @[Mux.scala 27:72]
  wire  _T_3001 = btb_rd_addr_f == 8'haa; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_3343 = _T_3001 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3598 = _T_3597 | _T_3343; // @[Mux.scala 27:72]
  wire  _T_3003 = btb_rd_addr_f == 8'hab; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_3344 = _T_3003 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3599 = _T_3598 | _T_3344; // @[Mux.scala 27:72]
  wire  _T_3005 = btb_rd_addr_f == 8'hac; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_3345 = _T_3005 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3600 = _T_3599 | _T_3345; // @[Mux.scala 27:72]
  wire  _T_3007 = btb_rd_addr_f == 8'had; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_3346 = _T_3007 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3601 = _T_3600 | _T_3346; // @[Mux.scala 27:72]
  wire  _T_3009 = btb_rd_addr_f == 8'hae; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_3347 = _T_3009 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3602 = _T_3601 | _T_3347; // @[Mux.scala 27:72]
  wire  _T_3011 = btb_rd_addr_f == 8'haf; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_3348 = _T_3011 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3603 = _T_3602 | _T_3348; // @[Mux.scala 27:72]
  wire  _T_3013 = btb_rd_addr_f == 8'hb0; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_3349 = _T_3013 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3604 = _T_3603 | _T_3349; // @[Mux.scala 27:72]
  wire  _T_3015 = btb_rd_addr_f == 8'hb1; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_3350 = _T_3015 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3605 = _T_3604 | _T_3350; // @[Mux.scala 27:72]
  wire  _T_3017 = btb_rd_addr_f == 8'hb2; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_3351 = _T_3017 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3606 = _T_3605 | _T_3351; // @[Mux.scala 27:72]
  wire  _T_3019 = btb_rd_addr_f == 8'hb3; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_3352 = _T_3019 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3607 = _T_3606 | _T_3352; // @[Mux.scala 27:72]
  wire  _T_3021 = btb_rd_addr_f == 8'hb4; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_3353 = _T_3021 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3608 = _T_3607 | _T_3353; // @[Mux.scala 27:72]
  wire  _T_3023 = btb_rd_addr_f == 8'hb5; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_3354 = _T_3023 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3609 = _T_3608 | _T_3354; // @[Mux.scala 27:72]
  wire  _T_3025 = btb_rd_addr_f == 8'hb6; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_3355 = _T_3025 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3610 = _T_3609 | _T_3355; // @[Mux.scala 27:72]
  wire  _T_3027 = btb_rd_addr_f == 8'hb7; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_3356 = _T_3027 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3611 = _T_3610 | _T_3356; // @[Mux.scala 27:72]
  wire  _T_3029 = btb_rd_addr_f == 8'hb8; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_3357 = _T_3029 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3612 = _T_3611 | _T_3357; // @[Mux.scala 27:72]
  wire  _T_3031 = btb_rd_addr_f == 8'hb9; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_3358 = _T_3031 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3613 = _T_3612 | _T_3358; // @[Mux.scala 27:72]
  wire  _T_3033 = btb_rd_addr_f == 8'hba; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_3359 = _T_3033 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3614 = _T_3613 | _T_3359; // @[Mux.scala 27:72]
  wire  _T_3035 = btb_rd_addr_f == 8'hbb; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_3360 = _T_3035 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3615 = _T_3614 | _T_3360; // @[Mux.scala 27:72]
  wire  _T_3037 = btb_rd_addr_f == 8'hbc; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_3361 = _T_3037 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3616 = _T_3615 | _T_3361; // @[Mux.scala 27:72]
  wire  _T_3039 = btb_rd_addr_f == 8'hbd; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_3362 = _T_3039 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3617 = _T_3616 | _T_3362; // @[Mux.scala 27:72]
  wire  _T_3041 = btb_rd_addr_f == 8'hbe; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_3363 = _T_3041 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3618 = _T_3617 | _T_3363; // @[Mux.scala 27:72]
  wire  _T_3043 = btb_rd_addr_f == 8'hbf; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_3364 = _T_3043 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3619 = _T_3618 | _T_3364; // @[Mux.scala 27:72]
  wire  _T_3045 = btb_rd_addr_f == 8'hc0; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_3365 = _T_3045 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3620 = _T_3619 | _T_3365; // @[Mux.scala 27:72]
  wire  _T_3047 = btb_rd_addr_f == 8'hc1; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_3366 = _T_3047 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3621 = _T_3620 | _T_3366; // @[Mux.scala 27:72]
  wire  _T_3049 = btb_rd_addr_f == 8'hc2; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_3367 = _T_3049 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3622 = _T_3621 | _T_3367; // @[Mux.scala 27:72]
  wire  _T_3051 = btb_rd_addr_f == 8'hc3; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_3368 = _T_3051 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3623 = _T_3622 | _T_3368; // @[Mux.scala 27:72]
  wire  _T_3053 = btb_rd_addr_f == 8'hc4; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_3369 = _T_3053 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3624 = _T_3623 | _T_3369; // @[Mux.scala 27:72]
  wire  _T_3055 = btb_rd_addr_f == 8'hc5; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_3370 = _T_3055 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3625 = _T_3624 | _T_3370; // @[Mux.scala 27:72]
  wire  _T_3057 = btb_rd_addr_f == 8'hc6; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_3371 = _T_3057 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3626 = _T_3625 | _T_3371; // @[Mux.scala 27:72]
  wire  _T_3059 = btb_rd_addr_f == 8'hc7; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_3372 = _T_3059 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3627 = _T_3626 | _T_3372; // @[Mux.scala 27:72]
  wire  _T_3061 = btb_rd_addr_f == 8'hc8; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_3373 = _T_3061 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3628 = _T_3627 | _T_3373; // @[Mux.scala 27:72]
  wire  _T_3063 = btb_rd_addr_f == 8'hc9; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_3374 = _T_3063 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3629 = _T_3628 | _T_3374; // @[Mux.scala 27:72]
  wire  _T_3065 = btb_rd_addr_f == 8'hca; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_3375 = _T_3065 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3630 = _T_3629 | _T_3375; // @[Mux.scala 27:72]
  wire  _T_3067 = btb_rd_addr_f == 8'hcb; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_3376 = _T_3067 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3631 = _T_3630 | _T_3376; // @[Mux.scala 27:72]
  wire  _T_3069 = btb_rd_addr_f == 8'hcc; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_3377 = _T_3069 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3632 = _T_3631 | _T_3377; // @[Mux.scala 27:72]
  wire  _T_3071 = btb_rd_addr_f == 8'hcd; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_3378 = _T_3071 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3633 = _T_3632 | _T_3378; // @[Mux.scala 27:72]
  wire  _T_3073 = btb_rd_addr_f == 8'hce; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_3379 = _T_3073 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3634 = _T_3633 | _T_3379; // @[Mux.scala 27:72]
  wire  _T_3075 = btb_rd_addr_f == 8'hcf; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_3380 = _T_3075 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3635 = _T_3634 | _T_3380; // @[Mux.scala 27:72]
  wire  _T_3077 = btb_rd_addr_f == 8'hd0; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_3381 = _T_3077 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3636 = _T_3635 | _T_3381; // @[Mux.scala 27:72]
  wire  _T_3079 = btb_rd_addr_f == 8'hd1; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_3382 = _T_3079 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3637 = _T_3636 | _T_3382; // @[Mux.scala 27:72]
  wire  _T_3081 = btb_rd_addr_f == 8'hd2; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_3383 = _T_3081 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3638 = _T_3637 | _T_3383; // @[Mux.scala 27:72]
  wire  _T_3083 = btb_rd_addr_f == 8'hd3; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_3384 = _T_3083 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3639 = _T_3638 | _T_3384; // @[Mux.scala 27:72]
  wire  _T_3085 = btb_rd_addr_f == 8'hd4; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_3385 = _T_3085 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3640 = _T_3639 | _T_3385; // @[Mux.scala 27:72]
  wire  _T_3087 = btb_rd_addr_f == 8'hd5; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_3386 = _T_3087 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3641 = _T_3640 | _T_3386; // @[Mux.scala 27:72]
  wire  _T_3089 = btb_rd_addr_f == 8'hd6; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_3387 = _T_3089 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3642 = _T_3641 | _T_3387; // @[Mux.scala 27:72]
  wire  _T_3091 = btb_rd_addr_f == 8'hd7; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_3388 = _T_3091 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3643 = _T_3642 | _T_3388; // @[Mux.scala 27:72]
  wire  _T_3093 = btb_rd_addr_f == 8'hd8; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_3389 = _T_3093 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3644 = _T_3643 | _T_3389; // @[Mux.scala 27:72]
  wire  _T_3095 = btb_rd_addr_f == 8'hd9; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_3390 = _T_3095 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3645 = _T_3644 | _T_3390; // @[Mux.scala 27:72]
  wire  _T_3097 = btb_rd_addr_f == 8'hda; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_3391 = _T_3097 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3646 = _T_3645 | _T_3391; // @[Mux.scala 27:72]
  wire  _T_3099 = btb_rd_addr_f == 8'hdb; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_3392 = _T_3099 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3647 = _T_3646 | _T_3392; // @[Mux.scala 27:72]
  wire  _T_3101 = btb_rd_addr_f == 8'hdc; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_3393 = _T_3101 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3648 = _T_3647 | _T_3393; // @[Mux.scala 27:72]
  wire  _T_3103 = btb_rd_addr_f == 8'hdd; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_3394 = _T_3103 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3649 = _T_3648 | _T_3394; // @[Mux.scala 27:72]
  wire  _T_3105 = btb_rd_addr_f == 8'hde; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_3395 = _T_3105 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3650 = _T_3649 | _T_3395; // @[Mux.scala 27:72]
  wire  _T_3107 = btb_rd_addr_f == 8'hdf; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_3396 = _T_3107 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3651 = _T_3650 | _T_3396; // @[Mux.scala 27:72]
  wire  _T_3109 = btb_rd_addr_f == 8'he0; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_3397 = _T_3109 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3652 = _T_3651 | _T_3397; // @[Mux.scala 27:72]
  wire  _T_3111 = btb_rd_addr_f == 8'he1; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_3398 = _T_3111 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3653 = _T_3652 | _T_3398; // @[Mux.scala 27:72]
  wire  _T_3113 = btb_rd_addr_f == 8'he2; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_3399 = _T_3113 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3654 = _T_3653 | _T_3399; // @[Mux.scala 27:72]
  wire  _T_3115 = btb_rd_addr_f == 8'he3; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_3400 = _T_3115 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3655 = _T_3654 | _T_3400; // @[Mux.scala 27:72]
  wire  _T_3117 = btb_rd_addr_f == 8'he4; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_3401 = _T_3117 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3656 = _T_3655 | _T_3401; // @[Mux.scala 27:72]
  wire  _T_3119 = btb_rd_addr_f == 8'he5; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_3402 = _T_3119 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3657 = _T_3656 | _T_3402; // @[Mux.scala 27:72]
  wire  _T_3121 = btb_rd_addr_f == 8'he6; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_3403 = _T_3121 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3658 = _T_3657 | _T_3403; // @[Mux.scala 27:72]
  wire  _T_3123 = btb_rd_addr_f == 8'he7; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_3404 = _T_3123 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3659 = _T_3658 | _T_3404; // @[Mux.scala 27:72]
  wire  _T_3125 = btb_rd_addr_f == 8'he8; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_3405 = _T_3125 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3660 = _T_3659 | _T_3405; // @[Mux.scala 27:72]
  wire  _T_3127 = btb_rd_addr_f == 8'he9; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_3406 = _T_3127 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3661 = _T_3660 | _T_3406; // @[Mux.scala 27:72]
  wire  _T_3129 = btb_rd_addr_f == 8'hea; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_3407 = _T_3129 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3662 = _T_3661 | _T_3407; // @[Mux.scala 27:72]
  wire  _T_3131 = btb_rd_addr_f == 8'heb; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_3408 = _T_3131 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3663 = _T_3662 | _T_3408; // @[Mux.scala 27:72]
  wire  _T_3133 = btb_rd_addr_f == 8'hec; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_3409 = _T_3133 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3664 = _T_3663 | _T_3409; // @[Mux.scala 27:72]
  wire  _T_3135 = btb_rd_addr_f == 8'hed; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_3410 = _T_3135 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3665 = _T_3664 | _T_3410; // @[Mux.scala 27:72]
  wire  _T_3137 = btb_rd_addr_f == 8'hee; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_3411 = _T_3137 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3666 = _T_3665 | _T_3411; // @[Mux.scala 27:72]
  wire  _T_3139 = btb_rd_addr_f == 8'hef; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_3412 = _T_3139 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3667 = _T_3666 | _T_3412; // @[Mux.scala 27:72]
  wire  _T_3141 = btb_rd_addr_f == 8'hf0; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_3413 = _T_3141 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3668 = _T_3667 | _T_3413; // @[Mux.scala 27:72]
  wire  _T_3143 = btb_rd_addr_f == 8'hf1; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_3414 = _T_3143 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3669 = _T_3668 | _T_3414; // @[Mux.scala 27:72]
  wire  _T_3145 = btb_rd_addr_f == 8'hf2; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_3415 = _T_3145 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3670 = _T_3669 | _T_3415; // @[Mux.scala 27:72]
  wire  _T_3147 = btb_rd_addr_f == 8'hf3; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_3416 = _T_3147 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3671 = _T_3670 | _T_3416; // @[Mux.scala 27:72]
  wire  _T_3149 = btb_rd_addr_f == 8'hf4; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_3417 = _T_3149 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3672 = _T_3671 | _T_3417; // @[Mux.scala 27:72]
  wire  _T_3151 = btb_rd_addr_f == 8'hf5; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_3418 = _T_3151 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3673 = _T_3672 | _T_3418; // @[Mux.scala 27:72]
  wire  _T_3153 = btb_rd_addr_f == 8'hf6; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_3419 = _T_3153 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3674 = _T_3673 | _T_3419; // @[Mux.scala 27:72]
  wire  _T_3155 = btb_rd_addr_f == 8'hf7; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_3420 = _T_3155 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3675 = _T_3674 | _T_3420; // @[Mux.scala 27:72]
  wire  _T_3157 = btb_rd_addr_f == 8'hf8; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_3421 = _T_3157 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3676 = _T_3675 | _T_3421; // @[Mux.scala 27:72]
  wire  _T_3159 = btb_rd_addr_f == 8'hf9; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_3422 = _T_3159 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3677 = _T_3676 | _T_3422; // @[Mux.scala 27:72]
  wire  _T_3161 = btb_rd_addr_f == 8'hfa; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_3423 = _T_3161 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3678 = _T_3677 | _T_3423; // @[Mux.scala 27:72]
  wire  _T_3163 = btb_rd_addr_f == 8'hfb; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_3424 = _T_3163 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3679 = _T_3678 | _T_3424; // @[Mux.scala 27:72]
  wire  _T_3165 = btb_rd_addr_f == 8'hfc; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_3425 = _T_3165 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3680 = _T_3679 | _T_3425; // @[Mux.scala 27:72]
  wire  _T_3167 = btb_rd_addr_f == 8'hfd; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_3426 = _T_3167 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3681 = _T_3680 | _T_3426; // @[Mux.scala 27:72]
  wire  _T_3169 = btb_rd_addr_f == 8'hfe; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_3427 = _T_3169 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_3682 = _T_3681 | _T_3427; // @[Mux.scala 27:72]
  wire  _T_3171 = btb_rd_addr_f == 8'hff; // @[ifu_bp_ctl.scala 436:80]
  reg [21:0] btb_bank0_rd_data_way0_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_3428 = _T_3171 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_f = _T_3682 | _T_3428; // @[Mux.scala 27:72]
  wire [4:0] _T_29 = io_ifc_fetch_addr_f[13:9] ^ io_ifc_fetch_addr_f[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_f = _T_29 ^ io_ifc_fetch_addr_f[23:19]; // @[lib.scala 42:111]
  wire  _T_46 = btb_bank0_rd_data_way0_f[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 144:98]
  wire  _T_47 = btb_bank0_rd_data_way0_f[0] & _T_46; // @[ifu_bp_ctl.scala 144:55]
  wire  _T_19 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_f; // @[ifu_bp_ctl.scala 125:72]
  wire  branch_error_collision_f = dec_tlu_error_wb & _T_19; // @[ifu_bp_ctl.scala 125:51]
  wire  branch_error_bank_conflict_f = branch_error_collision_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 129:63]
  wire  _T_48 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & branch_error_bank_conflict_f; // @[ifu_bp_ctl.scala 145:22]
  wire  _T_49 = ~_T_48; // @[ifu_bp_ctl.scala 145:5]
  wire  _T_50 = _T_47 & _T_49; // @[ifu_bp_ctl.scala 144:118]
  wire  _T_51 = _T_50 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 145:54]
  wire  tag_match_way0_f = _T_51 & _T; // @[ifu_bp_ctl.scala 145:75]
  wire  _T_82 = btb_bank0_rd_data_way0_f[3] ^ btb_bank0_rd_data_way0_f[4]; // @[ifu_bp_ctl.scala 159:90]
  wire  _T_83 = tag_match_way0_f & _T_82; // @[ifu_bp_ctl.scala 159:56]
  wire  _T_87 = ~_T_82; // @[ifu_bp_ctl.scala 160:24]
  wire  _T_88 = tag_match_way0_f & _T_87; // @[ifu_bp_ctl.scala 160:22]
  wire [1:0] tag_match_way0_expanded_f = {_T_83,_T_88}; // @[Cat.scala 29:58]
  wire [21:0] _T_129 = tag_match_way0_expanded_f[1] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_0; // @[Reg.scala 27:20]
  wire [21:0] _T_4197 = _T_2661 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_1; // @[Reg.scala 27:20]
  wire [21:0] _T_4198 = _T_2663 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4453 = _T_4197 | _T_4198; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_2; // @[Reg.scala 27:20]
  wire [21:0] _T_4199 = _T_2665 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4454 = _T_4453 | _T_4199; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_3; // @[Reg.scala 27:20]
  wire [21:0] _T_4200 = _T_2667 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4455 = _T_4454 | _T_4200; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_4; // @[Reg.scala 27:20]
  wire [21:0] _T_4201 = _T_2669 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4456 = _T_4455 | _T_4201; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_5; // @[Reg.scala 27:20]
  wire [21:0] _T_4202 = _T_2671 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4457 = _T_4456 | _T_4202; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_6; // @[Reg.scala 27:20]
  wire [21:0] _T_4203 = _T_2673 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4458 = _T_4457 | _T_4203; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_7; // @[Reg.scala 27:20]
  wire [21:0] _T_4204 = _T_2675 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4459 = _T_4458 | _T_4204; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_8; // @[Reg.scala 27:20]
  wire [21:0] _T_4205 = _T_2677 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4460 = _T_4459 | _T_4205; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_9; // @[Reg.scala 27:20]
  wire [21:0] _T_4206 = _T_2679 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4461 = _T_4460 | _T_4206; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_10; // @[Reg.scala 27:20]
  wire [21:0] _T_4207 = _T_2681 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4462 = _T_4461 | _T_4207; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_11; // @[Reg.scala 27:20]
  wire [21:0] _T_4208 = _T_2683 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4463 = _T_4462 | _T_4208; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_12; // @[Reg.scala 27:20]
  wire [21:0] _T_4209 = _T_2685 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4464 = _T_4463 | _T_4209; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_13; // @[Reg.scala 27:20]
  wire [21:0] _T_4210 = _T_2687 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4465 = _T_4464 | _T_4210; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_14; // @[Reg.scala 27:20]
  wire [21:0] _T_4211 = _T_2689 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4466 = _T_4465 | _T_4211; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_15; // @[Reg.scala 27:20]
  wire [21:0] _T_4212 = _T_2691 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4467 = _T_4466 | _T_4212; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_16; // @[Reg.scala 27:20]
  wire [21:0] _T_4213 = _T_2693 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4468 = _T_4467 | _T_4213; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_17; // @[Reg.scala 27:20]
  wire [21:0] _T_4214 = _T_2695 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4469 = _T_4468 | _T_4214; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_18; // @[Reg.scala 27:20]
  wire [21:0] _T_4215 = _T_2697 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4470 = _T_4469 | _T_4215; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_19; // @[Reg.scala 27:20]
  wire [21:0] _T_4216 = _T_2699 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4471 = _T_4470 | _T_4216; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_20; // @[Reg.scala 27:20]
  wire [21:0] _T_4217 = _T_2701 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4472 = _T_4471 | _T_4217; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_21; // @[Reg.scala 27:20]
  wire [21:0] _T_4218 = _T_2703 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4473 = _T_4472 | _T_4218; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_22; // @[Reg.scala 27:20]
  wire [21:0] _T_4219 = _T_2705 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4474 = _T_4473 | _T_4219; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_23; // @[Reg.scala 27:20]
  wire [21:0] _T_4220 = _T_2707 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4475 = _T_4474 | _T_4220; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_24; // @[Reg.scala 27:20]
  wire [21:0] _T_4221 = _T_2709 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4476 = _T_4475 | _T_4221; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_25; // @[Reg.scala 27:20]
  wire [21:0] _T_4222 = _T_2711 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4477 = _T_4476 | _T_4222; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_26; // @[Reg.scala 27:20]
  wire [21:0] _T_4223 = _T_2713 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4478 = _T_4477 | _T_4223; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_27; // @[Reg.scala 27:20]
  wire [21:0] _T_4224 = _T_2715 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4479 = _T_4478 | _T_4224; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_28; // @[Reg.scala 27:20]
  wire [21:0] _T_4225 = _T_2717 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4480 = _T_4479 | _T_4225; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_29; // @[Reg.scala 27:20]
  wire [21:0] _T_4226 = _T_2719 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4481 = _T_4480 | _T_4226; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_30; // @[Reg.scala 27:20]
  wire [21:0] _T_4227 = _T_2721 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4482 = _T_4481 | _T_4227; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_31; // @[Reg.scala 27:20]
  wire [21:0] _T_4228 = _T_2723 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4483 = _T_4482 | _T_4228; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_32; // @[Reg.scala 27:20]
  wire [21:0] _T_4229 = _T_2725 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4484 = _T_4483 | _T_4229; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_33; // @[Reg.scala 27:20]
  wire [21:0] _T_4230 = _T_2727 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4485 = _T_4484 | _T_4230; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_34; // @[Reg.scala 27:20]
  wire [21:0] _T_4231 = _T_2729 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4486 = _T_4485 | _T_4231; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_35; // @[Reg.scala 27:20]
  wire [21:0] _T_4232 = _T_2731 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4487 = _T_4486 | _T_4232; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_36; // @[Reg.scala 27:20]
  wire [21:0] _T_4233 = _T_2733 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4488 = _T_4487 | _T_4233; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_37; // @[Reg.scala 27:20]
  wire [21:0] _T_4234 = _T_2735 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4489 = _T_4488 | _T_4234; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_38; // @[Reg.scala 27:20]
  wire [21:0] _T_4235 = _T_2737 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4490 = _T_4489 | _T_4235; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_39; // @[Reg.scala 27:20]
  wire [21:0] _T_4236 = _T_2739 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4491 = _T_4490 | _T_4236; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_40; // @[Reg.scala 27:20]
  wire [21:0] _T_4237 = _T_2741 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4492 = _T_4491 | _T_4237; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_41; // @[Reg.scala 27:20]
  wire [21:0] _T_4238 = _T_2743 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4493 = _T_4492 | _T_4238; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_42; // @[Reg.scala 27:20]
  wire [21:0] _T_4239 = _T_2745 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4494 = _T_4493 | _T_4239; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_43; // @[Reg.scala 27:20]
  wire [21:0] _T_4240 = _T_2747 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4495 = _T_4494 | _T_4240; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_44; // @[Reg.scala 27:20]
  wire [21:0] _T_4241 = _T_2749 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4496 = _T_4495 | _T_4241; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_45; // @[Reg.scala 27:20]
  wire [21:0] _T_4242 = _T_2751 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4497 = _T_4496 | _T_4242; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_46; // @[Reg.scala 27:20]
  wire [21:0] _T_4243 = _T_2753 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4498 = _T_4497 | _T_4243; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_47; // @[Reg.scala 27:20]
  wire [21:0] _T_4244 = _T_2755 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4499 = _T_4498 | _T_4244; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_48; // @[Reg.scala 27:20]
  wire [21:0] _T_4245 = _T_2757 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4500 = _T_4499 | _T_4245; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_49; // @[Reg.scala 27:20]
  wire [21:0] _T_4246 = _T_2759 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4501 = _T_4500 | _T_4246; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_50; // @[Reg.scala 27:20]
  wire [21:0] _T_4247 = _T_2761 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4502 = _T_4501 | _T_4247; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_51; // @[Reg.scala 27:20]
  wire [21:0] _T_4248 = _T_2763 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4503 = _T_4502 | _T_4248; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_52; // @[Reg.scala 27:20]
  wire [21:0] _T_4249 = _T_2765 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4504 = _T_4503 | _T_4249; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_53; // @[Reg.scala 27:20]
  wire [21:0] _T_4250 = _T_2767 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4505 = _T_4504 | _T_4250; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_54; // @[Reg.scala 27:20]
  wire [21:0] _T_4251 = _T_2769 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4506 = _T_4505 | _T_4251; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_55; // @[Reg.scala 27:20]
  wire [21:0] _T_4252 = _T_2771 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4507 = _T_4506 | _T_4252; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_56; // @[Reg.scala 27:20]
  wire [21:0] _T_4253 = _T_2773 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4508 = _T_4507 | _T_4253; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_57; // @[Reg.scala 27:20]
  wire [21:0] _T_4254 = _T_2775 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4509 = _T_4508 | _T_4254; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_58; // @[Reg.scala 27:20]
  wire [21:0] _T_4255 = _T_2777 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4510 = _T_4509 | _T_4255; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_59; // @[Reg.scala 27:20]
  wire [21:0] _T_4256 = _T_2779 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4511 = _T_4510 | _T_4256; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_60; // @[Reg.scala 27:20]
  wire [21:0] _T_4257 = _T_2781 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4512 = _T_4511 | _T_4257; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_61; // @[Reg.scala 27:20]
  wire [21:0] _T_4258 = _T_2783 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4513 = _T_4512 | _T_4258; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_62; // @[Reg.scala 27:20]
  wire [21:0] _T_4259 = _T_2785 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4514 = _T_4513 | _T_4259; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_63; // @[Reg.scala 27:20]
  wire [21:0] _T_4260 = _T_2787 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4515 = _T_4514 | _T_4260; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_64; // @[Reg.scala 27:20]
  wire [21:0] _T_4261 = _T_2789 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4516 = _T_4515 | _T_4261; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_65; // @[Reg.scala 27:20]
  wire [21:0] _T_4262 = _T_2791 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4517 = _T_4516 | _T_4262; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_66; // @[Reg.scala 27:20]
  wire [21:0] _T_4263 = _T_2793 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4518 = _T_4517 | _T_4263; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_67; // @[Reg.scala 27:20]
  wire [21:0] _T_4264 = _T_2795 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4519 = _T_4518 | _T_4264; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_68; // @[Reg.scala 27:20]
  wire [21:0] _T_4265 = _T_2797 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4520 = _T_4519 | _T_4265; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_69; // @[Reg.scala 27:20]
  wire [21:0] _T_4266 = _T_2799 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4521 = _T_4520 | _T_4266; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_70; // @[Reg.scala 27:20]
  wire [21:0] _T_4267 = _T_2801 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4522 = _T_4521 | _T_4267; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_71; // @[Reg.scala 27:20]
  wire [21:0] _T_4268 = _T_2803 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4523 = _T_4522 | _T_4268; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_72; // @[Reg.scala 27:20]
  wire [21:0] _T_4269 = _T_2805 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4524 = _T_4523 | _T_4269; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_73; // @[Reg.scala 27:20]
  wire [21:0] _T_4270 = _T_2807 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4525 = _T_4524 | _T_4270; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_74; // @[Reg.scala 27:20]
  wire [21:0] _T_4271 = _T_2809 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4526 = _T_4525 | _T_4271; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_75; // @[Reg.scala 27:20]
  wire [21:0] _T_4272 = _T_2811 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4527 = _T_4526 | _T_4272; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_76; // @[Reg.scala 27:20]
  wire [21:0] _T_4273 = _T_2813 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4528 = _T_4527 | _T_4273; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_77; // @[Reg.scala 27:20]
  wire [21:0] _T_4274 = _T_2815 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4529 = _T_4528 | _T_4274; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_78; // @[Reg.scala 27:20]
  wire [21:0] _T_4275 = _T_2817 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4530 = _T_4529 | _T_4275; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_79; // @[Reg.scala 27:20]
  wire [21:0] _T_4276 = _T_2819 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4531 = _T_4530 | _T_4276; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_80; // @[Reg.scala 27:20]
  wire [21:0] _T_4277 = _T_2821 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4532 = _T_4531 | _T_4277; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_81; // @[Reg.scala 27:20]
  wire [21:0] _T_4278 = _T_2823 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4533 = _T_4532 | _T_4278; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_82; // @[Reg.scala 27:20]
  wire [21:0] _T_4279 = _T_2825 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4534 = _T_4533 | _T_4279; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_83; // @[Reg.scala 27:20]
  wire [21:0] _T_4280 = _T_2827 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4535 = _T_4534 | _T_4280; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_84; // @[Reg.scala 27:20]
  wire [21:0] _T_4281 = _T_2829 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4536 = _T_4535 | _T_4281; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_85; // @[Reg.scala 27:20]
  wire [21:0] _T_4282 = _T_2831 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4537 = _T_4536 | _T_4282; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_86; // @[Reg.scala 27:20]
  wire [21:0] _T_4283 = _T_2833 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4538 = _T_4537 | _T_4283; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_87; // @[Reg.scala 27:20]
  wire [21:0] _T_4284 = _T_2835 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4539 = _T_4538 | _T_4284; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_88; // @[Reg.scala 27:20]
  wire [21:0] _T_4285 = _T_2837 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4540 = _T_4539 | _T_4285; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_89; // @[Reg.scala 27:20]
  wire [21:0] _T_4286 = _T_2839 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4541 = _T_4540 | _T_4286; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_90; // @[Reg.scala 27:20]
  wire [21:0] _T_4287 = _T_2841 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4542 = _T_4541 | _T_4287; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_91; // @[Reg.scala 27:20]
  wire [21:0] _T_4288 = _T_2843 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4543 = _T_4542 | _T_4288; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_92; // @[Reg.scala 27:20]
  wire [21:0] _T_4289 = _T_2845 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4544 = _T_4543 | _T_4289; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_93; // @[Reg.scala 27:20]
  wire [21:0] _T_4290 = _T_2847 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4545 = _T_4544 | _T_4290; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_94; // @[Reg.scala 27:20]
  wire [21:0] _T_4291 = _T_2849 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4546 = _T_4545 | _T_4291; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_95; // @[Reg.scala 27:20]
  wire [21:0] _T_4292 = _T_2851 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4547 = _T_4546 | _T_4292; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_96; // @[Reg.scala 27:20]
  wire [21:0] _T_4293 = _T_2853 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4548 = _T_4547 | _T_4293; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_97; // @[Reg.scala 27:20]
  wire [21:0] _T_4294 = _T_2855 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4549 = _T_4548 | _T_4294; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_98; // @[Reg.scala 27:20]
  wire [21:0] _T_4295 = _T_2857 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4550 = _T_4549 | _T_4295; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_99; // @[Reg.scala 27:20]
  wire [21:0] _T_4296 = _T_2859 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4551 = _T_4550 | _T_4296; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_100; // @[Reg.scala 27:20]
  wire [21:0] _T_4297 = _T_2861 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4552 = _T_4551 | _T_4297; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_101; // @[Reg.scala 27:20]
  wire [21:0] _T_4298 = _T_2863 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4553 = _T_4552 | _T_4298; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_102; // @[Reg.scala 27:20]
  wire [21:0] _T_4299 = _T_2865 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4554 = _T_4553 | _T_4299; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_103; // @[Reg.scala 27:20]
  wire [21:0] _T_4300 = _T_2867 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4555 = _T_4554 | _T_4300; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_104; // @[Reg.scala 27:20]
  wire [21:0] _T_4301 = _T_2869 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4556 = _T_4555 | _T_4301; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_105; // @[Reg.scala 27:20]
  wire [21:0] _T_4302 = _T_2871 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4557 = _T_4556 | _T_4302; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_106; // @[Reg.scala 27:20]
  wire [21:0] _T_4303 = _T_2873 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4558 = _T_4557 | _T_4303; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_107; // @[Reg.scala 27:20]
  wire [21:0] _T_4304 = _T_2875 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4559 = _T_4558 | _T_4304; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_108; // @[Reg.scala 27:20]
  wire [21:0] _T_4305 = _T_2877 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4560 = _T_4559 | _T_4305; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_109; // @[Reg.scala 27:20]
  wire [21:0] _T_4306 = _T_2879 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4561 = _T_4560 | _T_4306; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_110; // @[Reg.scala 27:20]
  wire [21:0] _T_4307 = _T_2881 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4562 = _T_4561 | _T_4307; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_111; // @[Reg.scala 27:20]
  wire [21:0] _T_4308 = _T_2883 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4563 = _T_4562 | _T_4308; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_112; // @[Reg.scala 27:20]
  wire [21:0] _T_4309 = _T_2885 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4564 = _T_4563 | _T_4309; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_113; // @[Reg.scala 27:20]
  wire [21:0] _T_4310 = _T_2887 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4565 = _T_4564 | _T_4310; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_114; // @[Reg.scala 27:20]
  wire [21:0] _T_4311 = _T_2889 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4566 = _T_4565 | _T_4311; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_115; // @[Reg.scala 27:20]
  wire [21:0] _T_4312 = _T_2891 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4567 = _T_4566 | _T_4312; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_116; // @[Reg.scala 27:20]
  wire [21:0] _T_4313 = _T_2893 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4568 = _T_4567 | _T_4313; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_117; // @[Reg.scala 27:20]
  wire [21:0] _T_4314 = _T_2895 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4569 = _T_4568 | _T_4314; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_118; // @[Reg.scala 27:20]
  wire [21:0] _T_4315 = _T_2897 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4570 = _T_4569 | _T_4315; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_119; // @[Reg.scala 27:20]
  wire [21:0] _T_4316 = _T_2899 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4571 = _T_4570 | _T_4316; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_120; // @[Reg.scala 27:20]
  wire [21:0] _T_4317 = _T_2901 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4572 = _T_4571 | _T_4317; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_121; // @[Reg.scala 27:20]
  wire [21:0] _T_4318 = _T_2903 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4573 = _T_4572 | _T_4318; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_122; // @[Reg.scala 27:20]
  wire [21:0] _T_4319 = _T_2905 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4574 = _T_4573 | _T_4319; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_123; // @[Reg.scala 27:20]
  wire [21:0] _T_4320 = _T_2907 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4575 = _T_4574 | _T_4320; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_124; // @[Reg.scala 27:20]
  wire [21:0] _T_4321 = _T_2909 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4576 = _T_4575 | _T_4321; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_125; // @[Reg.scala 27:20]
  wire [21:0] _T_4322 = _T_2911 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4577 = _T_4576 | _T_4322; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_126; // @[Reg.scala 27:20]
  wire [21:0] _T_4323 = _T_2913 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4578 = _T_4577 | _T_4323; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_127; // @[Reg.scala 27:20]
  wire [21:0] _T_4324 = _T_2915 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4579 = _T_4578 | _T_4324; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_128; // @[Reg.scala 27:20]
  wire [21:0] _T_4325 = _T_2917 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4580 = _T_4579 | _T_4325; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_129; // @[Reg.scala 27:20]
  wire [21:0] _T_4326 = _T_2919 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4581 = _T_4580 | _T_4326; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_130; // @[Reg.scala 27:20]
  wire [21:0] _T_4327 = _T_2921 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4582 = _T_4581 | _T_4327; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_131; // @[Reg.scala 27:20]
  wire [21:0] _T_4328 = _T_2923 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4583 = _T_4582 | _T_4328; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_132; // @[Reg.scala 27:20]
  wire [21:0] _T_4329 = _T_2925 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4584 = _T_4583 | _T_4329; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_133; // @[Reg.scala 27:20]
  wire [21:0] _T_4330 = _T_2927 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4585 = _T_4584 | _T_4330; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_134; // @[Reg.scala 27:20]
  wire [21:0] _T_4331 = _T_2929 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4586 = _T_4585 | _T_4331; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_135; // @[Reg.scala 27:20]
  wire [21:0] _T_4332 = _T_2931 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4587 = _T_4586 | _T_4332; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_136; // @[Reg.scala 27:20]
  wire [21:0] _T_4333 = _T_2933 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4588 = _T_4587 | _T_4333; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_137; // @[Reg.scala 27:20]
  wire [21:0] _T_4334 = _T_2935 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4589 = _T_4588 | _T_4334; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_138; // @[Reg.scala 27:20]
  wire [21:0] _T_4335 = _T_2937 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4590 = _T_4589 | _T_4335; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_139; // @[Reg.scala 27:20]
  wire [21:0] _T_4336 = _T_2939 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4591 = _T_4590 | _T_4336; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_140; // @[Reg.scala 27:20]
  wire [21:0] _T_4337 = _T_2941 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4592 = _T_4591 | _T_4337; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_141; // @[Reg.scala 27:20]
  wire [21:0] _T_4338 = _T_2943 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4593 = _T_4592 | _T_4338; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_142; // @[Reg.scala 27:20]
  wire [21:0] _T_4339 = _T_2945 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4594 = _T_4593 | _T_4339; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_143; // @[Reg.scala 27:20]
  wire [21:0] _T_4340 = _T_2947 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4595 = _T_4594 | _T_4340; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_144; // @[Reg.scala 27:20]
  wire [21:0] _T_4341 = _T_2949 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4596 = _T_4595 | _T_4341; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_145; // @[Reg.scala 27:20]
  wire [21:0] _T_4342 = _T_2951 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4597 = _T_4596 | _T_4342; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_146; // @[Reg.scala 27:20]
  wire [21:0] _T_4343 = _T_2953 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4598 = _T_4597 | _T_4343; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_147; // @[Reg.scala 27:20]
  wire [21:0] _T_4344 = _T_2955 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4599 = _T_4598 | _T_4344; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_148; // @[Reg.scala 27:20]
  wire [21:0] _T_4345 = _T_2957 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4600 = _T_4599 | _T_4345; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_149; // @[Reg.scala 27:20]
  wire [21:0] _T_4346 = _T_2959 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4601 = _T_4600 | _T_4346; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_150; // @[Reg.scala 27:20]
  wire [21:0] _T_4347 = _T_2961 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4602 = _T_4601 | _T_4347; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_151; // @[Reg.scala 27:20]
  wire [21:0] _T_4348 = _T_2963 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4603 = _T_4602 | _T_4348; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_152; // @[Reg.scala 27:20]
  wire [21:0] _T_4349 = _T_2965 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4604 = _T_4603 | _T_4349; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_153; // @[Reg.scala 27:20]
  wire [21:0] _T_4350 = _T_2967 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4605 = _T_4604 | _T_4350; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_154; // @[Reg.scala 27:20]
  wire [21:0] _T_4351 = _T_2969 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4606 = _T_4605 | _T_4351; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_155; // @[Reg.scala 27:20]
  wire [21:0] _T_4352 = _T_2971 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4607 = _T_4606 | _T_4352; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_156; // @[Reg.scala 27:20]
  wire [21:0] _T_4353 = _T_2973 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4608 = _T_4607 | _T_4353; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_157; // @[Reg.scala 27:20]
  wire [21:0] _T_4354 = _T_2975 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4609 = _T_4608 | _T_4354; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_158; // @[Reg.scala 27:20]
  wire [21:0] _T_4355 = _T_2977 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4610 = _T_4609 | _T_4355; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_159; // @[Reg.scala 27:20]
  wire [21:0] _T_4356 = _T_2979 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4611 = _T_4610 | _T_4356; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_160; // @[Reg.scala 27:20]
  wire [21:0] _T_4357 = _T_2981 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4612 = _T_4611 | _T_4357; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_161; // @[Reg.scala 27:20]
  wire [21:0] _T_4358 = _T_2983 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4613 = _T_4612 | _T_4358; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_162; // @[Reg.scala 27:20]
  wire [21:0] _T_4359 = _T_2985 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4614 = _T_4613 | _T_4359; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_163; // @[Reg.scala 27:20]
  wire [21:0] _T_4360 = _T_2987 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4615 = _T_4614 | _T_4360; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_164; // @[Reg.scala 27:20]
  wire [21:0] _T_4361 = _T_2989 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4616 = _T_4615 | _T_4361; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_165; // @[Reg.scala 27:20]
  wire [21:0] _T_4362 = _T_2991 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4617 = _T_4616 | _T_4362; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_166; // @[Reg.scala 27:20]
  wire [21:0] _T_4363 = _T_2993 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4618 = _T_4617 | _T_4363; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_167; // @[Reg.scala 27:20]
  wire [21:0] _T_4364 = _T_2995 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4619 = _T_4618 | _T_4364; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_168; // @[Reg.scala 27:20]
  wire [21:0] _T_4365 = _T_2997 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4620 = _T_4619 | _T_4365; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_169; // @[Reg.scala 27:20]
  wire [21:0] _T_4366 = _T_2999 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4621 = _T_4620 | _T_4366; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_170; // @[Reg.scala 27:20]
  wire [21:0] _T_4367 = _T_3001 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4622 = _T_4621 | _T_4367; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_171; // @[Reg.scala 27:20]
  wire [21:0] _T_4368 = _T_3003 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4623 = _T_4622 | _T_4368; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_172; // @[Reg.scala 27:20]
  wire [21:0] _T_4369 = _T_3005 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4624 = _T_4623 | _T_4369; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_173; // @[Reg.scala 27:20]
  wire [21:0] _T_4370 = _T_3007 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4625 = _T_4624 | _T_4370; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_174; // @[Reg.scala 27:20]
  wire [21:0] _T_4371 = _T_3009 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4626 = _T_4625 | _T_4371; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_175; // @[Reg.scala 27:20]
  wire [21:0] _T_4372 = _T_3011 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4627 = _T_4626 | _T_4372; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_176; // @[Reg.scala 27:20]
  wire [21:0] _T_4373 = _T_3013 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4628 = _T_4627 | _T_4373; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_177; // @[Reg.scala 27:20]
  wire [21:0] _T_4374 = _T_3015 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4629 = _T_4628 | _T_4374; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_178; // @[Reg.scala 27:20]
  wire [21:0] _T_4375 = _T_3017 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4630 = _T_4629 | _T_4375; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_179; // @[Reg.scala 27:20]
  wire [21:0] _T_4376 = _T_3019 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4631 = _T_4630 | _T_4376; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_180; // @[Reg.scala 27:20]
  wire [21:0] _T_4377 = _T_3021 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4632 = _T_4631 | _T_4377; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_181; // @[Reg.scala 27:20]
  wire [21:0] _T_4378 = _T_3023 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4633 = _T_4632 | _T_4378; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_182; // @[Reg.scala 27:20]
  wire [21:0] _T_4379 = _T_3025 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4634 = _T_4633 | _T_4379; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_183; // @[Reg.scala 27:20]
  wire [21:0] _T_4380 = _T_3027 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4635 = _T_4634 | _T_4380; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_184; // @[Reg.scala 27:20]
  wire [21:0] _T_4381 = _T_3029 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4636 = _T_4635 | _T_4381; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_185; // @[Reg.scala 27:20]
  wire [21:0] _T_4382 = _T_3031 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4637 = _T_4636 | _T_4382; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_186; // @[Reg.scala 27:20]
  wire [21:0] _T_4383 = _T_3033 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4638 = _T_4637 | _T_4383; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_187; // @[Reg.scala 27:20]
  wire [21:0] _T_4384 = _T_3035 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4639 = _T_4638 | _T_4384; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_188; // @[Reg.scala 27:20]
  wire [21:0] _T_4385 = _T_3037 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4640 = _T_4639 | _T_4385; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_189; // @[Reg.scala 27:20]
  wire [21:0] _T_4386 = _T_3039 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4641 = _T_4640 | _T_4386; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_190; // @[Reg.scala 27:20]
  wire [21:0] _T_4387 = _T_3041 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4642 = _T_4641 | _T_4387; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_191; // @[Reg.scala 27:20]
  wire [21:0] _T_4388 = _T_3043 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4643 = _T_4642 | _T_4388; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_192; // @[Reg.scala 27:20]
  wire [21:0] _T_4389 = _T_3045 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4644 = _T_4643 | _T_4389; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_193; // @[Reg.scala 27:20]
  wire [21:0] _T_4390 = _T_3047 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4645 = _T_4644 | _T_4390; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_194; // @[Reg.scala 27:20]
  wire [21:0] _T_4391 = _T_3049 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4646 = _T_4645 | _T_4391; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_195; // @[Reg.scala 27:20]
  wire [21:0] _T_4392 = _T_3051 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4647 = _T_4646 | _T_4392; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_196; // @[Reg.scala 27:20]
  wire [21:0] _T_4393 = _T_3053 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4648 = _T_4647 | _T_4393; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_197; // @[Reg.scala 27:20]
  wire [21:0] _T_4394 = _T_3055 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4649 = _T_4648 | _T_4394; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_198; // @[Reg.scala 27:20]
  wire [21:0] _T_4395 = _T_3057 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4650 = _T_4649 | _T_4395; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_199; // @[Reg.scala 27:20]
  wire [21:0] _T_4396 = _T_3059 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4651 = _T_4650 | _T_4396; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_200; // @[Reg.scala 27:20]
  wire [21:0] _T_4397 = _T_3061 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4652 = _T_4651 | _T_4397; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_201; // @[Reg.scala 27:20]
  wire [21:0] _T_4398 = _T_3063 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4653 = _T_4652 | _T_4398; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_202; // @[Reg.scala 27:20]
  wire [21:0] _T_4399 = _T_3065 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4654 = _T_4653 | _T_4399; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_203; // @[Reg.scala 27:20]
  wire [21:0] _T_4400 = _T_3067 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4655 = _T_4654 | _T_4400; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_204; // @[Reg.scala 27:20]
  wire [21:0] _T_4401 = _T_3069 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4656 = _T_4655 | _T_4401; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_205; // @[Reg.scala 27:20]
  wire [21:0] _T_4402 = _T_3071 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4657 = _T_4656 | _T_4402; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_206; // @[Reg.scala 27:20]
  wire [21:0] _T_4403 = _T_3073 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4658 = _T_4657 | _T_4403; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_207; // @[Reg.scala 27:20]
  wire [21:0] _T_4404 = _T_3075 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4659 = _T_4658 | _T_4404; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_208; // @[Reg.scala 27:20]
  wire [21:0] _T_4405 = _T_3077 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4660 = _T_4659 | _T_4405; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_209; // @[Reg.scala 27:20]
  wire [21:0] _T_4406 = _T_3079 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4661 = _T_4660 | _T_4406; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_210; // @[Reg.scala 27:20]
  wire [21:0] _T_4407 = _T_3081 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4662 = _T_4661 | _T_4407; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_211; // @[Reg.scala 27:20]
  wire [21:0] _T_4408 = _T_3083 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4663 = _T_4662 | _T_4408; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_212; // @[Reg.scala 27:20]
  wire [21:0] _T_4409 = _T_3085 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4664 = _T_4663 | _T_4409; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_213; // @[Reg.scala 27:20]
  wire [21:0] _T_4410 = _T_3087 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4665 = _T_4664 | _T_4410; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_214; // @[Reg.scala 27:20]
  wire [21:0] _T_4411 = _T_3089 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4666 = _T_4665 | _T_4411; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_215; // @[Reg.scala 27:20]
  wire [21:0] _T_4412 = _T_3091 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4667 = _T_4666 | _T_4412; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_216; // @[Reg.scala 27:20]
  wire [21:0] _T_4413 = _T_3093 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4668 = _T_4667 | _T_4413; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_217; // @[Reg.scala 27:20]
  wire [21:0] _T_4414 = _T_3095 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4669 = _T_4668 | _T_4414; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_218; // @[Reg.scala 27:20]
  wire [21:0] _T_4415 = _T_3097 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4670 = _T_4669 | _T_4415; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_219; // @[Reg.scala 27:20]
  wire [21:0] _T_4416 = _T_3099 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4671 = _T_4670 | _T_4416; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_220; // @[Reg.scala 27:20]
  wire [21:0] _T_4417 = _T_3101 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4672 = _T_4671 | _T_4417; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_221; // @[Reg.scala 27:20]
  wire [21:0] _T_4418 = _T_3103 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4673 = _T_4672 | _T_4418; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_222; // @[Reg.scala 27:20]
  wire [21:0] _T_4419 = _T_3105 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4674 = _T_4673 | _T_4419; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_223; // @[Reg.scala 27:20]
  wire [21:0] _T_4420 = _T_3107 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4675 = _T_4674 | _T_4420; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_224; // @[Reg.scala 27:20]
  wire [21:0] _T_4421 = _T_3109 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4676 = _T_4675 | _T_4421; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_225; // @[Reg.scala 27:20]
  wire [21:0] _T_4422 = _T_3111 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4677 = _T_4676 | _T_4422; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_226; // @[Reg.scala 27:20]
  wire [21:0] _T_4423 = _T_3113 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4678 = _T_4677 | _T_4423; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_227; // @[Reg.scala 27:20]
  wire [21:0] _T_4424 = _T_3115 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4679 = _T_4678 | _T_4424; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_228; // @[Reg.scala 27:20]
  wire [21:0] _T_4425 = _T_3117 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4680 = _T_4679 | _T_4425; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_229; // @[Reg.scala 27:20]
  wire [21:0] _T_4426 = _T_3119 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4681 = _T_4680 | _T_4426; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_230; // @[Reg.scala 27:20]
  wire [21:0] _T_4427 = _T_3121 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4682 = _T_4681 | _T_4427; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_231; // @[Reg.scala 27:20]
  wire [21:0] _T_4428 = _T_3123 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4683 = _T_4682 | _T_4428; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_232; // @[Reg.scala 27:20]
  wire [21:0] _T_4429 = _T_3125 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4684 = _T_4683 | _T_4429; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_233; // @[Reg.scala 27:20]
  wire [21:0] _T_4430 = _T_3127 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4685 = _T_4684 | _T_4430; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_234; // @[Reg.scala 27:20]
  wire [21:0] _T_4431 = _T_3129 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4686 = _T_4685 | _T_4431; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_235; // @[Reg.scala 27:20]
  wire [21:0] _T_4432 = _T_3131 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4687 = _T_4686 | _T_4432; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_236; // @[Reg.scala 27:20]
  wire [21:0] _T_4433 = _T_3133 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4688 = _T_4687 | _T_4433; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_237; // @[Reg.scala 27:20]
  wire [21:0] _T_4434 = _T_3135 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4689 = _T_4688 | _T_4434; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_238; // @[Reg.scala 27:20]
  wire [21:0] _T_4435 = _T_3137 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4690 = _T_4689 | _T_4435; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_239; // @[Reg.scala 27:20]
  wire [21:0] _T_4436 = _T_3139 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4691 = _T_4690 | _T_4436; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_240; // @[Reg.scala 27:20]
  wire [21:0] _T_4437 = _T_3141 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4692 = _T_4691 | _T_4437; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_241; // @[Reg.scala 27:20]
  wire [21:0] _T_4438 = _T_3143 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4693 = _T_4692 | _T_4438; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_242; // @[Reg.scala 27:20]
  wire [21:0] _T_4439 = _T_3145 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4694 = _T_4693 | _T_4439; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_243; // @[Reg.scala 27:20]
  wire [21:0] _T_4440 = _T_3147 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4695 = _T_4694 | _T_4440; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_244; // @[Reg.scala 27:20]
  wire [21:0] _T_4441 = _T_3149 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4696 = _T_4695 | _T_4441; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_245; // @[Reg.scala 27:20]
  wire [21:0] _T_4442 = _T_3151 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4697 = _T_4696 | _T_4442; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_246; // @[Reg.scala 27:20]
  wire [21:0] _T_4443 = _T_3153 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4698 = _T_4697 | _T_4443; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_247; // @[Reg.scala 27:20]
  wire [21:0] _T_4444 = _T_3155 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4699 = _T_4698 | _T_4444; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_248; // @[Reg.scala 27:20]
  wire [21:0] _T_4445 = _T_3157 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4700 = _T_4699 | _T_4445; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_249; // @[Reg.scala 27:20]
  wire [21:0] _T_4446 = _T_3159 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4701 = _T_4700 | _T_4446; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_250; // @[Reg.scala 27:20]
  wire [21:0] _T_4447 = _T_3161 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4702 = _T_4701 | _T_4447; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_251; // @[Reg.scala 27:20]
  wire [21:0] _T_4448 = _T_3163 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4703 = _T_4702 | _T_4448; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_252; // @[Reg.scala 27:20]
  wire [21:0] _T_4449 = _T_3165 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4704 = _T_4703 | _T_4449; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_253; // @[Reg.scala 27:20]
  wire [21:0] _T_4450 = _T_3167 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4705 = _T_4704 | _T_4450; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_254; // @[Reg.scala 27:20]
  wire [21:0] _T_4451 = _T_3169 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_4706 = _T_4705 | _T_4451; // @[Mux.scala 27:72]
  reg [21:0] btb_bank0_rd_data_way1_out_255; // @[Reg.scala 27:20]
  wire [21:0] _T_4452 = _T_3171 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_f = _T_4706 | _T_4452; // @[Mux.scala 27:72]
  wire  _T_55 = btb_bank0_rd_data_way1_f[21:17] == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 148:98]
  wire  _T_56 = btb_bank0_rd_data_way1_f[0] & _T_55; // @[ifu_bp_ctl.scala 148:55]
  wire  _T_59 = _T_56 & _T_49; // @[ifu_bp_ctl.scala 148:118]
  wire  _T_60 = _T_59 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 149:54]
  wire  tag_match_way1_f = _T_60 & _T; // @[ifu_bp_ctl.scala 149:75]
  wire  _T_91 = btb_bank0_rd_data_way1_f[3] ^ btb_bank0_rd_data_way1_f[4]; // @[ifu_bp_ctl.scala 162:90]
  wire  _T_92 = tag_match_way1_f & _T_91; // @[ifu_bp_ctl.scala 162:56]
  wire  _T_96 = ~_T_91; // @[ifu_bp_ctl.scala 163:24]
  wire  _T_97 = tag_match_way1_f & _T_96; // @[ifu_bp_ctl.scala 163:22]
  wire [1:0] tag_match_way1_expanded_f = {_T_92,_T_97}; // @[Cat.scala 29:58]
  wire [21:0] _T_130 = tag_match_way1_expanded_f[1] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0o_rd_data_f = _T_129 | _T_130; // @[Mux.scala 27:72]
  wire [21:0] _T_149 = _T_147 ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4709 = btb_rd_addr_p1_f == 8'h0; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5221 = _T_4709 ? btb_bank0_rd_data_way0_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire  _T_4711 = btb_rd_addr_p1_f == 8'h1; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5222 = _T_4711 ? btb_bank0_rd_data_way0_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5477 = _T_5221 | _T_5222; // @[Mux.scala 27:72]
  wire  _T_4713 = btb_rd_addr_p1_f == 8'h2; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5223 = _T_4713 ? btb_bank0_rd_data_way0_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5478 = _T_5477 | _T_5223; // @[Mux.scala 27:72]
  wire  _T_4715 = btb_rd_addr_p1_f == 8'h3; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5224 = _T_4715 ? btb_bank0_rd_data_way0_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5479 = _T_5478 | _T_5224; // @[Mux.scala 27:72]
  wire  _T_4717 = btb_rd_addr_p1_f == 8'h4; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5225 = _T_4717 ? btb_bank0_rd_data_way0_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5480 = _T_5479 | _T_5225; // @[Mux.scala 27:72]
  wire  _T_4719 = btb_rd_addr_p1_f == 8'h5; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5226 = _T_4719 ? btb_bank0_rd_data_way0_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5481 = _T_5480 | _T_5226; // @[Mux.scala 27:72]
  wire  _T_4721 = btb_rd_addr_p1_f == 8'h6; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5227 = _T_4721 ? btb_bank0_rd_data_way0_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5482 = _T_5481 | _T_5227; // @[Mux.scala 27:72]
  wire  _T_4723 = btb_rd_addr_p1_f == 8'h7; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5228 = _T_4723 ? btb_bank0_rd_data_way0_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5483 = _T_5482 | _T_5228; // @[Mux.scala 27:72]
  wire  _T_4725 = btb_rd_addr_p1_f == 8'h8; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5229 = _T_4725 ? btb_bank0_rd_data_way0_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5484 = _T_5483 | _T_5229; // @[Mux.scala 27:72]
  wire  _T_4727 = btb_rd_addr_p1_f == 8'h9; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5230 = _T_4727 ? btb_bank0_rd_data_way0_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5485 = _T_5484 | _T_5230; // @[Mux.scala 27:72]
  wire  _T_4729 = btb_rd_addr_p1_f == 8'ha; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5231 = _T_4729 ? btb_bank0_rd_data_way0_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5486 = _T_5485 | _T_5231; // @[Mux.scala 27:72]
  wire  _T_4731 = btb_rd_addr_p1_f == 8'hb; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5232 = _T_4731 ? btb_bank0_rd_data_way0_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5487 = _T_5486 | _T_5232; // @[Mux.scala 27:72]
  wire  _T_4733 = btb_rd_addr_p1_f == 8'hc; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5233 = _T_4733 ? btb_bank0_rd_data_way0_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5488 = _T_5487 | _T_5233; // @[Mux.scala 27:72]
  wire  _T_4735 = btb_rd_addr_p1_f == 8'hd; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5234 = _T_4735 ? btb_bank0_rd_data_way0_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5489 = _T_5488 | _T_5234; // @[Mux.scala 27:72]
  wire  _T_4737 = btb_rd_addr_p1_f == 8'he; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5235 = _T_4737 ? btb_bank0_rd_data_way0_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5490 = _T_5489 | _T_5235; // @[Mux.scala 27:72]
  wire  _T_4739 = btb_rd_addr_p1_f == 8'hf; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5236 = _T_4739 ? btb_bank0_rd_data_way0_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5491 = _T_5490 | _T_5236; // @[Mux.scala 27:72]
  wire  _T_4741 = btb_rd_addr_p1_f == 8'h10; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5237 = _T_4741 ? btb_bank0_rd_data_way0_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5492 = _T_5491 | _T_5237; // @[Mux.scala 27:72]
  wire  _T_4743 = btb_rd_addr_p1_f == 8'h11; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5238 = _T_4743 ? btb_bank0_rd_data_way0_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5493 = _T_5492 | _T_5238; // @[Mux.scala 27:72]
  wire  _T_4745 = btb_rd_addr_p1_f == 8'h12; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5239 = _T_4745 ? btb_bank0_rd_data_way0_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5494 = _T_5493 | _T_5239; // @[Mux.scala 27:72]
  wire  _T_4747 = btb_rd_addr_p1_f == 8'h13; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5240 = _T_4747 ? btb_bank0_rd_data_way0_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5495 = _T_5494 | _T_5240; // @[Mux.scala 27:72]
  wire  _T_4749 = btb_rd_addr_p1_f == 8'h14; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5241 = _T_4749 ? btb_bank0_rd_data_way0_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5496 = _T_5495 | _T_5241; // @[Mux.scala 27:72]
  wire  _T_4751 = btb_rd_addr_p1_f == 8'h15; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5242 = _T_4751 ? btb_bank0_rd_data_way0_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5497 = _T_5496 | _T_5242; // @[Mux.scala 27:72]
  wire  _T_4753 = btb_rd_addr_p1_f == 8'h16; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5243 = _T_4753 ? btb_bank0_rd_data_way0_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5498 = _T_5497 | _T_5243; // @[Mux.scala 27:72]
  wire  _T_4755 = btb_rd_addr_p1_f == 8'h17; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5244 = _T_4755 ? btb_bank0_rd_data_way0_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5499 = _T_5498 | _T_5244; // @[Mux.scala 27:72]
  wire  _T_4757 = btb_rd_addr_p1_f == 8'h18; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5245 = _T_4757 ? btb_bank0_rd_data_way0_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5500 = _T_5499 | _T_5245; // @[Mux.scala 27:72]
  wire  _T_4759 = btb_rd_addr_p1_f == 8'h19; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5246 = _T_4759 ? btb_bank0_rd_data_way0_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5501 = _T_5500 | _T_5246; // @[Mux.scala 27:72]
  wire  _T_4761 = btb_rd_addr_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5247 = _T_4761 ? btb_bank0_rd_data_way0_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5502 = _T_5501 | _T_5247; // @[Mux.scala 27:72]
  wire  _T_4763 = btb_rd_addr_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5248 = _T_4763 ? btb_bank0_rd_data_way0_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5503 = _T_5502 | _T_5248; // @[Mux.scala 27:72]
  wire  _T_4765 = btb_rd_addr_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5249 = _T_4765 ? btb_bank0_rd_data_way0_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5504 = _T_5503 | _T_5249; // @[Mux.scala 27:72]
  wire  _T_4767 = btb_rd_addr_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5250 = _T_4767 ? btb_bank0_rd_data_way0_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5505 = _T_5504 | _T_5250; // @[Mux.scala 27:72]
  wire  _T_4769 = btb_rd_addr_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5251 = _T_4769 ? btb_bank0_rd_data_way0_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5506 = _T_5505 | _T_5251; // @[Mux.scala 27:72]
  wire  _T_4771 = btb_rd_addr_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5252 = _T_4771 ? btb_bank0_rd_data_way0_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5507 = _T_5506 | _T_5252; // @[Mux.scala 27:72]
  wire  _T_4773 = btb_rd_addr_p1_f == 8'h20; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5253 = _T_4773 ? btb_bank0_rd_data_way0_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5508 = _T_5507 | _T_5253; // @[Mux.scala 27:72]
  wire  _T_4775 = btb_rd_addr_p1_f == 8'h21; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5254 = _T_4775 ? btb_bank0_rd_data_way0_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5509 = _T_5508 | _T_5254; // @[Mux.scala 27:72]
  wire  _T_4777 = btb_rd_addr_p1_f == 8'h22; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5255 = _T_4777 ? btb_bank0_rd_data_way0_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5510 = _T_5509 | _T_5255; // @[Mux.scala 27:72]
  wire  _T_4779 = btb_rd_addr_p1_f == 8'h23; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5256 = _T_4779 ? btb_bank0_rd_data_way0_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5511 = _T_5510 | _T_5256; // @[Mux.scala 27:72]
  wire  _T_4781 = btb_rd_addr_p1_f == 8'h24; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5257 = _T_4781 ? btb_bank0_rd_data_way0_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5512 = _T_5511 | _T_5257; // @[Mux.scala 27:72]
  wire  _T_4783 = btb_rd_addr_p1_f == 8'h25; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5258 = _T_4783 ? btb_bank0_rd_data_way0_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5513 = _T_5512 | _T_5258; // @[Mux.scala 27:72]
  wire  _T_4785 = btb_rd_addr_p1_f == 8'h26; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5259 = _T_4785 ? btb_bank0_rd_data_way0_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5514 = _T_5513 | _T_5259; // @[Mux.scala 27:72]
  wire  _T_4787 = btb_rd_addr_p1_f == 8'h27; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5260 = _T_4787 ? btb_bank0_rd_data_way0_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5515 = _T_5514 | _T_5260; // @[Mux.scala 27:72]
  wire  _T_4789 = btb_rd_addr_p1_f == 8'h28; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5261 = _T_4789 ? btb_bank0_rd_data_way0_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5516 = _T_5515 | _T_5261; // @[Mux.scala 27:72]
  wire  _T_4791 = btb_rd_addr_p1_f == 8'h29; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5262 = _T_4791 ? btb_bank0_rd_data_way0_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5517 = _T_5516 | _T_5262; // @[Mux.scala 27:72]
  wire  _T_4793 = btb_rd_addr_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5263 = _T_4793 ? btb_bank0_rd_data_way0_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5518 = _T_5517 | _T_5263; // @[Mux.scala 27:72]
  wire  _T_4795 = btb_rd_addr_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5264 = _T_4795 ? btb_bank0_rd_data_way0_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5519 = _T_5518 | _T_5264; // @[Mux.scala 27:72]
  wire  _T_4797 = btb_rd_addr_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5265 = _T_4797 ? btb_bank0_rd_data_way0_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5520 = _T_5519 | _T_5265; // @[Mux.scala 27:72]
  wire  _T_4799 = btb_rd_addr_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5266 = _T_4799 ? btb_bank0_rd_data_way0_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5521 = _T_5520 | _T_5266; // @[Mux.scala 27:72]
  wire  _T_4801 = btb_rd_addr_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5267 = _T_4801 ? btb_bank0_rd_data_way0_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5522 = _T_5521 | _T_5267; // @[Mux.scala 27:72]
  wire  _T_4803 = btb_rd_addr_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5268 = _T_4803 ? btb_bank0_rd_data_way0_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5523 = _T_5522 | _T_5268; // @[Mux.scala 27:72]
  wire  _T_4805 = btb_rd_addr_p1_f == 8'h30; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5269 = _T_4805 ? btb_bank0_rd_data_way0_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5524 = _T_5523 | _T_5269; // @[Mux.scala 27:72]
  wire  _T_4807 = btb_rd_addr_p1_f == 8'h31; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5270 = _T_4807 ? btb_bank0_rd_data_way0_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5525 = _T_5524 | _T_5270; // @[Mux.scala 27:72]
  wire  _T_4809 = btb_rd_addr_p1_f == 8'h32; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5271 = _T_4809 ? btb_bank0_rd_data_way0_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5526 = _T_5525 | _T_5271; // @[Mux.scala 27:72]
  wire  _T_4811 = btb_rd_addr_p1_f == 8'h33; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5272 = _T_4811 ? btb_bank0_rd_data_way0_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5527 = _T_5526 | _T_5272; // @[Mux.scala 27:72]
  wire  _T_4813 = btb_rd_addr_p1_f == 8'h34; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5273 = _T_4813 ? btb_bank0_rd_data_way0_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5528 = _T_5527 | _T_5273; // @[Mux.scala 27:72]
  wire  _T_4815 = btb_rd_addr_p1_f == 8'h35; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5274 = _T_4815 ? btb_bank0_rd_data_way0_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5529 = _T_5528 | _T_5274; // @[Mux.scala 27:72]
  wire  _T_4817 = btb_rd_addr_p1_f == 8'h36; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5275 = _T_4817 ? btb_bank0_rd_data_way0_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5530 = _T_5529 | _T_5275; // @[Mux.scala 27:72]
  wire  _T_4819 = btb_rd_addr_p1_f == 8'h37; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5276 = _T_4819 ? btb_bank0_rd_data_way0_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5531 = _T_5530 | _T_5276; // @[Mux.scala 27:72]
  wire  _T_4821 = btb_rd_addr_p1_f == 8'h38; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5277 = _T_4821 ? btb_bank0_rd_data_way0_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5532 = _T_5531 | _T_5277; // @[Mux.scala 27:72]
  wire  _T_4823 = btb_rd_addr_p1_f == 8'h39; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5278 = _T_4823 ? btb_bank0_rd_data_way0_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5533 = _T_5532 | _T_5278; // @[Mux.scala 27:72]
  wire  _T_4825 = btb_rd_addr_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5279 = _T_4825 ? btb_bank0_rd_data_way0_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5534 = _T_5533 | _T_5279; // @[Mux.scala 27:72]
  wire  _T_4827 = btb_rd_addr_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5280 = _T_4827 ? btb_bank0_rd_data_way0_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5535 = _T_5534 | _T_5280; // @[Mux.scala 27:72]
  wire  _T_4829 = btb_rd_addr_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5281 = _T_4829 ? btb_bank0_rd_data_way0_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5536 = _T_5535 | _T_5281; // @[Mux.scala 27:72]
  wire  _T_4831 = btb_rd_addr_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5282 = _T_4831 ? btb_bank0_rd_data_way0_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5537 = _T_5536 | _T_5282; // @[Mux.scala 27:72]
  wire  _T_4833 = btb_rd_addr_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5283 = _T_4833 ? btb_bank0_rd_data_way0_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5538 = _T_5537 | _T_5283; // @[Mux.scala 27:72]
  wire  _T_4835 = btb_rd_addr_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5284 = _T_4835 ? btb_bank0_rd_data_way0_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5539 = _T_5538 | _T_5284; // @[Mux.scala 27:72]
  wire  _T_4837 = btb_rd_addr_p1_f == 8'h40; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5285 = _T_4837 ? btb_bank0_rd_data_way0_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5540 = _T_5539 | _T_5285; // @[Mux.scala 27:72]
  wire  _T_4839 = btb_rd_addr_p1_f == 8'h41; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5286 = _T_4839 ? btb_bank0_rd_data_way0_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5541 = _T_5540 | _T_5286; // @[Mux.scala 27:72]
  wire  _T_4841 = btb_rd_addr_p1_f == 8'h42; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5287 = _T_4841 ? btb_bank0_rd_data_way0_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5542 = _T_5541 | _T_5287; // @[Mux.scala 27:72]
  wire  _T_4843 = btb_rd_addr_p1_f == 8'h43; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5288 = _T_4843 ? btb_bank0_rd_data_way0_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5543 = _T_5542 | _T_5288; // @[Mux.scala 27:72]
  wire  _T_4845 = btb_rd_addr_p1_f == 8'h44; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5289 = _T_4845 ? btb_bank0_rd_data_way0_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5544 = _T_5543 | _T_5289; // @[Mux.scala 27:72]
  wire  _T_4847 = btb_rd_addr_p1_f == 8'h45; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5290 = _T_4847 ? btb_bank0_rd_data_way0_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5545 = _T_5544 | _T_5290; // @[Mux.scala 27:72]
  wire  _T_4849 = btb_rd_addr_p1_f == 8'h46; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5291 = _T_4849 ? btb_bank0_rd_data_way0_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5546 = _T_5545 | _T_5291; // @[Mux.scala 27:72]
  wire  _T_4851 = btb_rd_addr_p1_f == 8'h47; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5292 = _T_4851 ? btb_bank0_rd_data_way0_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5547 = _T_5546 | _T_5292; // @[Mux.scala 27:72]
  wire  _T_4853 = btb_rd_addr_p1_f == 8'h48; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5293 = _T_4853 ? btb_bank0_rd_data_way0_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5548 = _T_5547 | _T_5293; // @[Mux.scala 27:72]
  wire  _T_4855 = btb_rd_addr_p1_f == 8'h49; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5294 = _T_4855 ? btb_bank0_rd_data_way0_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5549 = _T_5548 | _T_5294; // @[Mux.scala 27:72]
  wire  _T_4857 = btb_rd_addr_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5295 = _T_4857 ? btb_bank0_rd_data_way0_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5550 = _T_5549 | _T_5295; // @[Mux.scala 27:72]
  wire  _T_4859 = btb_rd_addr_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5296 = _T_4859 ? btb_bank0_rd_data_way0_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5551 = _T_5550 | _T_5296; // @[Mux.scala 27:72]
  wire  _T_4861 = btb_rd_addr_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5297 = _T_4861 ? btb_bank0_rd_data_way0_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5552 = _T_5551 | _T_5297; // @[Mux.scala 27:72]
  wire  _T_4863 = btb_rd_addr_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5298 = _T_4863 ? btb_bank0_rd_data_way0_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5553 = _T_5552 | _T_5298; // @[Mux.scala 27:72]
  wire  _T_4865 = btb_rd_addr_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5299 = _T_4865 ? btb_bank0_rd_data_way0_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5554 = _T_5553 | _T_5299; // @[Mux.scala 27:72]
  wire  _T_4867 = btb_rd_addr_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5300 = _T_4867 ? btb_bank0_rd_data_way0_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5555 = _T_5554 | _T_5300; // @[Mux.scala 27:72]
  wire  _T_4869 = btb_rd_addr_p1_f == 8'h50; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5301 = _T_4869 ? btb_bank0_rd_data_way0_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5556 = _T_5555 | _T_5301; // @[Mux.scala 27:72]
  wire  _T_4871 = btb_rd_addr_p1_f == 8'h51; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5302 = _T_4871 ? btb_bank0_rd_data_way0_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5557 = _T_5556 | _T_5302; // @[Mux.scala 27:72]
  wire  _T_4873 = btb_rd_addr_p1_f == 8'h52; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5303 = _T_4873 ? btb_bank0_rd_data_way0_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5558 = _T_5557 | _T_5303; // @[Mux.scala 27:72]
  wire  _T_4875 = btb_rd_addr_p1_f == 8'h53; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5304 = _T_4875 ? btb_bank0_rd_data_way0_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5559 = _T_5558 | _T_5304; // @[Mux.scala 27:72]
  wire  _T_4877 = btb_rd_addr_p1_f == 8'h54; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5305 = _T_4877 ? btb_bank0_rd_data_way0_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5560 = _T_5559 | _T_5305; // @[Mux.scala 27:72]
  wire  _T_4879 = btb_rd_addr_p1_f == 8'h55; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5306 = _T_4879 ? btb_bank0_rd_data_way0_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5561 = _T_5560 | _T_5306; // @[Mux.scala 27:72]
  wire  _T_4881 = btb_rd_addr_p1_f == 8'h56; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5307 = _T_4881 ? btb_bank0_rd_data_way0_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5562 = _T_5561 | _T_5307; // @[Mux.scala 27:72]
  wire  _T_4883 = btb_rd_addr_p1_f == 8'h57; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5308 = _T_4883 ? btb_bank0_rd_data_way0_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5563 = _T_5562 | _T_5308; // @[Mux.scala 27:72]
  wire  _T_4885 = btb_rd_addr_p1_f == 8'h58; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5309 = _T_4885 ? btb_bank0_rd_data_way0_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5564 = _T_5563 | _T_5309; // @[Mux.scala 27:72]
  wire  _T_4887 = btb_rd_addr_p1_f == 8'h59; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5310 = _T_4887 ? btb_bank0_rd_data_way0_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5565 = _T_5564 | _T_5310; // @[Mux.scala 27:72]
  wire  _T_4889 = btb_rd_addr_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5311 = _T_4889 ? btb_bank0_rd_data_way0_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5566 = _T_5565 | _T_5311; // @[Mux.scala 27:72]
  wire  _T_4891 = btb_rd_addr_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5312 = _T_4891 ? btb_bank0_rd_data_way0_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5567 = _T_5566 | _T_5312; // @[Mux.scala 27:72]
  wire  _T_4893 = btb_rd_addr_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5313 = _T_4893 ? btb_bank0_rd_data_way0_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5568 = _T_5567 | _T_5313; // @[Mux.scala 27:72]
  wire  _T_4895 = btb_rd_addr_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5314 = _T_4895 ? btb_bank0_rd_data_way0_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5569 = _T_5568 | _T_5314; // @[Mux.scala 27:72]
  wire  _T_4897 = btb_rd_addr_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5315 = _T_4897 ? btb_bank0_rd_data_way0_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5570 = _T_5569 | _T_5315; // @[Mux.scala 27:72]
  wire  _T_4899 = btb_rd_addr_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5316 = _T_4899 ? btb_bank0_rd_data_way0_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5571 = _T_5570 | _T_5316; // @[Mux.scala 27:72]
  wire  _T_4901 = btb_rd_addr_p1_f == 8'h60; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5317 = _T_4901 ? btb_bank0_rd_data_way0_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5572 = _T_5571 | _T_5317; // @[Mux.scala 27:72]
  wire  _T_4903 = btb_rd_addr_p1_f == 8'h61; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5318 = _T_4903 ? btb_bank0_rd_data_way0_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5573 = _T_5572 | _T_5318; // @[Mux.scala 27:72]
  wire  _T_4905 = btb_rd_addr_p1_f == 8'h62; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5319 = _T_4905 ? btb_bank0_rd_data_way0_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5574 = _T_5573 | _T_5319; // @[Mux.scala 27:72]
  wire  _T_4907 = btb_rd_addr_p1_f == 8'h63; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5320 = _T_4907 ? btb_bank0_rd_data_way0_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5575 = _T_5574 | _T_5320; // @[Mux.scala 27:72]
  wire  _T_4909 = btb_rd_addr_p1_f == 8'h64; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5321 = _T_4909 ? btb_bank0_rd_data_way0_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5576 = _T_5575 | _T_5321; // @[Mux.scala 27:72]
  wire  _T_4911 = btb_rd_addr_p1_f == 8'h65; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5322 = _T_4911 ? btb_bank0_rd_data_way0_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5577 = _T_5576 | _T_5322; // @[Mux.scala 27:72]
  wire  _T_4913 = btb_rd_addr_p1_f == 8'h66; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5323 = _T_4913 ? btb_bank0_rd_data_way0_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5578 = _T_5577 | _T_5323; // @[Mux.scala 27:72]
  wire  _T_4915 = btb_rd_addr_p1_f == 8'h67; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5324 = _T_4915 ? btb_bank0_rd_data_way0_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5579 = _T_5578 | _T_5324; // @[Mux.scala 27:72]
  wire  _T_4917 = btb_rd_addr_p1_f == 8'h68; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5325 = _T_4917 ? btb_bank0_rd_data_way0_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5580 = _T_5579 | _T_5325; // @[Mux.scala 27:72]
  wire  _T_4919 = btb_rd_addr_p1_f == 8'h69; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5326 = _T_4919 ? btb_bank0_rd_data_way0_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5581 = _T_5580 | _T_5326; // @[Mux.scala 27:72]
  wire  _T_4921 = btb_rd_addr_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5327 = _T_4921 ? btb_bank0_rd_data_way0_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5582 = _T_5581 | _T_5327; // @[Mux.scala 27:72]
  wire  _T_4923 = btb_rd_addr_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5328 = _T_4923 ? btb_bank0_rd_data_way0_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5583 = _T_5582 | _T_5328; // @[Mux.scala 27:72]
  wire  _T_4925 = btb_rd_addr_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5329 = _T_4925 ? btb_bank0_rd_data_way0_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5584 = _T_5583 | _T_5329; // @[Mux.scala 27:72]
  wire  _T_4927 = btb_rd_addr_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5330 = _T_4927 ? btb_bank0_rd_data_way0_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5585 = _T_5584 | _T_5330; // @[Mux.scala 27:72]
  wire  _T_4929 = btb_rd_addr_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5331 = _T_4929 ? btb_bank0_rd_data_way0_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5586 = _T_5585 | _T_5331; // @[Mux.scala 27:72]
  wire  _T_4931 = btb_rd_addr_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5332 = _T_4931 ? btb_bank0_rd_data_way0_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5587 = _T_5586 | _T_5332; // @[Mux.scala 27:72]
  wire  _T_4933 = btb_rd_addr_p1_f == 8'h70; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5333 = _T_4933 ? btb_bank0_rd_data_way0_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5588 = _T_5587 | _T_5333; // @[Mux.scala 27:72]
  wire  _T_4935 = btb_rd_addr_p1_f == 8'h71; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5334 = _T_4935 ? btb_bank0_rd_data_way0_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5589 = _T_5588 | _T_5334; // @[Mux.scala 27:72]
  wire  _T_4937 = btb_rd_addr_p1_f == 8'h72; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5335 = _T_4937 ? btb_bank0_rd_data_way0_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5590 = _T_5589 | _T_5335; // @[Mux.scala 27:72]
  wire  _T_4939 = btb_rd_addr_p1_f == 8'h73; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5336 = _T_4939 ? btb_bank0_rd_data_way0_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5591 = _T_5590 | _T_5336; // @[Mux.scala 27:72]
  wire  _T_4941 = btb_rd_addr_p1_f == 8'h74; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5337 = _T_4941 ? btb_bank0_rd_data_way0_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5592 = _T_5591 | _T_5337; // @[Mux.scala 27:72]
  wire  _T_4943 = btb_rd_addr_p1_f == 8'h75; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5338 = _T_4943 ? btb_bank0_rd_data_way0_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5593 = _T_5592 | _T_5338; // @[Mux.scala 27:72]
  wire  _T_4945 = btb_rd_addr_p1_f == 8'h76; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5339 = _T_4945 ? btb_bank0_rd_data_way0_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5594 = _T_5593 | _T_5339; // @[Mux.scala 27:72]
  wire  _T_4947 = btb_rd_addr_p1_f == 8'h77; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5340 = _T_4947 ? btb_bank0_rd_data_way0_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5595 = _T_5594 | _T_5340; // @[Mux.scala 27:72]
  wire  _T_4949 = btb_rd_addr_p1_f == 8'h78; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5341 = _T_4949 ? btb_bank0_rd_data_way0_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5596 = _T_5595 | _T_5341; // @[Mux.scala 27:72]
  wire  _T_4951 = btb_rd_addr_p1_f == 8'h79; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5342 = _T_4951 ? btb_bank0_rd_data_way0_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5597 = _T_5596 | _T_5342; // @[Mux.scala 27:72]
  wire  _T_4953 = btb_rd_addr_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5343 = _T_4953 ? btb_bank0_rd_data_way0_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5598 = _T_5597 | _T_5343; // @[Mux.scala 27:72]
  wire  _T_4955 = btb_rd_addr_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5344 = _T_4955 ? btb_bank0_rd_data_way0_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5599 = _T_5598 | _T_5344; // @[Mux.scala 27:72]
  wire  _T_4957 = btb_rd_addr_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5345 = _T_4957 ? btb_bank0_rd_data_way0_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5600 = _T_5599 | _T_5345; // @[Mux.scala 27:72]
  wire  _T_4959 = btb_rd_addr_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5346 = _T_4959 ? btb_bank0_rd_data_way0_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5601 = _T_5600 | _T_5346; // @[Mux.scala 27:72]
  wire  _T_4961 = btb_rd_addr_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5347 = _T_4961 ? btb_bank0_rd_data_way0_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5602 = _T_5601 | _T_5347; // @[Mux.scala 27:72]
  wire  _T_4963 = btb_rd_addr_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5348 = _T_4963 ? btb_bank0_rd_data_way0_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5603 = _T_5602 | _T_5348; // @[Mux.scala 27:72]
  wire  _T_4965 = btb_rd_addr_p1_f == 8'h80; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5349 = _T_4965 ? btb_bank0_rd_data_way0_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5604 = _T_5603 | _T_5349; // @[Mux.scala 27:72]
  wire  _T_4967 = btb_rd_addr_p1_f == 8'h81; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5350 = _T_4967 ? btb_bank0_rd_data_way0_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5605 = _T_5604 | _T_5350; // @[Mux.scala 27:72]
  wire  _T_4969 = btb_rd_addr_p1_f == 8'h82; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5351 = _T_4969 ? btb_bank0_rd_data_way0_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5606 = _T_5605 | _T_5351; // @[Mux.scala 27:72]
  wire  _T_4971 = btb_rd_addr_p1_f == 8'h83; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5352 = _T_4971 ? btb_bank0_rd_data_way0_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5607 = _T_5606 | _T_5352; // @[Mux.scala 27:72]
  wire  _T_4973 = btb_rd_addr_p1_f == 8'h84; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5353 = _T_4973 ? btb_bank0_rd_data_way0_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5608 = _T_5607 | _T_5353; // @[Mux.scala 27:72]
  wire  _T_4975 = btb_rd_addr_p1_f == 8'h85; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5354 = _T_4975 ? btb_bank0_rd_data_way0_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5609 = _T_5608 | _T_5354; // @[Mux.scala 27:72]
  wire  _T_4977 = btb_rd_addr_p1_f == 8'h86; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5355 = _T_4977 ? btb_bank0_rd_data_way0_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5610 = _T_5609 | _T_5355; // @[Mux.scala 27:72]
  wire  _T_4979 = btb_rd_addr_p1_f == 8'h87; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5356 = _T_4979 ? btb_bank0_rd_data_way0_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5611 = _T_5610 | _T_5356; // @[Mux.scala 27:72]
  wire  _T_4981 = btb_rd_addr_p1_f == 8'h88; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5357 = _T_4981 ? btb_bank0_rd_data_way0_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5612 = _T_5611 | _T_5357; // @[Mux.scala 27:72]
  wire  _T_4983 = btb_rd_addr_p1_f == 8'h89; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5358 = _T_4983 ? btb_bank0_rd_data_way0_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5613 = _T_5612 | _T_5358; // @[Mux.scala 27:72]
  wire  _T_4985 = btb_rd_addr_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5359 = _T_4985 ? btb_bank0_rd_data_way0_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5614 = _T_5613 | _T_5359; // @[Mux.scala 27:72]
  wire  _T_4987 = btb_rd_addr_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5360 = _T_4987 ? btb_bank0_rd_data_way0_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5615 = _T_5614 | _T_5360; // @[Mux.scala 27:72]
  wire  _T_4989 = btb_rd_addr_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5361 = _T_4989 ? btb_bank0_rd_data_way0_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5616 = _T_5615 | _T_5361; // @[Mux.scala 27:72]
  wire  _T_4991 = btb_rd_addr_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5362 = _T_4991 ? btb_bank0_rd_data_way0_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5617 = _T_5616 | _T_5362; // @[Mux.scala 27:72]
  wire  _T_4993 = btb_rd_addr_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5363 = _T_4993 ? btb_bank0_rd_data_way0_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5618 = _T_5617 | _T_5363; // @[Mux.scala 27:72]
  wire  _T_4995 = btb_rd_addr_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5364 = _T_4995 ? btb_bank0_rd_data_way0_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5619 = _T_5618 | _T_5364; // @[Mux.scala 27:72]
  wire  _T_4997 = btb_rd_addr_p1_f == 8'h90; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5365 = _T_4997 ? btb_bank0_rd_data_way0_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5620 = _T_5619 | _T_5365; // @[Mux.scala 27:72]
  wire  _T_4999 = btb_rd_addr_p1_f == 8'h91; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5366 = _T_4999 ? btb_bank0_rd_data_way0_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5621 = _T_5620 | _T_5366; // @[Mux.scala 27:72]
  wire  _T_5001 = btb_rd_addr_p1_f == 8'h92; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5367 = _T_5001 ? btb_bank0_rd_data_way0_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5622 = _T_5621 | _T_5367; // @[Mux.scala 27:72]
  wire  _T_5003 = btb_rd_addr_p1_f == 8'h93; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5368 = _T_5003 ? btb_bank0_rd_data_way0_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5623 = _T_5622 | _T_5368; // @[Mux.scala 27:72]
  wire  _T_5005 = btb_rd_addr_p1_f == 8'h94; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5369 = _T_5005 ? btb_bank0_rd_data_way0_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5624 = _T_5623 | _T_5369; // @[Mux.scala 27:72]
  wire  _T_5007 = btb_rd_addr_p1_f == 8'h95; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5370 = _T_5007 ? btb_bank0_rd_data_way0_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5625 = _T_5624 | _T_5370; // @[Mux.scala 27:72]
  wire  _T_5009 = btb_rd_addr_p1_f == 8'h96; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5371 = _T_5009 ? btb_bank0_rd_data_way0_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5626 = _T_5625 | _T_5371; // @[Mux.scala 27:72]
  wire  _T_5011 = btb_rd_addr_p1_f == 8'h97; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5372 = _T_5011 ? btb_bank0_rd_data_way0_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5627 = _T_5626 | _T_5372; // @[Mux.scala 27:72]
  wire  _T_5013 = btb_rd_addr_p1_f == 8'h98; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5373 = _T_5013 ? btb_bank0_rd_data_way0_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5628 = _T_5627 | _T_5373; // @[Mux.scala 27:72]
  wire  _T_5015 = btb_rd_addr_p1_f == 8'h99; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5374 = _T_5015 ? btb_bank0_rd_data_way0_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5629 = _T_5628 | _T_5374; // @[Mux.scala 27:72]
  wire  _T_5017 = btb_rd_addr_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5375 = _T_5017 ? btb_bank0_rd_data_way0_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5630 = _T_5629 | _T_5375; // @[Mux.scala 27:72]
  wire  _T_5019 = btb_rd_addr_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5376 = _T_5019 ? btb_bank0_rd_data_way0_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5631 = _T_5630 | _T_5376; // @[Mux.scala 27:72]
  wire  _T_5021 = btb_rd_addr_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5377 = _T_5021 ? btb_bank0_rd_data_way0_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5632 = _T_5631 | _T_5377; // @[Mux.scala 27:72]
  wire  _T_5023 = btb_rd_addr_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5378 = _T_5023 ? btb_bank0_rd_data_way0_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5633 = _T_5632 | _T_5378; // @[Mux.scala 27:72]
  wire  _T_5025 = btb_rd_addr_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5379 = _T_5025 ? btb_bank0_rd_data_way0_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5634 = _T_5633 | _T_5379; // @[Mux.scala 27:72]
  wire  _T_5027 = btb_rd_addr_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5380 = _T_5027 ? btb_bank0_rd_data_way0_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5635 = _T_5634 | _T_5380; // @[Mux.scala 27:72]
  wire  _T_5029 = btb_rd_addr_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5381 = _T_5029 ? btb_bank0_rd_data_way0_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5636 = _T_5635 | _T_5381; // @[Mux.scala 27:72]
  wire  _T_5031 = btb_rd_addr_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5382 = _T_5031 ? btb_bank0_rd_data_way0_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5637 = _T_5636 | _T_5382; // @[Mux.scala 27:72]
  wire  _T_5033 = btb_rd_addr_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5383 = _T_5033 ? btb_bank0_rd_data_way0_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5638 = _T_5637 | _T_5383; // @[Mux.scala 27:72]
  wire  _T_5035 = btb_rd_addr_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5384 = _T_5035 ? btb_bank0_rd_data_way0_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5639 = _T_5638 | _T_5384; // @[Mux.scala 27:72]
  wire  _T_5037 = btb_rd_addr_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5385 = _T_5037 ? btb_bank0_rd_data_way0_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5640 = _T_5639 | _T_5385; // @[Mux.scala 27:72]
  wire  _T_5039 = btb_rd_addr_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5386 = _T_5039 ? btb_bank0_rd_data_way0_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5641 = _T_5640 | _T_5386; // @[Mux.scala 27:72]
  wire  _T_5041 = btb_rd_addr_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5387 = _T_5041 ? btb_bank0_rd_data_way0_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5642 = _T_5641 | _T_5387; // @[Mux.scala 27:72]
  wire  _T_5043 = btb_rd_addr_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5388 = _T_5043 ? btb_bank0_rd_data_way0_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5643 = _T_5642 | _T_5388; // @[Mux.scala 27:72]
  wire  _T_5045 = btb_rd_addr_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5389 = _T_5045 ? btb_bank0_rd_data_way0_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5644 = _T_5643 | _T_5389; // @[Mux.scala 27:72]
  wire  _T_5047 = btb_rd_addr_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5390 = _T_5047 ? btb_bank0_rd_data_way0_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5645 = _T_5644 | _T_5390; // @[Mux.scala 27:72]
  wire  _T_5049 = btb_rd_addr_p1_f == 8'haa; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5391 = _T_5049 ? btb_bank0_rd_data_way0_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5646 = _T_5645 | _T_5391; // @[Mux.scala 27:72]
  wire  _T_5051 = btb_rd_addr_p1_f == 8'hab; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5392 = _T_5051 ? btb_bank0_rd_data_way0_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5647 = _T_5646 | _T_5392; // @[Mux.scala 27:72]
  wire  _T_5053 = btb_rd_addr_p1_f == 8'hac; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5393 = _T_5053 ? btb_bank0_rd_data_way0_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5648 = _T_5647 | _T_5393; // @[Mux.scala 27:72]
  wire  _T_5055 = btb_rd_addr_p1_f == 8'had; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5394 = _T_5055 ? btb_bank0_rd_data_way0_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5649 = _T_5648 | _T_5394; // @[Mux.scala 27:72]
  wire  _T_5057 = btb_rd_addr_p1_f == 8'hae; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5395 = _T_5057 ? btb_bank0_rd_data_way0_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5650 = _T_5649 | _T_5395; // @[Mux.scala 27:72]
  wire  _T_5059 = btb_rd_addr_p1_f == 8'haf; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5396 = _T_5059 ? btb_bank0_rd_data_way0_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5651 = _T_5650 | _T_5396; // @[Mux.scala 27:72]
  wire  _T_5061 = btb_rd_addr_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5397 = _T_5061 ? btb_bank0_rd_data_way0_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5652 = _T_5651 | _T_5397; // @[Mux.scala 27:72]
  wire  _T_5063 = btb_rd_addr_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5398 = _T_5063 ? btb_bank0_rd_data_way0_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5653 = _T_5652 | _T_5398; // @[Mux.scala 27:72]
  wire  _T_5065 = btb_rd_addr_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5399 = _T_5065 ? btb_bank0_rd_data_way0_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5654 = _T_5653 | _T_5399; // @[Mux.scala 27:72]
  wire  _T_5067 = btb_rd_addr_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5400 = _T_5067 ? btb_bank0_rd_data_way0_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5655 = _T_5654 | _T_5400; // @[Mux.scala 27:72]
  wire  _T_5069 = btb_rd_addr_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5401 = _T_5069 ? btb_bank0_rd_data_way0_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5656 = _T_5655 | _T_5401; // @[Mux.scala 27:72]
  wire  _T_5071 = btb_rd_addr_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5402 = _T_5071 ? btb_bank0_rd_data_way0_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5657 = _T_5656 | _T_5402; // @[Mux.scala 27:72]
  wire  _T_5073 = btb_rd_addr_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5403 = _T_5073 ? btb_bank0_rd_data_way0_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5658 = _T_5657 | _T_5403; // @[Mux.scala 27:72]
  wire  _T_5075 = btb_rd_addr_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5404 = _T_5075 ? btb_bank0_rd_data_way0_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5659 = _T_5658 | _T_5404; // @[Mux.scala 27:72]
  wire  _T_5077 = btb_rd_addr_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5405 = _T_5077 ? btb_bank0_rd_data_way0_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5660 = _T_5659 | _T_5405; // @[Mux.scala 27:72]
  wire  _T_5079 = btb_rd_addr_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5406 = _T_5079 ? btb_bank0_rd_data_way0_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5661 = _T_5660 | _T_5406; // @[Mux.scala 27:72]
  wire  _T_5081 = btb_rd_addr_p1_f == 8'hba; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5407 = _T_5081 ? btb_bank0_rd_data_way0_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5662 = _T_5661 | _T_5407; // @[Mux.scala 27:72]
  wire  _T_5083 = btb_rd_addr_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5408 = _T_5083 ? btb_bank0_rd_data_way0_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5663 = _T_5662 | _T_5408; // @[Mux.scala 27:72]
  wire  _T_5085 = btb_rd_addr_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5409 = _T_5085 ? btb_bank0_rd_data_way0_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5664 = _T_5663 | _T_5409; // @[Mux.scala 27:72]
  wire  _T_5087 = btb_rd_addr_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5410 = _T_5087 ? btb_bank0_rd_data_way0_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5665 = _T_5664 | _T_5410; // @[Mux.scala 27:72]
  wire  _T_5089 = btb_rd_addr_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5411 = _T_5089 ? btb_bank0_rd_data_way0_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5666 = _T_5665 | _T_5411; // @[Mux.scala 27:72]
  wire  _T_5091 = btb_rd_addr_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5412 = _T_5091 ? btb_bank0_rd_data_way0_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5667 = _T_5666 | _T_5412; // @[Mux.scala 27:72]
  wire  _T_5093 = btb_rd_addr_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5413 = _T_5093 ? btb_bank0_rd_data_way0_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5668 = _T_5667 | _T_5413; // @[Mux.scala 27:72]
  wire  _T_5095 = btb_rd_addr_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5414 = _T_5095 ? btb_bank0_rd_data_way0_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5669 = _T_5668 | _T_5414; // @[Mux.scala 27:72]
  wire  _T_5097 = btb_rd_addr_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5415 = _T_5097 ? btb_bank0_rd_data_way0_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5670 = _T_5669 | _T_5415; // @[Mux.scala 27:72]
  wire  _T_5099 = btb_rd_addr_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5416 = _T_5099 ? btb_bank0_rd_data_way0_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5671 = _T_5670 | _T_5416; // @[Mux.scala 27:72]
  wire  _T_5101 = btb_rd_addr_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5417 = _T_5101 ? btb_bank0_rd_data_way0_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5672 = _T_5671 | _T_5417; // @[Mux.scala 27:72]
  wire  _T_5103 = btb_rd_addr_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5418 = _T_5103 ? btb_bank0_rd_data_way0_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5673 = _T_5672 | _T_5418; // @[Mux.scala 27:72]
  wire  _T_5105 = btb_rd_addr_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5419 = _T_5105 ? btb_bank0_rd_data_way0_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5674 = _T_5673 | _T_5419; // @[Mux.scala 27:72]
  wire  _T_5107 = btb_rd_addr_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5420 = _T_5107 ? btb_bank0_rd_data_way0_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5675 = _T_5674 | _T_5420; // @[Mux.scala 27:72]
  wire  _T_5109 = btb_rd_addr_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5421 = _T_5109 ? btb_bank0_rd_data_way0_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5676 = _T_5675 | _T_5421; // @[Mux.scala 27:72]
  wire  _T_5111 = btb_rd_addr_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5422 = _T_5111 ? btb_bank0_rd_data_way0_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5677 = _T_5676 | _T_5422; // @[Mux.scala 27:72]
  wire  _T_5113 = btb_rd_addr_p1_f == 8'hca; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5423 = _T_5113 ? btb_bank0_rd_data_way0_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5678 = _T_5677 | _T_5423; // @[Mux.scala 27:72]
  wire  _T_5115 = btb_rd_addr_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5424 = _T_5115 ? btb_bank0_rd_data_way0_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5679 = _T_5678 | _T_5424; // @[Mux.scala 27:72]
  wire  _T_5117 = btb_rd_addr_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5425 = _T_5117 ? btb_bank0_rd_data_way0_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5680 = _T_5679 | _T_5425; // @[Mux.scala 27:72]
  wire  _T_5119 = btb_rd_addr_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5426 = _T_5119 ? btb_bank0_rd_data_way0_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5681 = _T_5680 | _T_5426; // @[Mux.scala 27:72]
  wire  _T_5121 = btb_rd_addr_p1_f == 8'hce; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5427 = _T_5121 ? btb_bank0_rd_data_way0_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5682 = _T_5681 | _T_5427; // @[Mux.scala 27:72]
  wire  _T_5123 = btb_rd_addr_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5428 = _T_5123 ? btb_bank0_rd_data_way0_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5683 = _T_5682 | _T_5428; // @[Mux.scala 27:72]
  wire  _T_5125 = btb_rd_addr_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5429 = _T_5125 ? btb_bank0_rd_data_way0_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5684 = _T_5683 | _T_5429; // @[Mux.scala 27:72]
  wire  _T_5127 = btb_rd_addr_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5430 = _T_5127 ? btb_bank0_rd_data_way0_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5685 = _T_5684 | _T_5430; // @[Mux.scala 27:72]
  wire  _T_5129 = btb_rd_addr_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5431 = _T_5129 ? btb_bank0_rd_data_way0_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5686 = _T_5685 | _T_5431; // @[Mux.scala 27:72]
  wire  _T_5131 = btb_rd_addr_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5432 = _T_5131 ? btb_bank0_rd_data_way0_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5687 = _T_5686 | _T_5432; // @[Mux.scala 27:72]
  wire  _T_5133 = btb_rd_addr_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5433 = _T_5133 ? btb_bank0_rd_data_way0_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5688 = _T_5687 | _T_5433; // @[Mux.scala 27:72]
  wire  _T_5135 = btb_rd_addr_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5434 = _T_5135 ? btb_bank0_rd_data_way0_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5689 = _T_5688 | _T_5434; // @[Mux.scala 27:72]
  wire  _T_5137 = btb_rd_addr_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5435 = _T_5137 ? btb_bank0_rd_data_way0_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5690 = _T_5689 | _T_5435; // @[Mux.scala 27:72]
  wire  _T_5139 = btb_rd_addr_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5436 = _T_5139 ? btb_bank0_rd_data_way0_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5691 = _T_5690 | _T_5436; // @[Mux.scala 27:72]
  wire  _T_5141 = btb_rd_addr_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5437 = _T_5141 ? btb_bank0_rd_data_way0_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5692 = _T_5691 | _T_5437; // @[Mux.scala 27:72]
  wire  _T_5143 = btb_rd_addr_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5438 = _T_5143 ? btb_bank0_rd_data_way0_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5693 = _T_5692 | _T_5438; // @[Mux.scala 27:72]
  wire  _T_5145 = btb_rd_addr_p1_f == 8'hda; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5439 = _T_5145 ? btb_bank0_rd_data_way0_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5694 = _T_5693 | _T_5439; // @[Mux.scala 27:72]
  wire  _T_5147 = btb_rd_addr_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5440 = _T_5147 ? btb_bank0_rd_data_way0_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5695 = _T_5694 | _T_5440; // @[Mux.scala 27:72]
  wire  _T_5149 = btb_rd_addr_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5441 = _T_5149 ? btb_bank0_rd_data_way0_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5696 = _T_5695 | _T_5441; // @[Mux.scala 27:72]
  wire  _T_5151 = btb_rd_addr_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5442 = _T_5151 ? btb_bank0_rd_data_way0_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5697 = _T_5696 | _T_5442; // @[Mux.scala 27:72]
  wire  _T_5153 = btb_rd_addr_p1_f == 8'hde; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5443 = _T_5153 ? btb_bank0_rd_data_way0_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5698 = _T_5697 | _T_5443; // @[Mux.scala 27:72]
  wire  _T_5155 = btb_rd_addr_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5444 = _T_5155 ? btb_bank0_rd_data_way0_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5699 = _T_5698 | _T_5444; // @[Mux.scala 27:72]
  wire  _T_5157 = btb_rd_addr_p1_f == 8'he0; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5445 = _T_5157 ? btb_bank0_rd_data_way0_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5700 = _T_5699 | _T_5445; // @[Mux.scala 27:72]
  wire  _T_5159 = btb_rd_addr_p1_f == 8'he1; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5446 = _T_5159 ? btb_bank0_rd_data_way0_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5701 = _T_5700 | _T_5446; // @[Mux.scala 27:72]
  wire  _T_5161 = btb_rd_addr_p1_f == 8'he2; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5447 = _T_5161 ? btb_bank0_rd_data_way0_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5702 = _T_5701 | _T_5447; // @[Mux.scala 27:72]
  wire  _T_5163 = btb_rd_addr_p1_f == 8'he3; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5448 = _T_5163 ? btb_bank0_rd_data_way0_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5703 = _T_5702 | _T_5448; // @[Mux.scala 27:72]
  wire  _T_5165 = btb_rd_addr_p1_f == 8'he4; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5449 = _T_5165 ? btb_bank0_rd_data_way0_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5704 = _T_5703 | _T_5449; // @[Mux.scala 27:72]
  wire  _T_5167 = btb_rd_addr_p1_f == 8'he5; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5450 = _T_5167 ? btb_bank0_rd_data_way0_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5705 = _T_5704 | _T_5450; // @[Mux.scala 27:72]
  wire  _T_5169 = btb_rd_addr_p1_f == 8'he6; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5451 = _T_5169 ? btb_bank0_rd_data_way0_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5706 = _T_5705 | _T_5451; // @[Mux.scala 27:72]
  wire  _T_5171 = btb_rd_addr_p1_f == 8'he7; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5452 = _T_5171 ? btb_bank0_rd_data_way0_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5707 = _T_5706 | _T_5452; // @[Mux.scala 27:72]
  wire  _T_5173 = btb_rd_addr_p1_f == 8'he8; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5453 = _T_5173 ? btb_bank0_rd_data_way0_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5708 = _T_5707 | _T_5453; // @[Mux.scala 27:72]
  wire  _T_5175 = btb_rd_addr_p1_f == 8'he9; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5454 = _T_5175 ? btb_bank0_rd_data_way0_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5709 = _T_5708 | _T_5454; // @[Mux.scala 27:72]
  wire  _T_5177 = btb_rd_addr_p1_f == 8'hea; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5455 = _T_5177 ? btb_bank0_rd_data_way0_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5710 = _T_5709 | _T_5455; // @[Mux.scala 27:72]
  wire  _T_5179 = btb_rd_addr_p1_f == 8'heb; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5456 = _T_5179 ? btb_bank0_rd_data_way0_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5711 = _T_5710 | _T_5456; // @[Mux.scala 27:72]
  wire  _T_5181 = btb_rd_addr_p1_f == 8'hec; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5457 = _T_5181 ? btb_bank0_rd_data_way0_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5712 = _T_5711 | _T_5457; // @[Mux.scala 27:72]
  wire  _T_5183 = btb_rd_addr_p1_f == 8'hed; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5458 = _T_5183 ? btb_bank0_rd_data_way0_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5713 = _T_5712 | _T_5458; // @[Mux.scala 27:72]
  wire  _T_5185 = btb_rd_addr_p1_f == 8'hee; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5459 = _T_5185 ? btb_bank0_rd_data_way0_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5714 = _T_5713 | _T_5459; // @[Mux.scala 27:72]
  wire  _T_5187 = btb_rd_addr_p1_f == 8'hef; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5460 = _T_5187 ? btb_bank0_rd_data_way0_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5715 = _T_5714 | _T_5460; // @[Mux.scala 27:72]
  wire  _T_5189 = btb_rd_addr_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5461 = _T_5189 ? btb_bank0_rd_data_way0_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5716 = _T_5715 | _T_5461; // @[Mux.scala 27:72]
  wire  _T_5191 = btb_rd_addr_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5462 = _T_5191 ? btb_bank0_rd_data_way0_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5717 = _T_5716 | _T_5462; // @[Mux.scala 27:72]
  wire  _T_5193 = btb_rd_addr_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5463 = _T_5193 ? btb_bank0_rd_data_way0_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5718 = _T_5717 | _T_5463; // @[Mux.scala 27:72]
  wire  _T_5195 = btb_rd_addr_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5464 = _T_5195 ? btb_bank0_rd_data_way0_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5719 = _T_5718 | _T_5464; // @[Mux.scala 27:72]
  wire  _T_5197 = btb_rd_addr_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5465 = _T_5197 ? btb_bank0_rd_data_way0_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5720 = _T_5719 | _T_5465; // @[Mux.scala 27:72]
  wire  _T_5199 = btb_rd_addr_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5466 = _T_5199 ? btb_bank0_rd_data_way0_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5721 = _T_5720 | _T_5466; // @[Mux.scala 27:72]
  wire  _T_5201 = btb_rd_addr_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5467 = _T_5201 ? btb_bank0_rd_data_way0_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5722 = _T_5721 | _T_5467; // @[Mux.scala 27:72]
  wire  _T_5203 = btb_rd_addr_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5468 = _T_5203 ? btb_bank0_rd_data_way0_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5723 = _T_5722 | _T_5468; // @[Mux.scala 27:72]
  wire  _T_5205 = btb_rd_addr_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5469 = _T_5205 ? btb_bank0_rd_data_way0_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5724 = _T_5723 | _T_5469; // @[Mux.scala 27:72]
  wire  _T_5207 = btb_rd_addr_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5470 = _T_5207 ? btb_bank0_rd_data_way0_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5725 = _T_5724 | _T_5470; // @[Mux.scala 27:72]
  wire  _T_5209 = btb_rd_addr_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5471 = _T_5209 ? btb_bank0_rd_data_way0_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5726 = _T_5725 | _T_5471; // @[Mux.scala 27:72]
  wire  _T_5211 = btb_rd_addr_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5472 = _T_5211 ? btb_bank0_rd_data_way0_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5727 = _T_5726 | _T_5472; // @[Mux.scala 27:72]
  wire  _T_5213 = btb_rd_addr_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5473 = _T_5213 ? btb_bank0_rd_data_way0_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5728 = _T_5727 | _T_5473; // @[Mux.scala 27:72]
  wire  _T_5215 = btb_rd_addr_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5474 = _T_5215 ? btb_bank0_rd_data_way0_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5729 = _T_5728 | _T_5474; // @[Mux.scala 27:72]
  wire  _T_5217 = btb_rd_addr_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5475 = _T_5217 ? btb_bank0_rd_data_way0_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_5730 = _T_5729 | _T_5475; // @[Mux.scala 27:72]
  wire  _T_5219 = btb_rd_addr_p1_f == 8'hff; // @[ifu_bp_ctl.scala 439:86]
  wire [21:0] _T_5476 = _T_5219 ? btb_bank0_rd_data_way0_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way0_p1_f = _T_5730 | _T_5476; // @[Mux.scala 27:72]
  wire [4:0] _T_35 = _T_8[13:9] ^ _T_8[18:14]; // @[lib.scala 42:111]
  wire [4:0] fetch_rd_tag_p1_f = _T_35 ^ _T_8[23:19]; // @[lib.scala 42:111]
  wire  _T_64 = btb_bank0_rd_data_way0_p1_f[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 152:107]
  wire  _T_65 = btb_bank0_rd_data_way0_p1_f[0] & _T_64; // @[ifu_bp_ctl.scala 152:61]
  wire  _T_20 = io_exu_bp_exu_i0_br_index_r == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 126:75]
  wire  branch_error_collision_p1_f = dec_tlu_error_wb & _T_20; // @[ifu_bp_ctl.scala 126:54]
  wire  branch_error_bank_conflict_p1_f = branch_error_collision_p1_f & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 130:69]
  wire  _T_66 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & branch_error_bank_conflict_p1_f; // @[ifu_bp_ctl.scala 153:22]
  wire  _T_67 = ~_T_66; // @[ifu_bp_ctl.scala 153:5]
  wire  _T_68 = _T_65 & _T_67; // @[ifu_bp_ctl.scala 152:130]
  wire  _T_69 = _T_68 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 153:57]
  wire  tag_match_way0_p1_f = _T_69 & _T; // @[ifu_bp_ctl.scala 153:78]
  wire  _T_100 = btb_bank0_rd_data_way0_p1_f[3] ^ btb_bank0_rd_data_way0_p1_f[4]; // @[ifu_bp_ctl.scala 165:99]
  wire  _T_101 = tag_match_way0_p1_f & _T_100; // @[ifu_bp_ctl.scala 165:62]
  wire  _T_105 = ~_T_100; // @[ifu_bp_ctl.scala 166:27]
  wire  _T_106 = tag_match_way0_p1_f & _T_105; // @[ifu_bp_ctl.scala 166:25]
  wire [1:0] tag_match_way0_expanded_p1_f = {_T_101,_T_106}; // @[Cat.scala 29:58]
  wire [21:0] _T_136 = tag_match_way0_expanded_p1_f[0] ? btb_bank0_rd_data_way0_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6245 = _T_4709 ? btb_bank0_rd_data_way1_out_0 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6246 = _T_4711 ? btb_bank0_rd_data_way1_out_1 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6501 = _T_6245 | _T_6246; // @[Mux.scala 27:72]
  wire [21:0] _T_6247 = _T_4713 ? btb_bank0_rd_data_way1_out_2 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6502 = _T_6501 | _T_6247; // @[Mux.scala 27:72]
  wire [21:0] _T_6248 = _T_4715 ? btb_bank0_rd_data_way1_out_3 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6503 = _T_6502 | _T_6248; // @[Mux.scala 27:72]
  wire [21:0] _T_6249 = _T_4717 ? btb_bank0_rd_data_way1_out_4 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6504 = _T_6503 | _T_6249; // @[Mux.scala 27:72]
  wire [21:0] _T_6250 = _T_4719 ? btb_bank0_rd_data_way1_out_5 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6505 = _T_6504 | _T_6250; // @[Mux.scala 27:72]
  wire [21:0] _T_6251 = _T_4721 ? btb_bank0_rd_data_way1_out_6 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6506 = _T_6505 | _T_6251; // @[Mux.scala 27:72]
  wire [21:0] _T_6252 = _T_4723 ? btb_bank0_rd_data_way1_out_7 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6507 = _T_6506 | _T_6252; // @[Mux.scala 27:72]
  wire [21:0] _T_6253 = _T_4725 ? btb_bank0_rd_data_way1_out_8 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6508 = _T_6507 | _T_6253; // @[Mux.scala 27:72]
  wire [21:0] _T_6254 = _T_4727 ? btb_bank0_rd_data_way1_out_9 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6509 = _T_6508 | _T_6254; // @[Mux.scala 27:72]
  wire [21:0] _T_6255 = _T_4729 ? btb_bank0_rd_data_way1_out_10 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6510 = _T_6509 | _T_6255; // @[Mux.scala 27:72]
  wire [21:0] _T_6256 = _T_4731 ? btb_bank0_rd_data_way1_out_11 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6511 = _T_6510 | _T_6256; // @[Mux.scala 27:72]
  wire [21:0] _T_6257 = _T_4733 ? btb_bank0_rd_data_way1_out_12 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6512 = _T_6511 | _T_6257; // @[Mux.scala 27:72]
  wire [21:0] _T_6258 = _T_4735 ? btb_bank0_rd_data_way1_out_13 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6513 = _T_6512 | _T_6258; // @[Mux.scala 27:72]
  wire [21:0] _T_6259 = _T_4737 ? btb_bank0_rd_data_way1_out_14 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6514 = _T_6513 | _T_6259; // @[Mux.scala 27:72]
  wire [21:0] _T_6260 = _T_4739 ? btb_bank0_rd_data_way1_out_15 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6515 = _T_6514 | _T_6260; // @[Mux.scala 27:72]
  wire [21:0] _T_6261 = _T_4741 ? btb_bank0_rd_data_way1_out_16 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6516 = _T_6515 | _T_6261; // @[Mux.scala 27:72]
  wire [21:0] _T_6262 = _T_4743 ? btb_bank0_rd_data_way1_out_17 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6517 = _T_6516 | _T_6262; // @[Mux.scala 27:72]
  wire [21:0] _T_6263 = _T_4745 ? btb_bank0_rd_data_way1_out_18 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6518 = _T_6517 | _T_6263; // @[Mux.scala 27:72]
  wire [21:0] _T_6264 = _T_4747 ? btb_bank0_rd_data_way1_out_19 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6519 = _T_6518 | _T_6264; // @[Mux.scala 27:72]
  wire [21:0] _T_6265 = _T_4749 ? btb_bank0_rd_data_way1_out_20 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6520 = _T_6519 | _T_6265; // @[Mux.scala 27:72]
  wire [21:0] _T_6266 = _T_4751 ? btb_bank0_rd_data_way1_out_21 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6521 = _T_6520 | _T_6266; // @[Mux.scala 27:72]
  wire [21:0] _T_6267 = _T_4753 ? btb_bank0_rd_data_way1_out_22 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6522 = _T_6521 | _T_6267; // @[Mux.scala 27:72]
  wire [21:0] _T_6268 = _T_4755 ? btb_bank0_rd_data_way1_out_23 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6523 = _T_6522 | _T_6268; // @[Mux.scala 27:72]
  wire [21:0] _T_6269 = _T_4757 ? btb_bank0_rd_data_way1_out_24 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6524 = _T_6523 | _T_6269; // @[Mux.scala 27:72]
  wire [21:0] _T_6270 = _T_4759 ? btb_bank0_rd_data_way1_out_25 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6525 = _T_6524 | _T_6270; // @[Mux.scala 27:72]
  wire [21:0] _T_6271 = _T_4761 ? btb_bank0_rd_data_way1_out_26 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6526 = _T_6525 | _T_6271; // @[Mux.scala 27:72]
  wire [21:0] _T_6272 = _T_4763 ? btb_bank0_rd_data_way1_out_27 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6527 = _T_6526 | _T_6272; // @[Mux.scala 27:72]
  wire [21:0] _T_6273 = _T_4765 ? btb_bank0_rd_data_way1_out_28 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6528 = _T_6527 | _T_6273; // @[Mux.scala 27:72]
  wire [21:0] _T_6274 = _T_4767 ? btb_bank0_rd_data_way1_out_29 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6529 = _T_6528 | _T_6274; // @[Mux.scala 27:72]
  wire [21:0] _T_6275 = _T_4769 ? btb_bank0_rd_data_way1_out_30 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6530 = _T_6529 | _T_6275; // @[Mux.scala 27:72]
  wire [21:0] _T_6276 = _T_4771 ? btb_bank0_rd_data_way1_out_31 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6531 = _T_6530 | _T_6276; // @[Mux.scala 27:72]
  wire [21:0] _T_6277 = _T_4773 ? btb_bank0_rd_data_way1_out_32 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6532 = _T_6531 | _T_6277; // @[Mux.scala 27:72]
  wire [21:0] _T_6278 = _T_4775 ? btb_bank0_rd_data_way1_out_33 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6533 = _T_6532 | _T_6278; // @[Mux.scala 27:72]
  wire [21:0] _T_6279 = _T_4777 ? btb_bank0_rd_data_way1_out_34 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6534 = _T_6533 | _T_6279; // @[Mux.scala 27:72]
  wire [21:0] _T_6280 = _T_4779 ? btb_bank0_rd_data_way1_out_35 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6535 = _T_6534 | _T_6280; // @[Mux.scala 27:72]
  wire [21:0] _T_6281 = _T_4781 ? btb_bank0_rd_data_way1_out_36 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6536 = _T_6535 | _T_6281; // @[Mux.scala 27:72]
  wire [21:0] _T_6282 = _T_4783 ? btb_bank0_rd_data_way1_out_37 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6537 = _T_6536 | _T_6282; // @[Mux.scala 27:72]
  wire [21:0] _T_6283 = _T_4785 ? btb_bank0_rd_data_way1_out_38 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6538 = _T_6537 | _T_6283; // @[Mux.scala 27:72]
  wire [21:0] _T_6284 = _T_4787 ? btb_bank0_rd_data_way1_out_39 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6539 = _T_6538 | _T_6284; // @[Mux.scala 27:72]
  wire [21:0] _T_6285 = _T_4789 ? btb_bank0_rd_data_way1_out_40 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6540 = _T_6539 | _T_6285; // @[Mux.scala 27:72]
  wire [21:0] _T_6286 = _T_4791 ? btb_bank0_rd_data_way1_out_41 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6541 = _T_6540 | _T_6286; // @[Mux.scala 27:72]
  wire [21:0] _T_6287 = _T_4793 ? btb_bank0_rd_data_way1_out_42 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6542 = _T_6541 | _T_6287; // @[Mux.scala 27:72]
  wire [21:0] _T_6288 = _T_4795 ? btb_bank0_rd_data_way1_out_43 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6543 = _T_6542 | _T_6288; // @[Mux.scala 27:72]
  wire [21:0] _T_6289 = _T_4797 ? btb_bank0_rd_data_way1_out_44 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6544 = _T_6543 | _T_6289; // @[Mux.scala 27:72]
  wire [21:0] _T_6290 = _T_4799 ? btb_bank0_rd_data_way1_out_45 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6545 = _T_6544 | _T_6290; // @[Mux.scala 27:72]
  wire [21:0] _T_6291 = _T_4801 ? btb_bank0_rd_data_way1_out_46 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6546 = _T_6545 | _T_6291; // @[Mux.scala 27:72]
  wire [21:0] _T_6292 = _T_4803 ? btb_bank0_rd_data_way1_out_47 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6547 = _T_6546 | _T_6292; // @[Mux.scala 27:72]
  wire [21:0] _T_6293 = _T_4805 ? btb_bank0_rd_data_way1_out_48 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6548 = _T_6547 | _T_6293; // @[Mux.scala 27:72]
  wire [21:0] _T_6294 = _T_4807 ? btb_bank0_rd_data_way1_out_49 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6549 = _T_6548 | _T_6294; // @[Mux.scala 27:72]
  wire [21:0] _T_6295 = _T_4809 ? btb_bank0_rd_data_way1_out_50 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6550 = _T_6549 | _T_6295; // @[Mux.scala 27:72]
  wire [21:0] _T_6296 = _T_4811 ? btb_bank0_rd_data_way1_out_51 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6551 = _T_6550 | _T_6296; // @[Mux.scala 27:72]
  wire [21:0] _T_6297 = _T_4813 ? btb_bank0_rd_data_way1_out_52 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6552 = _T_6551 | _T_6297; // @[Mux.scala 27:72]
  wire [21:0] _T_6298 = _T_4815 ? btb_bank0_rd_data_way1_out_53 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6553 = _T_6552 | _T_6298; // @[Mux.scala 27:72]
  wire [21:0] _T_6299 = _T_4817 ? btb_bank0_rd_data_way1_out_54 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6554 = _T_6553 | _T_6299; // @[Mux.scala 27:72]
  wire [21:0] _T_6300 = _T_4819 ? btb_bank0_rd_data_way1_out_55 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6555 = _T_6554 | _T_6300; // @[Mux.scala 27:72]
  wire [21:0] _T_6301 = _T_4821 ? btb_bank0_rd_data_way1_out_56 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6556 = _T_6555 | _T_6301; // @[Mux.scala 27:72]
  wire [21:0] _T_6302 = _T_4823 ? btb_bank0_rd_data_way1_out_57 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6557 = _T_6556 | _T_6302; // @[Mux.scala 27:72]
  wire [21:0] _T_6303 = _T_4825 ? btb_bank0_rd_data_way1_out_58 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6558 = _T_6557 | _T_6303; // @[Mux.scala 27:72]
  wire [21:0] _T_6304 = _T_4827 ? btb_bank0_rd_data_way1_out_59 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6559 = _T_6558 | _T_6304; // @[Mux.scala 27:72]
  wire [21:0] _T_6305 = _T_4829 ? btb_bank0_rd_data_way1_out_60 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6560 = _T_6559 | _T_6305; // @[Mux.scala 27:72]
  wire [21:0] _T_6306 = _T_4831 ? btb_bank0_rd_data_way1_out_61 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6561 = _T_6560 | _T_6306; // @[Mux.scala 27:72]
  wire [21:0] _T_6307 = _T_4833 ? btb_bank0_rd_data_way1_out_62 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6562 = _T_6561 | _T_6307; // @[Mux.scala 27:72]
  wire [21:0] _T_6308 = _T_4835 ? btb_bank0_rd_data_way1_out_63 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6563 = _T_6562 | _T_6308; // @[Mux.scala 27:72]
  wire [21:0] _T_6309 = _T_4837 ? btb_bank0_rd_data_way1_out_64 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6564 = _T_6563 | _T_6309; // @[Mux.scala 27:72]
  wire [21:0] _T_6310 = _T_4839 ? btb_bank0_rd_data_way1_out_65 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6565 = _T_6564 | _T_6310; // @[Mux.scala 27:72]
  wire [21:0] _T_6311 = _T_4841 ? btb_bank0_rd_data_way1_out_66 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6566 = _T_6565 | _T_6311; // @[Mux.scala 27:72]
  wire [21:0] _T_6312 = _T_4843 ? btb_bank0_rd_data_way1_out_67 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6567 = _T_6566 | _T_6312; // @[Mux.scala 27:72]
  wire [21:0] _T_6313 = _T_4845 ? btb_bank0_rd_data_way1_out_68 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6568 = _T_6567 | _T_6313; // @[Mux.scala 27:72]
  wire [21:0] _T_6314 = _T_4847 ? btb_bank0_rd_data_way1_out_69 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6569 = _T_6568 | _T_6314; // @[Mux.scala 27:72]
  wire [21:0] _T_6315 = _T_4849 ? btb_bank0_rd_data_way1_out_70 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6570 = _T_6569 | _T_6315; // @[Mux.scala 27:72]
  wire [21:0] _T_6316 = _T_4851 ? btb_bank0_rd_data_way1_out_71 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6571 = _T_6570 | _T_6316; // @[Mux.scala 27:72]
  wire [21:0] _T_6317 = _T_4853 ? btb_bank0_rd_data_way1_out_72 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6572 = _T_6571 | _T_6317; // @[Mux.scala 27:72]
  wire [21:0] _T_6318 = _T_4855 ? btb_bank0_rd_data_way1_out_73 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6573 = _T_6572 | _T_6318; // @[Mux.scala 27:72]
  wire [21:0] _T_6319 = _T_4857 ? btb_bank0_rd_data_way1_out_74 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6574 = _T_6573 | _T_6319; // @[Mux.scala 27:72]
  wire [21:0] _T_6320 = _T_4859 ? btb_bank0_rd_data_way1_out_75 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6575 = _T_6574 | _T_6320; // @[Mux.scala 27:72]
  wire [21:0] _T_6321 = _T_4861 ? btb_bank0_rd_data_way1_out_76 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6576 = _T_6575 | _T_6321; // @[Mux.scala 27:72]
  wire [21:0] _T_6322 = _T_4863 ? btb_bank0_rd_data_way1_out_77 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6577 = _T_6576 | _T_6322; // @[Mux.scala 27:72]
  wire [21:0] _T_6323 = _T_4865 ? btb_bank0_rd_data_way1_out_78 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6578 = _T_6577 | _T_6323; // @[Mux.scala 27:72]
  wire [21:0] _T_6324 = _T_4867 ? btb_bank0_rd_data_way1_out_79 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6579 = _T_6578 | _T_6324; // @[Mux.scala 27:72]
  wire [21:0] _T_6325 = _T_4869 ? btb_bank0_rd_data_way1_out_80 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6580 = _T_6579 | _T_6325; // @[Mux.scala 27:72]
  wire [21:0] _T_6326 = _T_4871 ? btb_bank0_rd_data_way1_out_81 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6581 = _T_6580 | _T_6326; // @[Mux.scala 27:72]
  wire [21:0] _T_6327 = _T_4873 ? btb_bank0_rd_data_way1_out_82 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6582 = _T_6581 | _T_6327; // @[Mux.scala 27:72]
  wire [21:0] _T_6328 = _T_4875 ? btb_bank0_rd_data_way1_out_83 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6583 = _T_6582 | _T_6328; // @[Mux.scala 27:72]
  wire [21:0] _T_6329 = _T_4877 ? btb_bank0_rd_data_way1_out_84 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6584 = _T_6583 | _T_6329; // @[Mux.scala 27:72]
  wire [21:0] _T_6330 = _T_4879 ? btb_bank0_rd_data_way1_out_85 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6585 = _T_6584 | _T_6330; // @[Mux.scala 27:72]
  wire [21:0] _T_6331 = _T_4881 ? btb_bank0_rd_data_way1_out_86 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6586 = _T_6585 | _T_6331; // @[Mux.scala 27:72]
  wire [21:0] _T_6332 = _T_4883 ? btb_bank0_rd_data_way1_out_87 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6587 = _T_6586 | _T_6332; // @[Mux.scala 27:72]
  wire [21:0] _T_6333 = _T_4885 ? btb_bank0_rd_data_way1_out_88 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6588 = _T_6587 | _T_6333; // @[Mux.scala 27:72]
  wire [21:0] _T_6334 = _T_4887 ? btb_bank0_rd_data_way1_out_89 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6589 = _T_6588 | _T_6334; // @[Mux.scala 27:72]
  wire [21:0] _T_6335 = _T_4889 ? btb_bank0_rd_data_way1_out_90 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6590 = _T_6589 | _T_6335; // @[Mux.scala 27:72]
  wire [21:0] _T_6336 = _T_4891 ? btb_bank0_rd_data_way1_out_91 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6591 = _T_6590 | _T_6336; // @[Mux.scala 27:72]
  wire [21:0] _T_6337 = _T_4893 ? btb_bank0_rd_data_way1_out_92 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6592 = _T_6591 | _T_6337; // @[Mux.scala 27:72]
  wire [21:0] _T_6338 = _T_4895 ? btb_bank0_rd_data_way1_out_93 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6593 = _T_6592 | _T_6338; // @[Mux.scala 27:72]
  wire [21:0] _T_6339 = _T_4897 ? btb_bank0_rd_data_way1_out_94 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6594 = _T_6593 | _T_6339; // @[Mux.scala 27:72]
  wire [21:0] _T_6340 = _T_4899 ? btb_bank0_rd_data_way1_out_95 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6595 = _T_6594 | _T_6340; // @[Mux.scala 27:72]
  wire [21:0] _T_6341 = _T_4901 ? btb_bank0_rd_data_way1_out_96 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6596 = _T_6595 | _T_6341; // @[Mux.scala 27:72]
  wire [21:0] _T_6342 = _T_4903 ? btb_bank0_rd_data_way1_out_97 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6597 = _T_6596 | _T_6342; // @[Mux.scala 27:72]
  wire [21:0] _T_6343 = _T_4905 ? btb_bank0_rd_data_way1_out_98 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6598 = _T_6597 | _T_6343; // @[Mux.scala 27:72]
  wire [21:0] _T_6344 = _T_4907 ? btb_bank0_rd_data_way1_out_99 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6599 = _T_6598 | _T_6344; // @[Mux.scala 27:72]
  wire [21:0] _T_6345 = _T_4909 ? btb_bank0_rd_data_way1_out_100 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6600 = _T_6599 | _T_6345; // @[Mux.scala 27:72]
  wire [21:0] _T_6346 = _T_4911 ? btb_bank0_rd_data_way1_out_101 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6601 = _T_6600 | _T_6346; // @[Mux.scala 27:72]
  wire [21:0] _T_6347 = _T_4913 ? btb_bank0_rd_data_way1_out_102 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6602 = _T_6601 | _T_6347; // @[Mux.scala 27:72]
  wire [21:0] _T_6348 = _T_4915 ? btb_bank0_rd_data_way1_out_103 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6603 = _T_6602 | _T_6348; // @[Mux.scala 27:72]
  wire [21:0] _T_6349 = _T_4917 ? btb_bank0_rd_data_way1_out_104 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6604 = _T_6603 | _T_6349; // @[Mux.scala 27:72]
  wire [21:0] _T_6350 = _T_4919 ? btb_bank0_rd_data_way1_out_105 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6605 = _T_6604 | _T_6350; // @[Mux.scala 27:72]
  wire [21:0] _T_6351 = _T_4921 ? btb_bank0_rd_data_way1_out_106 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6606 = _T_6605 | _T_6351; // @[Mux.scala 27:72]
  wire [21:0] _T_6352 = _T_4923 ? btb_bank0_rd_data_way1_out_107 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6607 = _T_6606 | _T_6352; // @[Mux.scala 27:72]
  wire [21:0] _T_6353 = _T_4925 ? btb_bank0_rd_data_way1_out_108 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6608 = _T_6607 | _T_6353; // @[Mux.scala 27:72]
  wire [21:0] _T_6354 = _T_4927 ? btb_bank0_rd_data_way1_out_109 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6609 = _T_6608 | _T_6354; // @[Mux.scala 27:72]
  wire [21:0] _T_6355 = _T_4929 ? btb_bank0_rd_data_way1_out_110 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6610 = _T_6609 | _T_6355; // @[Mux.scala 27:72]
  wire [21:0] _T_6356 = _T_4931 ? btb_bank0_rd_data_way1_out_111 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6611 = _T_6610 | _T_6356; // @[Mux.scala 27:72]
  wire [21:0] _T_6357 = _T_4933 ? btb_bank0_rd_data_way1_out_112 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6612 = _T_6611 | _T_6357; // @[Mux.scala 27:72]
  wire [21:0] _T_6358 = _T_4935 ? btb_bank0_rd_data_way1_out_113 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6613 = _T_6612 | _T_6358; // @[Mux.scala 27:72]
  wire [21:0] _T_6359 = _T_4937 ? btb_bank0_rd_data_way1_out_114 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6614 = _T_6613 | _T_6359; // @[Mux.scala 27:72]
  wire [21:0] _T_6360 = _T_4939 ? btb_bank0_rd_data_way1_out_115 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6615 = _T_6614 | _T_6360; // @[Mux.scala 27:72]
  wire [21:0] _T_6361 = _T_4941 ? btb_bank0_rd_data_way1_out_116 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6616 = _T_6615 | _T_6361; // @[Mux.scala 27:72]
  wire [21:0] _T_6362 = _T_4943 ? btb_bank0_rd_data_way1_out_117 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6617 = _T_6616 | _T_6362; // @[Mux.scala 27:72]
  wire [21:0] _T_6363 = _T_4945 ? btb_bank0_rd_data_way1_out_118 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6618 = _T_6617 | _T_6363; // @[Mux.scala 27:72]
  wire [21:0] _T_6364 = _T_4947 ? btb_bank0_rd_data_way1_out_119 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6619 = _T_6618 | _T_6364; // @[Mux.scala 27:72]
  wire [21:0] _T_6365 = _T_4949 ? btb_bank0_rd_data_way1_out_120 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6620 = _T_6619 | _T_6365; // @[Mux.scala 27:72]
  wire [21:0] _T_6366 = _T_4951 ? btb_bank0_rd_data_way1_out_121 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6621 = _T_6620 | _T_6366; // @[Mux.scala 27:72]
  wire [21:0] _T_6367 = _T_4953 ? btb_bank0_rd_data_way1_out_122 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6622 = _T_6621 | _T_6367; // @[Mux.scala 27:72]
  wire [21:0] _T_6368 = _T_4955 ? btb_bank0_rd_data_way1_out_123 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6623 = _T_6622 | _T_6368; // @[Mux.scala 27:72]
  wire [21:0] _T_6369 = _T_4957 ? btb_bank0_rd_data_way1_out_124 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6624 = _T_6623 | _T_6369; // @[Mux.scala 27:72]
  wire [21:0] _T_6370 = _T_4959 ? btb_bank0_rd_data_way1_out_125 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6625 = _T_6624 | _T_6370; // @[Mux.scala 27:72]
  wire [21:0] _T_6371 = _T_4961 ? btb_bank0_rd_data_way1_out_126 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6626 = _T_6625 | _T_6371; // @[Mux.scala 27:72]
  wire [21:0] _T_6372 = _T_4963 ? btb_bank0_rd_data_way1_out_127 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6627 = _T_6626 | _T_6372; // @[Mux.scala 27:72]
  wire [21:0] _T_6373 = _T_4965 ? btb_bank0_rd_data_way1_out_128 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6628 = _T_6627 | _T_6373; // @[Mux.scala 27:72]
  wire [21:0] _T_6374 = _T_4967 ? btb_bank0_rd_data_way1_out_129 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6629 = _T_6628 | _T_6374; // @[Mux.scala 27:72]
  wire [21:0] _T_6375 = _T_4969 ? btb_bank0_rd_data_way1_out_130 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6630 = _T_6629 | _T_6375; // @[Mux.scala 27:72]
  wire [21:0] _T_6376 = _T_4971 ? btb_bank0_rd_data_way1_out_131 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6631 = _T_6630 | _T_6376; // @[Mux.scala 27:72]
  wire [21:0] _T_6377 = _T_4973 ? btb_bank0_rd_data_way1_out_132 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6632 = _T_6631 | _T_6377; // @[Mux.scala 27:72]
  wire [21:0] _T_6378 = _T_4975 ? btb_bank0_rd_data_way1_out_133 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6633 = _T_6632 | _T_6378; // @[Mux.scala 27:72]
  wire [21:0] _T_6379 = _T_4977 ? btb_bank0_rd_data_way1_out_134 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6634 = _T_6633 | _T_6379; // @[Mux.scala 27:72]
  wire [21:0] _T_6380 = _T_4979 ? btb_bank0_rd_data_way1_out_135 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6635 = _T_6634 | _T_6380; // @[Mux.scala 27:72]
  wire [21:0] _T_6381 = _T_4981 ? btb_bank0_rd_data_way1_out_136 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6636 = _T_6635 | _T_6381; // @[Mux.scala 27:72]
  wire [21:0] _T_6382 = _T_4983 ? btb_bank0_rd_data_way1_out_137 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6637 = _T_6636 | _T_6382; // @[Mux.scala 27:72]
  wire [21:0] _T_6383 = _T_4985 ? btb_bank0_rd_data_way1_out_138 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6638 = _T_6637 | _T_6383; // @[Mux.scala 27:72]
  wire [21:0] _T_6384 = _T_4987 ? btb_bank0_rd_data_way1_out_139 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6639 = _T_6638 | _T_6384; // @[Mux.scala 27:72]
  wire [21:0] _T_6385 = _T_4989 ? btb_bank0_rd_data_way1_out_140 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6640 = _T_6639 | _T_6385; // @[Mux.scala 27:72]
  wire [21:0] _T_6386 = _T_4991 ? btb_bank0_rd_data_way1_out_141 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6641 = _T_6640 | _T_6386; // @[Mux.scala 27:72]
  wire [21:0] _T_6387 = _T_4993 ? btb_bank0_rd_data_way1_out_142 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6642 = _T_6641 | _T_6387; // @[Mux.scala 27:72]
  wire [21:0] _T_6388 = _T_4995 ? btb_bank0_rd_data_way1_out_143 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6643 = _T_6642 | _T_6388; // @[Mux.scala 27:72]
  wire [21:0] _T_6389 = _T_4997 ? btb_bank0_rd_data_way1_out_144 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6644 = _T_6643 | _T_6389; // @[Mux.scala 27:72]
  wire [21:0] _T_6390 = _T_4999 ? btb_bank0_rd_data_way1_out_145 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6645 = _T_6644 | _T_6390; // @[Mux.scala 27:72]
  wire [21:0] _T_6391 = _T_5001 ? btb_bank0_rd_data_way1_out_146 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6646 = _T_6645 | _T_6391; // @[Mux.scala 27:72]
  wire [21:0] _T_6392 = _T_5003 ? btb_bank0_rd_data_way1_out_147 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6647 = _T_6646 | _T_6392; // @[Mux.scala 27:72]
  wire [21:0] _T_6393 = _T_5005 ? btb_bank0_rd_data_way1_out_148 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6648 = _T_6647 | _T_6393; // @[Mux.scala 27:72]
  wire [21:0] _T_6394 = _T_5007 ? btb_bank0_rd_data_way1_out_149 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6649 = _T_6648 | _T_6394; // @[Mux.scala 27:72]
  wire [21:0] _T_6395 = _T_5009 ? btb_bank0_rd_data_way1_out_150 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6650 = _T_6649 | _T_6395; // @[Mux.scala 27:72]
  wire [21:0] _T_6396 = _T_5011 ? btb_bank0_rd_data_way1_out_151 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6651 = _T_6650 | _T_6396; // @[Mux.scala 27:72]
  wire [21:0] _T_6397 = _T_5013 ? btb_bank0_rd_data_way1_out_152 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6652 = _T_6651 | _T_6397; // @[Mux.scala 27:72]
  wire [21:0] _T_6398 = _T_5015 ? btb_bank0_rd_data_way1_out_153 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6653 = _T_6652 | _T_6398; // @[Mux.scala 27:72]
  wire [21:0] _T_6399 = _T_5017 ? btb_bank0_rd_data_way1_out_154 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6654 = _T_6653 | _T_6399; // @[Mux.scala 27:72]
  wire [21:0] _T_6400 = _T_5019 ? btb_bank0_rd_data_way1_out_155 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6655 = _T_6654 | _T_6400; // @[Mux.scala 27:72]
  wire [21:0] _T_6401 = _T_5021 ? btb_bank0_rd_data_way1_out_156 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6656 = _T_6655 | _T_6401; // @[Mux.scala 27:72]
  wire [21:0] _T_6402 = _T_5023 ? btb_bank0_rd_data_way1_out_157 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6657 = _T_6656 | _T_6402; // @[Mux.scala 27:72]
  wire [21:0] _T_6403 = _T_5025 ? btb_bank0_rd_data_way1_out_158 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6658 = _T_6657 | _T_6403; // @[Mux.scala 27:72]
  wire [21:0] _T_6404 = _T_5027 ? btb_bank0_rd_data_way1_out_159 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6659 = _T_6658 | _T_6404; // @[Mux.scala 27:72]
  wire [21:0] _T_6405 = _T_5029 ? btb_bank0_rd_data_way1_out_160 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6660 = _T_6659 | _T_6405; // @[Mux.scala 27:72]
  wire [21:0] _T_6406 = _T_5031 ? btb_bank0_rd_data_way1_out_161 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6661 = _T_6660 | _T_6406; // @[Mux.scala 27:72]
  wire [21:0] _T_6407 = _T_5033 ? btb_bank0_rd_data_way1_out_162 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6662 = _T_6661 | _T_6407; // @[Mux.scala 27:72]
  wire [21:0] _T_6408 = _T_5035 ? btb_bank0_rd_data_way1_out_163 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6663 = _T_6662 | _T_6408; // @[Mux.scala 27:72]
  wire [21:0] _T_6409 = _T_5037 ? btb_bank0_rd_data_way1_out_164 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6664 = _T_6663 | _T_6409; // @[Mux.scala 27:72]
  wire [21:0] _T_6410 = _T_5039 ? btb_bank0_rd_data_way1_out_165 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6665 = _T_6664 | _T_6410; // @[Mux.scala 27:72]
  wire [21:0] _T_6411 = _T_5041 ? btb_bank0_rd_data_way1_out_166 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6666 = _T_6665 | _T_6411; // @[Mux.scala 27:72]
  wire [21:0] _T_6412 = _T_5043 ? btb_bank0_rd_data_way1_out_167 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6667 = _T_6666 | _T_6412; // @[Mux.scala 27:72]
  wire [21:0] _T_6413 = _T_5045 ? btb_bank0_rd_data_way1_out_168 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6668 = _T_6667 | _T_6413; // @[Mux.scala 27:72]
  wire [21:0] _T_6414 = _T_5047 ? btb_bank0_rd_data_way1_out_169 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6669 = _T_6668 | _T_6414; // @[Mux.scala 27:72]
  wire [21:0] _T_6415 = _T_5049 ? btb_bank0_rd_data_way1_out_170 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6670 = _T_6669 | _T_6415; // @[Mux.scala 27:72]
  wire [21:0] _T_6416 = _T_5051 ? btb_bank0_rd_data_way1_out_171 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6671 = _T_6670 | _T_6416; // @[Mux.scala 27:72]
  wire [21:0] _T_6417 = _T_5053 ? btb_bank0_rd_data_way1_out_172 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6672 = _T_6671 | _T_6417; // @[Mux.scala 27:72]
  wire [21:0] _T_6418 = _T_5055 ? btb_bank0_rd_data_way1_out_173 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6673 = _T_6672 | _T_6418; // @[Mux.scala 27:72]
  wire [21:0] _T_6419 = _T_5057 ? btb_bank0_rd_data_way1_out_174 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6674 = _T_6673 | _T_6419; // @[Mux.scala 27:72]
  wire [21:0] _T_6420 = _T_5059 ? btb_bank0_rd_data_way1_out_175 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6675 = _T_6674 | _T_6420; // @[Mux.scala 27:72]
  wire [21:0] _T_6421 = _T_5061 ? btb_bank0_rd_data_way1_out_176 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6676 = _T_6675 | _T_6421; // @[Mux.scala 27:72]
  wire [21:0] _T_6422 = _T_5063 ? btb_bank0_rd_data_way1_out_177 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6677 = _T_6676 | _T_6422; // @[Mux.scala 27:72]
  wire [21:0] _T_6423 = _T_5065 ? btb_bank0_rd_data_way1_out_178 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6678 = _T_6677 | _T_6423; // @[Mux.scala 27:72]
  wire [21:0] _T_6424 = _T_5067 ? btb_bank0_rd_data_way1_out_179 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6679 = _T_6678 | _T_6424; // @[Mux.scala 27:72]
  wire [21:0] _T_6425 = _T_5069 ? btb_bank0_rd_data_way1_out_180 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6680 = _T_6679 | _T_6425; // @[Mux.scala 27:72]
  wire [21:0] _T_6426 = _T_5071 ? btb_bank0_rd_data_way1_out_181 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6681 = _T_6680 | _T_6426; // @[Mux.scala 27:72]
  wire [21:0] _T_6427 = _T_5073 ? btb_bank0_rd_data_way1_out_182 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6682 = _T_6681 | _T_6427; // @[Mux.scala 27:72]
  wire [21:0] _T_6428 = _T_5075 ? btb_bank0_rd_data_way1_out_183 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6683 = _T_6682 | _T_6428; // @[Mux.scala 27:72]
  wire [21:0] _T_6429 = _T_5077 ? btb_bank0_rd_data_way1_out_184 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6684 = _T_6683 | _T_6429; // @[Mux.scala 27:72]
  wire [21:0] _T_6430 = _T_5079 ? btb_bank0_rd_data_way1_out_185 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6685 = _T_6684 | _T_6430; // @[Mux.scala 27:72]
  wire [21:0] _T_6431 = _T_5081 ? btb_bank0_rd_data_way1_out_186 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6686 = _T_6685 | _T_6431; // @[Mux.scala 27:72]
  wire [21:0] _T_6432 = _T_5083 ? btb_bank0_rd_data_way1_out_187 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6687 = _T_6686 | _T_6432; // @[Mux.scala 27:72]
  wire [21:0] _T_6433 = _T_5085 ? btb_bank0_rd_data_way1_out_188 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6688 = _T_6687 | _T_6433; // @[Mux.scala 27:72]
  wire [21:0] _T_6434 = _T_5087 ? btb_bank0_rd_data_way1_out_189 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6689 = _T_6688 | _T_6434; // @[Mux.scala 27:72]
  wire [21:0] _T_6435 = _T_5089 ? btb_bank0_rd_data_way1_out_190 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6690 = _T_6689 | _T_6435; // @[Mux.scala 27:72]
  wire [21:0] _T_6436 = _T_5091 ? btb_bank0_rd_data_way1_out_191 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6691 = _T_6690 | _T_6436; // @[Mux.scala 27:72]
  wire [21:0] _T_6437 = _T_5093 ? btb_bank0_rd_data_way1_out_192 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6692 = _T_6691 | _T_6437; // @[Mux.scala 27:72]
  wire [21:0] _T_6438 = _T_5095 ? btb_bank0_rd_data_way1_out_193 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6693 = _T_6692 | _T_6438; // @[Mux.scala 27:72]
  wire [21:0] _T_6439 = _T_5097 ? btb_bank0_rd_data_way1_out_194 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6694 = _T_6693 | _T_6439; // @[Mux.scala 27:72]
  wire [21:0] _T_6440 = _T_5099 ? btb_bank0_rd_data_way1_out_195 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6695 = _T_6694 | _T_6440; // @[Mux.scala 27:72]
  wire [21:0] _T_6441 = _T_5101 ? btb_bank0_rd_data_way1_out_196 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6696 = _T_6695 | _T_6441; // @[Mux.scala 27:72]
  wire [21:0] _T_6442 = _T_5103 ? btb_bank0_rd_data_way1_out_197 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6697 = _T_6696 | _T_6442; // @[Mux.scala 27:72]
  wire [21:0] _T_6443 = _T_5105 ? btb_bank0_rd_data_way1_out_198 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6698 = _T_6697 | _T_6443; // @[Mux.scala 27:72]
  wire [21:0] _T_6444 = _T_5107 ? btb_bank0_rd_data_way1_out_199 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6699 = _T_6698 | _T_6444; // @[Mux.scala 27:72]
  wire [21:0] _T_6445 = _T_5109 ? btb_bank0_rd_data_way1_out_200 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6700 = _T_6699 | _T_6445; // @[Mux.scala 27:72]
  wire [21:0] _T_6446 = _T_5111 ? btb_bank0_rd_data_way1_out_201 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6701 = _T_6700 | _T_6446; // @[Mux.scala 27:72]
  wire [21:0] _T_6447 = _T_5113 ? btb_bank0_rd_data_way1_out_202 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6702 = _T_6701 | _T_6447; // @[Mux.scala 27:72]
  wire [21:0] _T_6448 = _T_5115 ? btb_bank0_rd_data_way1_out_203 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6703 = _T_6702 | _T_6448; // @[Mux.scala 27:72]
  wire [21:0] _T_6449 = _T_5117 ? btb_bank0_rd_data_way1_out_204 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6704 = _T_6703 | _T_6449; // @[Mux.scala 27:72]
  wire [21:0] _T_6450 = _T_5119 ? btb_bank0_rd_data_way1_out_205 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6705 = _T_6704 | _T_6450; // @[Mux.scala 27:72]
  wire [21:0] _T_6451 = _T_5121 ? btb_bank0_rd_data_way1_out_206 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6706 = _T_6705 | _T_6451; // @[Mux.scala 27:72]
  wire [21:0] _T_6452 = _T_5123 ? btb_bank0_rd_data_way1_out_207 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6707 = _T_6706 | _T_6452; // @[Mux.scala 27:72]
  wire [21:0] _T_6453 = _T_5125 ? btb_bank0_rd_data_way1_out_208 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6708 = _T_6707 | _T_6453; // @[Mux.scala 27:72]
  wire [21:0] _T_6454 = _T_5127 ? btb_bank0_rd_data_way1_out_209 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6709 = _T_6708 | _T_6454; // @[Mux.scala 27:72]
  wire [21:0] _T_6455 = _T_5129 ? btb_bank0_rd_data_way1_out_210 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6710 = _T_6709 | _T_6455; // @[Mux.scala 27:72]
  wire [21:0] _T_6456 = _T_5131 ? btb_bank0_rd_data_way1_out_211 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6711 = _T_6710 | _T_6456; // @[Mux.scala 27:72]
  wire [21:0] _T_6457 = _T_5133 ? btb_bank0_rd_data_way1_out_212 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6712 = _T_6711 | _T_6457; // @[Mux.scala 27:72]
  wire [21:0] _T_6458 = _T_5135 ? btb_bank0_rd_data_way1_out_213 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6713 = _T_6712 | _T_6458; // @[Mux.scala 27:72]
  wire [21:0] _T_6459 = _T_5137 ? btb_bank0_rd_data_way1_out_214 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6714 = _T_6713 | _T_6459; // @[Mux.scala 27:72]
  wire [21:0] _T_6460 = _T_5139 ? btb_bank0_rd_data_way1_out_215 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6715 = _T_6714 | _T_6460; // @[Mux.scala 27:72]
  wire [21:0] _T_6461 = _T_5141 ? btb_bank0_rd_data_way1_out_216 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6716 = _T_6715 | _T_6461; // @[Mux.scala 27:72]
  wire [21:0] _T_6462 = _T_5143 ? btb_bank0_rd_data_way1_out_217 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6717 = _T_6716 | _T_6462; // @[Mux.scala 27:72]
  wire [21:0] _T_6463 = _T_5145 ? btb_bank0_rd_data_way1_out_218 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6718 = _T_6717 | _T_6463; // @[Mux.scala 27:72]
  wire [21:0] _T_6464 = _T_5147 ? btb_bank0_rd_data_way1_out_219 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6719 = _T_6718 | _T_6464; // @[Mux.scala 27:72]
  wire [21:0] _T_6465 = _T_5149 ? btb_bank0_rd_data_way1_out_220 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6720 = _T_6719 | _T_6465; // @[Mux.scala 27:72]
  wire [21:0] _T_6466 = _T_5151 ? btb_bank0_rd_data_way1_out_221 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6721 = _T_6720 | _T_6466; // @[Mux.scala 27:72]
  wire [21:0] _T_6467 = _T_5153 ? btb_bank0_rd_data_way1_out_222 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6722 = _T_6721 | _T_6467; // @[Mux.scala 27:72]
  wire [21:0] _T_6468 = _T_5155 ? btb_bank0_rd_data_way1_out_223 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6723 = _T_6722 | _T_6468; // @[Mux.scala 27:72]
  wire [21:0] _T_6469 = _T_5157 ? btb_bank0_rd_data_way1_out_224 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6724 = _T_6723 | _T_6469; // @[Mux.scala 27:72]
  wire [21:0] _T_6470 = _T_5159 ? btb_bank0_rd_data_way1_out_225 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6725 = _T_6724 | _T_6470; // @[Mux.scala 27:72]
  wire [21:0] _T_6471 = _T_5161 ? btb_bank0_rd_data_way1_out_226 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6726 = _T_6725 | _T_6471; // @[Mux.scala 27:72]
  wire [21:0] _T_6472 = _T_5163 ? btb_bank0_rd_data_way1_out_227 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6727 = _T_6726 | _T_6472; // @[Mux.scala 27:72]
  wire [21:0] _T_6473 = _T_5165 ? btb_bank0_rd_data_way1_out_228 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6728 = _T_6727 | _T_6473; // @[Mux.scala 27:72]
  wire [21:0] _T_6474 = _T_5167 ? btb_bank0_rd_data_way1_out_229 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6729 = _T_6728 | _T_6474; // @[Mux.scala 27:72]
  wire [21:0] _T_6475 = _T_5169 ? btb_bank0_rd_data_way1_out_230 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6730 = _T_6729 | _T_6475; // @[Mux.scala 27:72]
  wire [21:0] _T_6476 = _T_5171 ? btb_bank0_rd_data_way1_out_231 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6731 = _T_6730 | _T_6476; // @[Mux.scala 27:72]
  wire [21:0] _T_6477 = _T_5173 ? btb_bank0_rd_data_way1_out_232 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6732 = _T_6731 | _T_6477; // @[Mux.scala 27:72]
  wire [21:0] _T_6478 = _T_5175 ? btb_bank0_rd_data_way1_out_233 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6733 = _T_6732 | _T_6478; // @[Mux.scala 27:72]
  wire [21:0] _T_6479 = _T_5177 ? btb_bank0_rd_data_way1_out_234 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6734 = _T_6733 | _T_6479; // @[Mux.scala 27:72]
  wire [21:0] _T_6480 = _T_5179 ? btb_bank0_rd_data_way1_out_235 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6735 = _T_6734 | _T_6480; // @[Mux.scala 27:72]
  wire [21:0] _T_6481 = _T_5181 ? btb_bank0_rd_data_way1_out_236 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6736 = _T_6735 | _T_6481; // @[Mux.scala 27:72]
  wire [21:0] _T_6482 = _T_5183 ? btb_bank0_rd_data_way1_out_237 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6737 = _T_6736 | _T_6482; // @[Mux.scala 27:72]
  wire [21:0] _T_6483 = _T_5185 ? btb_bank0_rd_data_way1_out_238 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6738 = _T_6737 | _T_6483; // @[Mux.scala 27:72]
  wire [21:0] _T_6484 = _T_5187 ? btb_bank0_rd_data_way1_out_239 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6739 = _T_6738 | _T_6484; // @[Mux.scala 27:72]
  wire [21:0] _T_6485 = _T_5189 ? btb_bank0_rd_data_way1_out_240 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6740 = _T_6739 | _T_6485; // @[Mux.scala 27:72]
  wire [21:0] _T_6486 = _T_5191 ? btb_bank0_rd_data_way1_out_241 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6741 = _T_6740 | _T_6486; // @[Mux.scala 27:72]
  wire [21:0] _T_6487 = _T_5193 ? btb_bank0_rd_data_way1_out_242 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6742 = _T_6741 | _T_6487; // @[Mux.scala 27:72]
  wire [21:0] _T_6488 = _T_5195 ? btb_bank0_rd_data_way1_out_243 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6743 = _T_6742 | _T_6488; // @[Mux.scala 27:72]
  wire [21:0] _T_6489 = _T_5197 ? btb_bank0_rd_data_way1_out_244 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6744 = _T_6743 | _T_6489; // @[Mux.scala 27:72]
  wire [21:0] _T_6490 = _T_5199 ? btb_bank0_rd_data_way1_out_245 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6745 = _T_6744 | _T_6490; // @[Mux.scala 27:72]
  wire [21:0] _T_6491 = _T_5201 ? btb_bank0_rd_data_way1_out_246 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6746 = _T_6745 | _T_6491; // @[Mux.scala 27:72]
  wire [21:0] _T_6492 = _T_5203 ? btb_bank0_rd_data_way1_out_247 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6747 = _T_6746 | _T_6492; // @[Mux.scala 27:72]
  wire [21:0] _T_6493 = _T_5205 ? btb_bank0_rd_data_way1_out_248 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6748 = _T_6747 | _T_6493; // @[Mux.scala 27:72]
  wire [21:0] _T_6494 = _T_5207 ? btb_bank0_rd_data_way1_out_249 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6749 = _T_6748 | _T_6494; // @[Mux.scala 27:72]
  wire [21:0] _T_6495 = _T_5209 ? btb_bank0_rd_data_way1_out_250 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6750 = _T_6749 | _T_6495; // @[Mux.scala 27:72]
  wire [21:0] _T_6496 = _T_5211 ? btb_bank0_rd_data_way1_out_251 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6751 = _T_6750 | _T_6496; // @[Mux.scala 27:72]
  wire [21:0] _T_6497 = _T_5213 ? btb_bank0_rd_data_way1_out_252 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6752 = _T_6751 | _T_6497; // @[Mux.scala 27:72]
  wire [21:0] _T_6498 = _T_5215 ? btb_bank0_rd_data_way1_out_253 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6753 = _T_6752 | _T_6498; // @[Mux.scala 27:72]
  wire [21:0] _T_6499 = _T_5217 ? btb_bank0_rd_data_way1_out_254 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_6754 = _T_6753 | _T_6499; // @[Mux.scala 27:72]
  wire [21:0] _T_6500 = _T_5219 ? btb_bank0_rd_data_way1_out_255 : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0_rd_data_way1_p1_f = _T_6754 | _T_6500; // @[Mux.scala 27:72]
  wire  _T_73 = btb_bank0_rd_data_way1_p1_f[21:17] == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 155:107]
  wire  _T_74 = btb_bank0_rd_data_way1_p1_f[0] & _T_73; // @[ifu_bp_ctl.scala 155:61]
  wire  _T_77 = _T_74 & _T_67; // @[ifu_bp_ctl.scala 155:130]
  wire  _T_78 = _T_77 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 156:57]
  wire  tag_match_way1_p1_f = _T_78 & _T; // @[ifu_bp_ctl.scala 156:78]
  wire  _T_109 = btb_bank0_rd_data_way1_p1_f[3] ^ btb_bank0_rd_data_way1_p1_f[4]; // @[ifu_bp_ctl.scala 168:99]
  wire  _T_110 = tag_match_way1_p1_f & _T_109; // @[ifu_bp_ctl.scala 168:62]
  wire  _T_114 = ~_T_109; // @[ifu_bp_ctl.scala 169:27]
  wire  _T_115 = tag_match_way1_p1_f & _T_114; // @[ifu_bp_ctl.scala 169:25]
  wire [1:0] tag_match_way1_expanded_p1_f = {_T_110,_T_115}; // @[Cat.scala 29:58]
  wire [21:0] _T_137 = tag_match_way1_expanded_p1_f[0] ? btb_bank0_rd_data_way1_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_p1_f = _T_136 | _T_137; // @[Mux.scala 27:72]
  wire [21:0] _T_150 = io_ifc_fetch_addr_f[0] ? btb_bank0e_rd_data_p1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank1_rd_data_f = _T_149 | _T_150; // @[Mux.scala 27:72]
  wire  _T_236 = btb_vbank1_rd_data_f[2] | btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 280:59]
  wire [21:0] _T_122 = tag_match_way0_expanded_f[0] ? btb_bank0_rd_data_way0_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_123 = tag_match_way1_expanded_f[0] ? btb_bank0_rd_data_way1_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_bank0e_rd_data_f = _T_122 | _T_123; // @[Mux.scala 27:72]
  wire [21:0] _T_142 = _T_147 ? btb_bank0e_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] _T_143 = io_ifc_fetch_addr_f[0] ? btb_bank0o_rd_data_f : 22'h0; // @[Mux.scala 27:72]
  wire [21:0] btb_vbank0_rd_data_f = _T_142 | _T_143; // @[Mux.scala 27:72]
  wire  _T_239 = btb_vbank0_rd_data_f[2] | btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 281:59]
  wire [1:0] bht_force_taken_f = {_T_236,_T_239}; // @[Cat.scala 29:58]
  wire [9:0] _T_582 = {btb_rd_addr_f,2'h0}; // @[Cat.scala 29:58]
  reg [7:0] fghr; // @[Reg.scala 27:20]
  wire [7:0] bht_rd_addr_hashed_f = _T_582[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_22469 = bht_rd_addr_hashed_f == 8'h0; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_0; // @[Reg.scala 27:20]
  wire [1:0] _T_22981 = _T_22469 ? bht_bank_rd_data_out_1_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_22471 = bht_rd_addr_hashed_f == 8'h1; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_1; // @[Reg.scala 27:20]
  wire [1:0] _T_22982 = _T_22471 ? bht_bank_rd_data_out_1_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23237 = _T_22981 | _T_22982; // @[Mux.scala 27:72]
  wire  _T_22473 = bht_rd_addr_hashed_f == 8'h2; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_2; // @[Reg.scala 27:20]
  wire [1:0] _T_22983 = _T_22473 ? bht_bank_rd_data_out_1_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23238 = _T_23237 | _T_22983; // @[Mux.scala 27:72]
  wire  _T_22475 = bht_rd_addr_hashed_f == 8'h3; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_3; // @[Reg.scala 27:20]
  wire [1:0] _T_22984 = _T_22475 ? bht_bank_rd_data_out_1_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23239 = _T_23238 | _T_22984; // @[Mux.scala 27:72]
  wire  _T_22477 = bht_rd_addr_hashed_f == 8'h4; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_4; // @[Reg.scala 27:20]
  wire [1:0] _T_22985 = _T_22477 ? bht_bank_rd_data_out_1_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23240 = _T_23239 | _T_22985; // @[Mux.scala 27:72]
  wire  _T_22479 = bht_rd_addr_hashed_f == 8'h5; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_5; // @[Reg.scala 27:20]
  wire [1:0] _T_22986 = _T_22479 ? bht_bank_rd_data_out_1_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23241 = _T_23240 | _T_22986; // @[Mux.scala 27:72]
  wire  _T_22481 = bht_rd_addr_hashed_f == 8'h6; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_6; // @[Reg.scala 27:20]
  wire [1:0] _T_22987 = _T_22481 ? bht_bank_rd_data_out_1_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23242 = _T_23241 | _T_22987; // @[Mux.scala 27:72]
  wire  _T_22483 = bht_rd_addr_hashed_f == 8'h7; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_7; // @[Reg.scala 27:20]
  wire [1:0] _T_22988 = _T_22483 ? bht_bank_rd_data_out_1_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23243 = _T_23242 | _T_22988; // @[Mux.scala 27:72]
  wire  _T_22485 = bht_rd_addr_hashed_f == 8'h8; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_8; // @[Reg.scala 27:20]
  wire [1:0] _T_22989 = _T_22485 ? bht_bank_rd_data_out_1_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23244 = _T_23243 | _T_22989; // @[Mux.scala 27:72]
  wire  _T_22487 = bht_rd_addr_hashed_f == 8'h9; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_9; // @[Reg.scala 27:20]
  wire [1:0] _T_22990 = _T_22487 ? bht_bank_rd_data_out_1_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23245 = _T_23244 | _T_22990; // @[Mux.scala 27:72]
  wire  _T_22489 = bht_rd_addr_hashed_f == 8'ha; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_10; // @[Reg.scala 27:20]
  wire [1:0] _T_22991 = _T_22489 ? bht_bank_rd_data_out_1_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23246 = _T_23245 | _T_22991; // @[Mux.scala 27:72]
  wire  _T_22491 = bht_rd_addr_hashed_f == 8'hb; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_11; // @[Reg.scala 27:20]
  wire [1:0] _T_22992 = _T_22491 ? bht_bank_rd_data_out_1_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23247 = _T_23246 | _T_22992; // @[Mux.scala 27:72]
  wire  _T_22493 = bht_rd_addr_hashed_f == 8'hc; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_12; // @[Reg.scala 27:20]
  wire [1:0] _T_22993 = _T_22493 ? bht_bank_rd_data_out_1_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23248 = _T_23247 | _T_22993; // @[Mux.scala 27:72]
  wire  _T_22495 = bht_rd_addr_hashed_f == 8'hd; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_13; // @[Reg.scala 27:20]
  wire [1:0] _T_22994 = _T_22495 ? bht_bank_rd_data_out_1_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23249 = _T_23248 | _T_22994; // @[Mux.scala 27:72]
  wire  _T_22497 = bht_rd_addr_hashed_f == 8'he; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_14; // @[Reg.scala 27:20]
  wire [1:0] _T_22995 = _T_22497 ? bht_bank_rd_data_out_1_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23250 = _T_23249 | _T_22995; // @[Mux.scala 27:72]
  wire  _T_22499 = bht_rd_addr_hashed_f == 8'hf; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_15; // @[Reg.scala 27:20]
  wire [1:0] _T_22996 = _T_22499 ? bht_bank_rd_data_out_1_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23251 = _T_23250 | _T_22996; // @[Mux.scala 27:72]
  wire  _T_22501 = bht_rd_addr_hashed_f == 8'h10; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_16; // @[Reg.scala 27:20]
  wire [1:0] _T_22997 = _T_22501 ? bht_bank_rd_data_out_1_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23252 = _T_23251 | _T_22997; // @[Mux.scala 27:72]
  wire  _T_22503 = bht_rd_addr_hashed_f == 8'h11; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_17; // @[Reg.scala 27:20]
  wire [1:0] _T_22998 = _T_22503 ? bht_bank_rd_data_out_1_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23253 = _T_23252 | _T_22998; // @[Mux.scala 27:72]
  wire  _T_22505 = bht_rd_addr_hashed_f == 8'h12; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_18; // @[Reg.scala 27:20]
  wire [1:0] _T_22999 = _T_22505 ? bht_bank_rd_data_out_1_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23254 = _T_23253 | _T_22999; // @[Mux.scala 27:72]
  wire  _T_22507 = bht_rd_addr_hashed_f == 8'h13; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_19; // @[Reg.scala 27:20]
  wire [1:0] _T_23000 = _T_22507 ? bht_bank_rd_data_out_1_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23255 = _T_23254 | _T_23000; // @[Mux.scala 27:72]
  wire  _T_22509 = bht_rd_addr_hashed_f == 8'h14; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_20; // @[Reg.scala 27:20]
  wire [1:0] _T_23001 = _T_22509 ? bht_bank_rd_data_out_1_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23256 = _T_23255 | _T_23001; // @[Mux.scala 27:72]
  wire  _T_22511 = bht_rd_addr_hashed_f == 8'h15; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_21; // @[Reg.scala 27:20]
  wire [1:0] _T_23002 = _T_22511 ? bht_bank_rd_data_out_1_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23257 = _T_23256 | _T_23002; // @[Mux.scala 27:72]
  wire  _T_22513 = bht_rd_addr_hashed_f == 8'h16; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_22; // @[Reg.scala 27:20]
  wire [1:0] _T_23003 = _T_22513 ? bht_bank_rd_data_out_1_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23258 = _T_23257 | _T_23003; // @[Mux.scala 27:72]
  wire  _T_22515 = bht_rd_addr_hashed_f == 8'h17; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_23; // @[Reg.scala 27:20]
  wire [1:0] _T_23004 = _T_22515 ? bht_bank_rd_data_out_1_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23259 = _T_23258 | _T_23004; // @[Mux.scala 27:72]
  wire  _T_22517 = bht_rd_addr_hashed_f == 8'h18; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_24; // @[Reg.scala 27:20]
  wire [1:0] _T_23005 = _T_22517 ? bht_bank_rd_data_out_1_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23260 = _T_23259 | _T_23005; // @[Mux.scala 27:72]
  wire  _T_22519 = bht_rd_addr_hashed_f == 8'h19; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_25; // @[Reg.scala 27:20]
  wire [1:0] _T_23006 = _T_22519 ? bht_bank_rd_data_out_1_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23261 = _T_23260 | _T_23006; // @[Mux.scala 27:72]
  wire  _T_22521 = bht_rd_addr_hashed_f == 8'h1a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_26; // @[Reg.scala 27:20]
  wire [1:0] _T_23007 = _T_22521 ? bht_bank_rd_data_out_1_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23262 = _T_23261 | _T_23007; // @[Mux.scala 27:72]
  wire  _T_22523 = bht_rd_addr_hashed_f == 8'h1b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_27; // @[Reg.scala 27:20]
  wire [1:0] _T_23008 = _T_22523 ? bht_bank_rd_data_out_1_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23263 = _T_23262 | _T_23008; // @[Mux.scala 27:72]
  wire  _T_22525 = bht_rd_addr_hashed_f == 8'h1c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_28; // @[Reg.scala 27:20]
  wire [1:0] _T_23009 = _T_22525 ? bht_bank_rd_data_out_1_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23264 = _T_23263 | _T_23009; // @[Mux.scala 27:72]
  wire  _T_22527 = bht_rd_addr_hashed_f == 8'h1d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_29; // @[Reg.scala 27:20]
  wire [1:0] _T_23010 = _T_22527 ? bht_bank_rd_data_out_1_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23265 = _T_23264 | _T_23010; // @[Mux.scala 27:72]
  wire  _T_22529 = bht_rd_addr_hashed_f == 8'h1e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_30; // @[Reg.scala 27:20]
  wire [1:0] _T_23011 = _T_22529 ? bht_bank_rd_data_out_1_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23266 = _T_23265 | _T_23011; // @[Mux.scala 27:72]
  wire  _T_22531 = bht_rd_addr_hashed_f == 8'h1f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_31; // @[Reg.scala 27:20]
  wire [1:0] _T_23012 = _T_22531 ? bht_bank_rd_data_out_1_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23267 = _T_23266 | _T_23012; // @[Mux.scala 27:72]
  wire  _T_22533 = bht_rd_addr_hashed_f == 8'h20; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_32; // @[Reg.scala 27:20]
  wire [1:0] _T_23013 = _T_22533 ? bht_bank_rd_data_out_1_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23268 = _T_23267 | _T_23013; // @[Mux.scala 27:72]
  wire  _T_22535 = bht_rd_addr_hashed_f == 8'h21; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_33; // @[Reg.scala 27:20]
  wire [1:0] _T_23014 = _T_22535 ? bht_bank_rd_data_out_1_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23269 = _T_23268 | _T_23014; // @[Mux.scala 27:72]
  wire  _T_22537 = bht_rd_addr_hashed_f == 8'h22; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_34; // @[Reg.scala 27:20]
  wire [1:0] _T_23015 = _T_22537 ? bht_bank_rd_data_out_1_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23270 = _T_23269 | _T_23015; // @[Mux.scala 27:72]
  wire  _T_22539 = bht_rd_addr_hashed_f == 8'h23; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_35; // @[Reg.scala 27:20]
  wire [1:0] _T_23016 = _T_22539 ? bht_bank_rd_data_out_1_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23271 = _T_23270 | _T_23016; // @[Mux.scala 27:72]
  wire  _T_22541 = bht_rd_addr_hashed_f == 8'h24; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_36; // @[Reg.scala 27:20]
  wire [1:0] _T_23017 = _T_22541 ? bht_bank_rd_data_out_1_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23272 = _T_23271 | _T_23017; // @[Mux.scala 27:72]
  wire  _T_22543 = bht_rd_addr_hashed_f == 8'h25; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_37; // @[Reg.scala 27:20]
  wire [1:0] _T_23018 = _T_22543 ? bht_bank_rd_data_out_1_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23273 = _T_23272 | _T_23018; // @[Mux.scala 27:72]
  wire  _T_22545 = bht_rd_addr_hashed_f == 8'h26; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_38; // @[Reg.scala 27:20]
  wire [1:0] _T_23019 = _T_22545 ? bht_bank_rd_data_out_1_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23274 = _T_23273 | _T_23019; // @[Mux.scala 27:72]
  wire  _T_22547 = bht_rd_addr_hashed_f == 8'h27; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_39; // @[Reg.scala 27:20]
  wire [1:0] _T_23020 = _T_22547 ? bht_bank_rd_data_out_1_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23275 = _T_23274 | _T_23020; // @[Mux.scala 27:72]
  wire  _T_22549 = bht_rd_addr_hashed_f == 8'h28; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_40; // @[Reg.scala 27:20]
  wire [1:0] _T_23021 = _T_22549 ? bht_bank_rd_data_out_1_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23276 = _T_23275 | _T_23021; // @[Mux.scala 27:72]
  wire  _T_22551 = bht_rd_addr_hashed_f == 8'h29; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_41; // @[Reg.scala 27:20]
  wire [1:0] _T_23022 = _T_22551 ? bht_bank_rd_data_out_1_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23277 = _T_23276 | _T_23022; // @[Mux.scala 27:72]
  wire  _T_22553 = bht_rd_addr_hashed_f == 8'h2a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_42; // @[Reg.scala 27:20]
  wire [1:0] _T_23023 = _T_22553 ? bht_bank_rd_data_out_1_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23278 = _T_23277 | _T_23023; // @[Mux.scala 27:72]
  wire  _T_22555 = bht_rd_addr_hashed_f == 8'h2b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_43; // @[Reg.scala 27:20]
  wire [1:0] _T_23024 = _T_22555 ? bht_bank_rd_data_out_1_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23279 = _T_23278 | _T_23024; // @[Mux.scala 27:72]
  wire  _T_22557 = bht_rd_addr_hashed_f == 8'h2c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_44; // @[Reg.scala 27:20]
  wire [1:0] _T_23025 = _T_22557 ? bht_bank_rd_data_out_1_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23280 = _T_23279 | _T_23025; // @[Mux.scala 27:72]
  wire  _T_22559 = bht_rd_addr_hashed_f == 8'h2d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_45; // @[Reg.scala 27:20]
  wire [1:0] _T_23026 = _T_22559 ? bht_bank_rd_data_out_1_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23281 = _T_23280 | _T_23026; // @[Mux.scala 27:72]
  wire  _T_22561 = bht_rd_addr_hashed_f == 8'h2e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_46; // @[Reg.scala 27:20]
  wire [1:0] _T_23027 = _T_22561 ? bht_bank_rd_data_out_1_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23282 = _T_23281 | _T_23027; // @[Mux.scala 27:72]
  wire  _T_22563 = bht_rd_addr_hashed_f == 8'h2f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_47; // @[Reg.scala 27:20]
  wire [1:0] _T_23028 = _T_22563 ? bht_bank_rd_data_out_1_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23283 = _T_23282 | _T_23028; // @[Mux.scala 27:72]
  wire  _T_22565 = bht_rd_addr_hashed_f == 8'h30; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_48; // @[Reg.scala 27:20]
  wire [1:0] _T_23029 = _T_22565 ? bht_bank_rd_data_out_1_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23284 = _T_23283 | _T_23029; // @[Mux.scala 27:72]
  wire  _T_22567 = bht_rd_addr_hashed_f == 8'h31; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_49; // @[Reg.scala 27:20]
  wire [1:0] _T_23030 = _T_22567 ? bht_bank_rd_data_out_1_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23285 = _T_23284 | _T_23030; // @[Mux.scala 27:72]
  wire  _T_22569 = bht_rd_addr_hashed_f == 8'h32; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_50; // @[Reg.scala 27:20]
  wire [1:0] _T_23031 = _T_22569 ? bht_bank_rd_data_out_1_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23286 = _T_23285 | _T_23031; // @[Mux.scala 27:72]
  wire  _T_22571 = bht_rd_addr_hashed_f == 8'h33; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_51; // @[Reg.scala 27:20]
  wire [1:0] _T_23032 = _T_22571 ? bht_bank_rd_data_out_1_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23287 = _T_23286 | _T_23032; // @[Mux.scala 27:72]
  wire  _T_22573 = bht_rd_addr_hashed_f == 8'h34; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_52; // @[Reg.scala 27:20]
  wire [1:0] _T_23033 = _T_22573 ? bht_bank_rd_data_out_1_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23288 = _T_23287 | _T_23033; // @[Mux.scala 27:72]
  wire  _T_22575 = bht_rd_addr_hashed_f == 8'h35; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_53; // @[Reg.scala 27:20]
  wire [1:0] _T_23034 = _T_22575 ? bht_bank_rd_data_out_1_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23289 = _T_23288 | _T_23034; // @[Mux.scala 27:72]
  wire  _T_22577 = bht_rd_addr_hashed_f == 8'h36; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_54; // @[Reg.scala 27:20]
  wire [1:0] _T_23035 = _T_22577 ? bht_bank_rd_data_out_1_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23290 = _T_23289 | _T_23035; // @[Mux.scala 27:72]
  wire  _T_22579 = bht_rd_addr_hashed_f == 8'h37; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_55; // @[Reg.scala 27:20]
  wire [1:0] _T_23036 = _T_22579 ? bht_bank_rd_data_out_1_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23291 = _T_23290 | _T_23036; // @[Mux.scala 27:72]
  wire  _T_22581 = bht_rd_addr_hashed_f == 8'h38; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_56; // @[Reg.scala 27:20]
  wire [1:0] _T_23037 = _T_22581 ? bht_bank_rd_data_out_1_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23292 = _T_23291 | _T_23037; // @[Mux.scala 27:72]
  wire  _T_22583 = bht_rd_addr_hashed_f == 8'h39; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_57; // @[Reg.scala 27:20]
  wire [1:0] _T_23038 = _T_22583 ? bht_bank_rd_data_out_1_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23293 = _T_23292 | _T_23038; // @[Mux.scala 27:72]
  wire  _T_22585 = bht_rd_addr_hashed_f == 8'h3a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_58; // @[Reg.scala 27:20]
  wire [1:0] _T_23039 = _T_22585 ? bht_bank_rd_data_out_1_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23294 = _T_23293 | _T_23039; // @[Mux.scala 27:72]
  wire  _T_22587 = bht_rd_addr_hashed_f == 8'h3b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_59; // @[Reg.scala 27:20]
  wire [1:0] _T_23040 = _T_22587 ? bht_bank_rd_data_out_1_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23295 = _T_23294 | _T_23040; // @[Mux.scala 27:72]
  wire  _T_22589 = bht_rd_addr_hashed_f == 8'h3c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_60; // @[Reg.scala 27:20]
  wire [1:0] _T_23041 = _T_22589 ? bht_bank_rd_data_out_1_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23296 = _T_23295 | _T_23041; // @[Mux.scala 27:72]
  wire  _T_22591 = bht_rd_addr_hashed_f == 8'h3d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_61; // @[Reg.scala 27:20]
  wire [1:0] _T_23042 = _T_22591 ? bht_bank_rd_data_out_1_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23297 = _T_23296 | _T_23042; // @[Mux.scala 27:72]
  wire  _T_22593 = bht_rd_addr_hashed_f == 8'h3e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_62; // @[Reg.scala 27:20]
  wire [1:0] _T_23043 = _T_22593 ? bht_bank_rd_data_out_1_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23298 = _T_23297 | _T_23043; // @[Mux.scala 27:72]
  wire  _T_22595 = bht_rd_addr_hashed_f == 8'h3f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_63; // @[Reg.scala 27:20]
  wire [1:0] _T_23044 = _T_22595 ? bht_bank_rd_data_out_1_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23299 = _T_23298 | _T_23044; // @[Mux.scala 27:72]
  wire  _T_22597 = bht_rd_addr_hashed_f == 8'h40; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_64; // @[Reg.scala 27:20]
  wire [1:0] _T_23045 = _T_22597 ? bht_bank_rd_data_out_1_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23300 = _T_23299 | _T_23045; // @[Mux.scala 27:72]
  wire  _T_22599 = bht_rd_addr_hashed_f == 8'h41; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_65; // @[Reg.scala 27:20]
  wire [1:0] _T_23046 = _T_22599 ? bht_bank_rd_data_out_1_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23301 = _T_23300 | _T_23046; // @[Mux.scala 27:72]
  wire  _T_22601 = bht_rd_addr_hashed_f == 8'h42; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_66; // @[Reg.scala 27:20]
  wire [1:0] _T_23047 = _T_22601 ? bht_bank_rd_data_out_1_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23302 = _T_23301 | _T_23047; // @[Mux.scala 27:72]
  wire  _T_22603 = bht_rd_addr_hashed_f == 8'h43; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_67; // @[Reg.scala 27:20]
  wire [1:0] _T_23048 = _T_22603 ? bht_bank_rd_data_out_1_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23303 = _T_23302 | _T_23048; // @[Mux.scala 27:72]
  wire  _T_22605 = bht_rd_addr_hashed_f == 8'h44; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_68; // @[Reg.scala 27:20]
  wire [1:0] _T_23049 = _T_22605 ? bht_bank_rd_data_out_1_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23304 = _T_23303 | _T_23049; // @[Mux.scala 27:72]
  wire  _T_22607 = bht_rd_addr_hashed_f == 8'h45; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_69; // @[Reg.scala 27:20]
  wire [1:0] _T_23050 = _T_22607 ? bht_bank_rd_data_out_1_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23305 = _T_23304 | _T_23050; // @[Mux.scala 27:72]
  wire  _T_22609 = bht_rd_addr_hashed_f == 8'h46; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_70; // @[Reg.scala 27:20]
  wire [1:0] _T_23051 = _T_22609 ? bht_bank_rd_data_out_1_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23306 = _T_23305 | _T_23051; // @[Mux.scala 27:72]
  wire  _T_22611 = bht_rd_addr_hashed_f == 8'h47; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_71; // @[Reg.scala 27:20]
  wire [1:0] _T_23052 = _T_22611 ? bht_bank_rd_data_out_1_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23307 = _T_23306 | _T_23052; // @[Mux.scala 27:72]
  wire  _T_22613 = bht_rd_addr_hashed_f == 8'h48; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_72; // @[Reg.scala 27:20]
  wire [1:0] _T_23053 = _T_22613 ? bht_bank_rd_data_out_1_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23308 = _T_23307 | _T_23053; // @[Mux.scala 27:72]
  wire  _T_22615 = bht_rd_addr_hashed_f == 8'h49; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_73; // @[Reg.scala 27:20]
  wire [1:0] _T_23054 = _T_22615 ? bht_bank_rd_data_out_1_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23309 = _T_23308 | _T_23054; // @[Mux.scala 27:72]
  wire  _T_22617 = bht_rd_addr_hashed_f == 8'h4a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_74; // @[Reg.scala 27:20]
  wire [1:0] _T_23055 = _T_22617 ? bht_bank_rd_data_out_1_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23310 = _T_23309 | _T_23055; // @[Mux.scala 27:72]
  wire  _T_22619 = bht_rd_addr_hashed_f == 8'h4b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_75; // @[Reg.scala 27:20]
  wire [1:0] _T_23056 = _T_22619 ? bht_bank_rd_data_out_1_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23311 = _T_23310 | _T_23056; // @[Mux.scala 27:72]
  wire  _T_22621 = bht_rd_addr_hashed_f == 8'h4c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_76; // @[Reg.scala 27:20]
  wire [1:0] _T_23057 = _T_22621 ? bht_bank_rd_data_out_1_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23312 = _T_23311 | _T_23057; // @[Mux.scala 27:72]
  wire  _T_22623 = bht_rd_addr_hashed_f == 8'h4d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_77; // @[Reg.scala 27:20]
  wire [1:0] _T_23058 = _T_22623 ? bht_bank_rd_data_out_1_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23313 = _T_23312 | _T_23058; // @[Mux.scala 27:72]
  wire  _T_22625 = bht_rd_addr_hashed_f == 8'h4e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_78; // @[Reg.scala 27:20]
  wire [1:0] _T_23059 = _T_22625 ? bht_bank_rd_data_out_1_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23314 = _T_23313 | _T_23059; // @[Mux.scala 27:72]
  wire  _T_22627 = bht_rd_addr_hashed_f == 8'h4f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_79; // @[Reg.scala 27:20]
  wire [1:0] _T_23060 = _T_22627 ? bht_bank_rd_data_out_1_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23315 = _T_23314 | _T_23060; // @[Mux.scala 27:72]
  wire  _T_22629 = bht_rd_addr_hashed_f == 8'h50; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_80; // @[Reg.scala 27:20]
  wire [1:0] _T_23061 = _T_22629 ? bht_bank_rd_data_out_1_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23316 = _T_23315 | _T_23061; // @[Mux.scala 27:72]
  wire  _T_22631 = bht_rd_addr_hashed_f == 8'h51; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_81; // @[Reg.scala 27:20]
  wire [1:0] _T_23062 = _T_22631 ? bht_bank_rd_data_out_1_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23317 = _T_23316 | _T_23062; // @[Mux.scala 27:72]
  wire  _T_22633 = bht_rd_addr_hashed_f == 8'h52; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_82; // @[Reg.scala 27:20]
  wire [1:0] _T_23063 = _T_22633 ? bht_bank_rd_data_out_1_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23318 = _T_23317 | _T_23063; // @[Mux.scala 27:72]
  wire  _T_22635 = bht_rd_addr_hashed_f == 8'h53; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_83; // @[Reg.scala 27:20]
  wire [1:0] _T_23064 = _T_22635 ? bht_bank_rd_data_out_1_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23319 = _T_23318 | _T_23064; // @[Mux.scala 27:72]
  wire  _T_22637 = bht_rd_addr_hashed_f == 8'h54; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_84; // @[Reg.scala 27:20]
  wire [1:0] _T_23065 = _T_22637 ? bht_bank_rd_data_out_1_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23320 = _T_23319 | _T_23065; // @[Mux.scala 27:72]
  wire  _T_22639 = bht_rd_addr_hashed_f == 8'h55; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_85; // @[Reg.scala 27:20]
  wire [1:0] _T_23066 = _T_22639 ? bht_bank_rd_data_out_1_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23321 = _T_23320 | _T_23066; // @[Mux.scala 27:72]
  wire  _T_22641 = bht_rd_addr_hashed_f == 8'h56; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_86; // @[Reg.scala 27:20]
  wire [1:0] _T_23067 = _T_22641 ? bht_bank_rd_data_out_1_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23322 = _T_23321 | _T_23067; // @[Mux.scala 27:72]
  wire  _T_22643 = bht_rd_addr_hashed_f == 8'h57; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_87; // @[Reg.scala 27:20]
  wire [1:0] _T_23068 = _T_22643 ? bht_bank_rd_data_out_1_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23323 = _T_23322 | _T_23068; // @[Mux.scala 27:72]
  wire  _T_22645 = bht_rd_addr_hashed_f == 8'h58; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_88; // @[Reg.scala 27:20]
  wire [1:0] _T_23069 = _T_22645 ? bht_bank_rd_data_out_1_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23324 = _T_23323 | _T_23069; // @[Mux.scala 27:72]
  wire  _T_22647 = bht_rd_addr_hashed_f == 8'h59; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_89; // @[Reg.scala 27:20]
  wire [1:0] _T_23070 = _T_22647 ? bht_bank_rd_data_out_1_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23325 = _T_23324 | _T_23070; // @[Mux.scala 27:72]
  wire  _T_22649 = bht_rd_addr_hashed_f == 8'h5a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_90; // @[Reg.scala 27:20]
  wire [1:0] _T_23071 = _T_22649 ? bht_bank_rd_data_out_1_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23326 = _T_23325 | _T_23071; // @[Mux.scala 27:72]
  wire  _T_22651 = bht_rd_addr_hashed_f == 8'h5b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_91; // @[Reg.scala 27:20]
  wire [1:0] _T_23072 = _T_22651 ? bht_bank_rd_data_out_1_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23327 = _T_23326 | _T_23072; // @[Mux.scala 27:72]
  wire  _T_22653 = bht_rd_addr_hashed_f == 8'h5c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_92; // @[Reg.scala 27:20]
  wire [1:0] _T_23073 = _T_22653 ? bht_bank_rd_data_out_1_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23328 = _T_23327 | _T_23073; // @[Mux.scala 27:72]
  wire  _T_22655 = bht_rd_addr_hashed_f == 8'h5d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_93; // @[Reg.scala 27:20]
  wire [1:0] _T_23074 = _T_22655 ? bht_bank_rd_data_out_1_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23329 = _T_23328 | _T_23074; // @[Mux.scala 27:72]
  wire  _T_22657 = bht_rd_addr_hashed_f == 8'h5e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_94; // @[Reg.scala 27:20]
  wire [1:0] _T_23075 = _T_22657 ? bht_bank_rd_data_out_1_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23330 = _T_23329 | _T_23075; // @[Mux.scala 27:72]
  wire  _T_22659 = bht_rd_addr_hashed_f == 8'h5f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_95; // @[Reg.scala 27:20]
  wire [1:0] _T_23076 = _T_22659 ? bht_bank_rd_data_out_1_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23331 = _T_23330 | _T_23076; // @[Mux.scala 27:72]
  wire  _T_22661 = bht_rd_addr_hashed_f == 8'h60; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_96; // @[Reg.scala 27:20]
  wire [1:0] _T_23077 = _T_22661 ? bht_bank_rd_data_out_1_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23332 = _T_23331 | _T_23077; // @[Mux.scala 27:72]
  wire  _T_22663 = bht_rd_addr_hashed_f == 8'h61; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_97; // @[Reg.scala 27:20]
  wire [1:0] _T_23078 = _T_22663 ? bht_bank_rd_data_out_1_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23333 = _T_23332 | _T_23078; // @[Mux.scala 27:72]
  wire  _T_22665 = bht_rd_addr_hashed_f == 8'h62; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_98; // @[Reg.scala 27:20]
  wire [1:0] _T_23079 = _T_22665 ? bht_bank_rd_data_out_1_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23334 = _T_23333 | _T_23079; // @[Mux.scala 27:72]
  wire  _T_22667 = bht_rd_addr_hashed_f == 8'h63; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_99; // @[Reg.scala 27:20]
  wire [1:0] _T_23080 = _T_22667 ? bht_bank_rd_data_out_1_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23335 = _T_23334 | _T_23080; // @[Mux.scala 27:72]
  wire  _T_22669 = bht_rd_addr_hashed_f == 8'h64; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_100; // @[Reg.scala 27:20]
  wire [1:0] _T_23081 = _T_22669 ? bht_bank_rd_data_out_1_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23336 = _T_23335 | _T_23081; // @[Mux.scala 27:72]
  wire  _T_22671 = bht_rd_addr_hashed_f == 8'h65; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_101; // @[Reg.scala 27:20]
  wire [1:0] _T_23082 = _T_22671 ? bht_bank_rd_data_out_1_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23337 = _T_23336 | _T_23082; // @[Mux.scala 27:72]
  wire  _T_22673 = bht_rd_addr_hashed_f == 8'h66; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_102; // @[Reg.scala 27:20]
  wire [1:0] _T_23083 = _T_22673 ? bht_bank_rd_data_out_1_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23338 = _T_23337 | _T_23083; // @[Mux.scala 27:72]
  wire  _T_22675 = bht_rd_addr_hashed_f == 8'h67; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_103; // @[Reg.scala 27:20]
  wire [1:0] _T_23084 = _T_22675 ? bht_bank_rd_data_out_1_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23339 = _T_23338 | _T_23084; // @[Mux.scala 27:72]
  wire  _T_22677 = bht_rd_addr_hashed_f == 8'h68; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_104; // @[Reg.scala 27:20]
  wire [1:0] _T_23085 = _T_22677 ? bht_bank_rd_data_out_1_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23340 = _T_23339 | _T_23085; // @[Mux.scala 27:72]
  wire  _T_22679 = bht_rd_addr_hashed_f == 8'h69; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_105; // @[Reg.scala 27:20]
  wire [1:0] _T_23086 = _T_22679 ? bht_bank_rd_data_out_1_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23341 = _T_23340 | _T_23086; // @[Mux.scala 27:72]
  wire  _T_22681 = bht_rd_addr_hashed_f == 8'h6a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_106; // @[Reg.scala 27:20]
  wire [1:0] _T_23087 = _T_22681 ? bht_bank_rd_data_out_1_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23342 = _T_23341 | _T_23087; // @[Mux.scala 27:72]
  wire  _T_22683 = bht_rd_addr_hashed_f == 8'h6b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_107; // @[Reg.scala 27:20]
  wire [1:0] _T_23088 = _T_22683 ? bht_bank_rd_data_out_1_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23343 = _T_23342 | _T_23088; // @[Mux.scala 27:72]
  wire  _T_22685 = bht_rd_addr_hashed_f == 8'h6c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_108; // @[Reg.scala 27:20]
  wire [1:0] _T_23089 = _T_22685 ? bht_bank_rd_data_out_1_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23344 = _T_23343 | _T_23089; // @[Mux.scala 27:72]
  wire  _T_22687 = bht_rd_addr_hashed_f == 8'h6d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_109; // @[Reg.scala 27:20]
  wire [1:0] _T_23090 = _T_22687 ? bht_bank_rd_data_out_1_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23345 = _T_23344 | _T_23090; // @[Mux.scala 27:72]
  wire  _T_22689 = bht_rd_addr_hashed_f == 8'h6e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_110; // @[Reg.scala 27:20]
  wire [1:0] _T_23091 = _T_22689 ? bht_bank_rd_data_out_1_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23346 = _T_23345 | _T_23091; // @[Mux.scala 27:72]
  wire  _T_22691 = bht_rd_addr_hashed_f == 8'h6f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_111; // @[Reg.scala 27:20]
  wire [1:0] _T_23092 = _T_22691 ? bht_bank_rd_data_out_1_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23347 = _T_23346 | _T_23092; // @[Mux.scala 27:72]
  wire  _T_22693 = bht_rd_addr_hashed_f == 8'h70; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_112; // @[Reg.scala 27:20]
  wire [1:0] _T_23093 = _T_22693 ? bht_bank_rd_data_out_1_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23348 = _T_23347 | _T_23093; // @[Mux.scala 27:72]
  wire  _T_22695 = bht_rd_addr_hashed_f == 8'h71; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_113; // @[Reg.scala 27:20]
  wire [1:0] _T_23094 = _T_22695 ? bht_bank_rd_data_out_1_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23349 = _T_23348 | _T_23094; // @[Mux.scala 27:72]
  wire  _T_22697 = bht_rd_addr_hashed_f == 8'h72; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_114; // @[Reg.scala 27:20]
  wire [1:0] _T_23095 = _T_22697 ? bht_bank_rd_data_out_1_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23350 = _T_23349 | _T_23095; // @[Mux.scala 27:72]
  wire  _T_22699 = bht_rd_addr_hashed_f == 8'h73; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_115; // @[Reg.scala 27:20]
  wire [1:0] _T_23096 = _T_22699 ? bht_bank_rd_data_out_1_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23351 = _T_23350 | _T_23096; // @[Mux.scala 27:72]
  wire  _T_22701 = bht_rd_addr_hashed_f == 8'h74; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_116; // @[Reg.scala 27:20]
  wire [1:0] _T_23097 = _T_22701 ? bht_bank_rd_data_out_1_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23352 = _T_23351 | _T_23097; // @[Mux.scala 27:72]
  wire  _T_22703 = bht_rd_addr_hashed_f == 8'h75; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_117; // @[Reg.scala 27:20]
  wire [1:0] _T_23098 = _T_22703 ? bht_bank_rd_data_out_1_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23353 = _T_23352 | _T_23098; // @[Mux.scala 27:72]
  wire  _T_22705 = bht_rd_addr_hashed_f == 8'h76; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_118; // @[Reg.scala 27:20]
  wire [1:0] _T_23099 = _T_22705 ? bht_bank_rd_data_out_1_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23354 = _T_23353 | _T_23099; // @[Mux.scala 27:72]
  wire  _T_22707 = bht_rd_addr_hashed_f == 8'h77; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_119; // @[Reg.scala 27:20]
  wire [1:0] _T_23100 = _T_22707 ? bht_bank_rd_data_out_1_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23355 = _T_23354 | _T_23100; // @[Mux.scala 27:72]
  wire  _T_22709 = bht_rd_addr_hashed_f == 8'h78; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_120; // @[Reg.scala 27:20]
  wire [1:0] _T_23101 = _T_22709 ? bht_bank_rd_data_out_1_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23356 = _T_23355 | _T_23101; // @[Mux.scala 27:72]
  wire  _T_22711 = bht_rd_addr_hashed_f == 8'h79; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_121; // @[Reg.scala 27:20]
  wire [1:0] _T_23102 = _T_22711 ? bht_bank_rd_data_out_1_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23357 = _T_23356 | _T_23102; // @[Mux.scala 27:72]
  wire  _T_22713 = bht_rd_addr_hashed_f == 8'h7a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_122; // @[Reg.scala 27:20]
  wire [1:0] _T_23103 = _T_22713 ? bht_bank_rd_data_out_1_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23358 = _T_23357 | _T_23103; // @[Mux.scala 27:72]
  wire  _T_22715 = bht_rd_addr_hashed_f == 8'h7b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_123; // @[Reg.scala 27:20]
  wire [1:0] _T_23104 = _T_22715 ? bht_bank_rd_data_out_1_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23359 = _T_23358 | _T_23104; // @[Mux.scala 27:72]
  wire  _T_22717 = bht_rd_addr_hashed_f == 8'h7c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_124; // @[Reg.scala 27:20]
  wire [1:0] _T_23105 = _T_22717 ? bht_bank_rd_data_out_1_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23360 = _T_23359 | _T_23105; // @[Mux.scala 27:72]
  wire  _T_22719 = bht_rd_addr_hashed_f == 8'h7d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_125; // @[Reg.scala 27:20]
  wire [1:0] _T_23106 = _T_22719 ? bht_bank_rd_data_out_1_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23361 = _T_23360 | _T_23106; // @[Mux.scala 27:72]
  wire  _T_22721 = bht_rd_addr_hashed_f == 8'h7e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_126; // @[Reg.scala 27:20]
  wire [1:0] _T_23107 = _T_22721 ? bht_bank_rd_data_out_1_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23362 = _T_23361 | _T_23107; // @[Mux.scala 27:72]
  wire  _T_22723 = bht_rd_addr_hashed_f == 8'h7f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_127; // @[Reg.scala 27:20]
  wire [1:0] _T_23108 = _T_22723 ? bht_bank_rd_data_out_1_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23363 = _T_23362 | _T_23108; // @[Mux.scala 27:72]
  wire  _T_22725 = bht_rd_addr_hashed_f == 8'h80; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_128; // @[Reg.scala 27:20]
  wire [1:0] _T_23109 = _T_22725 ? bht_bank_rd_data_out_1_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23364 = _T_23363 | _T_23109; // @[Mux.scala 27:72]
  wire  _T_22727 = bht_rd_addr_hashed_f == 8'h81; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_129; // @[Reg.scala 27:20]
  wire [1:0] _T_23110 = _T_22727 ? bht_bank_rd_data_out_1_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23365 = _T_23364 | _T_23110; // @[Mux.scala 27:72]
  wire  _T_22729 = bht_rd_addr_hashed_f == 8'h82; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_130; // @[Reg.scala 27:20]
  wire [1:0] _T_23111 = _T_22729 ? bht_bank_rd_data_out_1_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23366 = _T_23365 | _T_23111; // @[Mux.scala 27:72]
  wire  _T_22731 = bht_rd_addr_hashed_f == 8'h83; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_131; // @[Reg.scala 27:20]
  wire [1:0] _T_23112 = _T_22731 ? bht_bank_rd_data_out_1_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23367 = _T_23366 | _T_23112; // @[Mux.scala 27:72]
  wire  _T_22733 = bht_rd_addr_hashed_f == 8'h84; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_132; // @[Reg.scala 27:20]
  wire [1:0] _T_23113 = _T_22733 ? bht_bank_rd_data_out_1_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23368 = _T_23367 | _T_23113; // @[Mux.scala 27:72]
  wire  _T_22735 = bht_rd_addr_hashed_f == 8'h85; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_133; // @[Reg.scala 27:20]
  wire [1:0] _T_23114 = _T_22735 ? bht_bank_rd_data_out_1_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23369 = _T_23368 | _T_23114; // @[Mux.scala 27:72]
  wire  _T_22737 = bht_rd_addr_hashed_f == 8'h86; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_134; // @[Reg.scala 27:20]
  wire [1:0] _T_23115 = _T_22737 ? bht_bank_rd_data_out_1_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23370 = _T_23369 | _T_23115; // @[Mux.scala 27:72]
  wire  _T_22739 = bht_rd_addr_hashed_f == 8'h87; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_135; // @[Reg.scala 27:20]
  wire [1:0] _T_23116 = _T_22739 ? bht_bank_rd_data_out_1_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23371 = _T_23370 | _T_23116; // @[Mux.scala 27:72]
  wire  _T_22741 = bht_rd_addr_hashed_f == 8'h88; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_136; // @[Reg.scala 27:20]
  wire [1:0] _T_23117 = _T_22741 ? bht_bank_rd_data_out_1_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23372 = _T_23371 | _T_23117; // @[Mux.scala 27:72]
  wire  _T_22743 = bht_rd_addr_hashed_f == 8'h89; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_137; // @[Reg.scala 27:20]
  wire [1:0] _T_23118 = _T_22743 ? bht_bank_rd_data_out_1_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23373 = _T_23372 | _T_23118; // @[Mux.scala 27:72]
  wire  _T_22745 = bht_rd_addr_hashed_f == 8'h8a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_138; // @[Reg.scala 27:20]
  wire [1:0] _T_23119 = _T_22745 ? bht_bank_rd_data_out_1_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23374 = _T_23373 | _T_23119; // @[Mux.scala 27:72]
  wire  _T_22747 = bht_rd_addr_hashed_f == 8'h8b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_139; // @[Reg.scala 27:20]
  wire [1:0] _T_23120 = _T_22747 ? bht_bank_rd_data_out_1_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23375 = _T_23374 | _T_23120; // @[Mux.scala 27:72]
  wire  _T_22749 = bht_rd_addr_hashed_f == 8'h8c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_140; // @[Reg.scala 27:20]
  wire [1:0] _T_23121 = _T_22749 ? bht_bank_rd_data_out_1_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23376 = _T_23375 | _T_23121; // @[Mux.scala 27:72]
  wire  _T_22751 = bht_rd_addr_hashed_f == 8'h8d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_141; // @[Reg.scala 27:20]
  wire [1:0] _T_23122 = _T_22751 ? bht_bank_rd_data_out_1_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23377 = _T_23376 | _T_23122; // @[Mux.scala 27:72]
  wire  _T_22753 = bht_rd_addr_hashed_f == 8'h8e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_142; // @[Reg.scala 27:20]
  wire [1:0] _T_23123 = _T_22753 ? bht_bank_rd_data_out_1_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23378 = _T_23377 | _T_23123; // @[Mux.scala 27:72]
  wire  _T_22755 = bht_rd_addr_hashed_f == 8'h8f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_143; // @[Reg.scala 27:20]
  wire [1:0] _T_23124 = _T_22755 ? bht_bank_rd_data_out_1_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23379 = _T_23378 | _T_23124; // @[Mux.scala 27:72]
  wire  _T_22757 = bht_rd_addr_hashed_f == 8'h90; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_144; // @[Reg.scala 27:20]
  wire [1:0] _T_23125 = _T_22757 ? bht_bank_rd_data_out_1_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23380 = _T_23379 | _T_23125; // @[Mux.scala 27:72]
  wire  _T_22759 = bht_rd_addr_hashed_f == 8'h91; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_145; // @[Reg.scala 27:20]
  wire [1:0] _T_23126 = _T_22759 ? bht_bank_rd_data_out_1_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23381 = _T_23380 | _T_23126; // @[Mux.scala 27:72]
  wire  _T_22761 = bht_rd_addr_hashed_f == 8'h92; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_146; // @[Reg.scala 27:20]
  wire [1:0] _T_23127 = _T_22761 ? bht_bank_rd_data_out_1_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23382 = _T_23381 | _T_23127; // @[Mux.scala 27:72]
  wire  _T_22763 = bht_rd_addr_hashed_f == 8'h93; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_147; // @[Reg.scala 27:20]
  wire [1:0] _T_23128 = _T_22763 ? bht_bank_rd_data_out_1_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23383 = _T_23382 | _T_23128; // @[Mux.scala 27:72]
  wire  _T_22765 = bht_rd_addr_hashed_f == 8'h94; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_148; // @[Reg.scala 27:20]
  wire [1:0] _T_23129 = _T_22765 ? bht_bank_rd_data_out_1_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23384 = _T_23383 | _T_23129; // @[Mux.scala 27:72]
  wire  _T_22767 = bht_rd_addr_hashed_f == 8'h95; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_149; // @[Reg.scala 27:20]
  wire [1:0] _T_23130 = _T_22767 ? bht_bank_rd_data_out_1_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23385 = _T_23384 | _T_23130; // @[Mux.scala 27:72]
  wire  _T_22769 = bht_rd_addr_hashed_f == 8'h96; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_150; // @[Reg.scala 27:20]
  wire [1:0] _T_23131 = _T_22769 ? bht_bank_rd_data_out_1_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23386 = _T_23385 | _T_23131; // @[Mux.scala 27:72]
  wire  _T_22771 = bht_rd_addr_hashed_f == 8'h97; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_151; // @[Reg.scala 27:20]
  wire [1:0] _T_23132 = _T_22771 ? bht_bank_rd_data_out_1_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23387 = _T_23386 | _T_23132; // @[Mux.scala 27:72]
  wire  _T_22773 = bht_rd_addr_hashed_f == 8'h98; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_152; // @[Reg.scala 27:20]
  wire [1:0] _T_23133 = _T_22773 ? bht_bank_rd_data_out_1_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23388 = _T_23387 | _T_23133; // @[Mux.scala 27:72]
  wire  _T_22775 = bht_rd_addr_hashed_f == 8'h99; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_153; // @[Reg.scala 27:20]
  wire [1:0] _T_23134 = _T_22775 ? bht_bank_rd_data_out_1_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23389 = _T_23388 | _T_23134; // @[Mux.scala 27:72]
  wire  _T_22777 = bht_rd_addr_hashed_f == 8'h9a; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_154; // @[Reg.scala 27:20]
  wire [1:0] _T_23135 = _T_22777 ? bht_bank_rd_data_out_1_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23390 = _T_23389 | _T_23135; // @[Mux.scala 27:72]
  wire  _T_22779 = bht_rd_addr_hashed_f == 8'h9b; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_155; // @[Reg.scala 27:20]
  wire [1:0] _T_23136 = _T_22779 ? bht_bank_rd_data_out_1_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23391 = _T_23390 | _T_23136; // @[Mux.scala 27:72]
  wire  _T_22781 = bht_rd_addr_hashed_f == 8'h9c; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_156; // @[Reg.scala 27:20]
  wire [1:0] _T_23137 = _T_22781 ? bht_bank_rd_data_out_1_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23392 = _T_23391 | _T_23137; // @[Mux.scala 27:72]
  wire  _T_22783 = bht_rd_addr_hashed_f == 8'h9d; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_157; // @[Reg.scala 27:20]
  wire [1:0] _T_23138 = _T_22783 ? bht_bank_rd_data_out_1_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23393 = _T_23392 | _T_23138; // @[Mux.scala 27:72]
  wire  _T_22785 = bht_rd_addr_hashed_f == 8'h9e; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_158; // @[Reg.scala 27:20]
  wire [1:0] _T_23139 = _T_22785 ? bht_bank_rd_data_out_1_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23394 = _T_23393 | _T_23139; // @[Mux.scala 27:72]
  wire  _T_22787 = bht_rd_addr_hashed_f == 8'h9f; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_159; // @[Reg.scala 27:20]
  wire [1:0] _T_23140 = _T_22787 ? bht_bank_rd_data_out_1_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23395 = _T_23394 | _T_23140; // @[Mux.scala 27:72]
  wire  _T_22789 = bht_rd_addr_hashed_f == 8'ha0; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_160; // @[Reg.scala 27:20]
  wire [1:0] _T_23141 = _T_22789 ? bht_bank_rd_data_out_1_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23396 = _T_23395 | _T_23141; // @[Mux.scala 27:72]
  wire  _T_22791 = bht_rd_addr_hashed_f == 8'ha1; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_161; // @[Reg.scala 27:20]
  wire [1:0] _T_23142 = _T_22791 ? bht_bank_rd_data_out_1_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23397 = _T_23396 | _T_23142; // @[Mux.scala 27:72]
  wire  _T_22793 = bht_rd_addr_hashed_f == 8'ha2; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_162; // @[Reg.scala 27:20]
  wire [1:0] _T_23143 = _T_22793 ? bht_bank_rd_data_out_1_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23398 = _T_23397 | _T_23143; // @[Mux.scala 27:72]
  wire  _T_22795 = bht_rd_addr_hashed_f == 8'ha3; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_163; // @[Reg.scala 27:20]
  wire [1:0] _T_23144 = _T_22795 ? bht_bank_rd_data_out_1_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23399 = _T_23398 | _T_23144; // @[Mux.scala 27:72]
  wire  _T_22797 = bht_rd_addr_hashed_f == 8'ha4; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_164; // @[Reg.scala 27:20]
  wire [1:0] _T_23145 = _T_22797 ? bht_bank_rd_data_out_1_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23400 = _T_23399 | _T_23145; // @[Mux.scala 27:72]
  wire  _T_22799 = bht_rd_addr_hashed_f == 8'ha5; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_165; // @[Reg.scala 27:20]
  wire [1:0] _T_23146 = _T_22799 ? bht_bank_rd_data_out_1_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23401 = _T_23400 | _T_23146; // @[Mux.scala 27:72]
  wire  _T_22801 = bht_rd_addr_hashed_f == 8'ha6; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_166; // @[Reg.scala 27:20]
  wire [1:0] _T_23147 = _T_22801 ? bht_bank_rd_data_out_1_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23402 = _T_23401 | _T_23147; // @[Mux.scala 27:72]
  wire  _T_22803 = bht_rd_addr_hashed_f == 8'ha7; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_167; // @[Reg.scala 27:20]
  wire [1:0] _T_23148 = _T_22803 ? bht_bank_rd_data_out_1_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23403 = _T_23402 | _T_23148; // @[Mux.scala 27:72]
  wire  _T_22805 = bht_rd_addr_hashed_f == 8'ha8; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_168; // @[Reg.scala 27:20]
  wire [1:0] _T_23149 = _T_22805 ? bht_bank_rd_data_out_1_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23404 = _T_23403 | _T_23149; // @[Mux.scala 27:72]
  wire  _T_22807 = bht_rd_addr_hashed_f == 8'ha9; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_169; // @[Reg.scala 27:20]
  wire [1:0] _T_23150 = _T_22807 ? bht_bank_rd_data_out_1_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23405 = _T_23404 | _T_23150; // @[Mux.scala 27:72]
  wire  _T_22809 = bht_rd_addr_hashed_f == 8'haa; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_170; // @[Reg.scala 27:20]
  wire [1:0] _T_23151 = _T_22809 ? bht_bank_rd_data_out_1_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23406 = _T_23405 | _T_23151; // @[Mux.scala 27:72]
  wire  _T_22811 = bht_rd_addr_hashed_f == 8'hab; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_171; // @[Reg.scala 27:20]
  wire [1:0] _T_23152 = _T_22811 ? bht_bank_rd_data_out_1_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23407 = _T_23406 | _T_23152; // @[Mux.scala 27:72]
  wire  _T_22813 = bht_rd_addr_hashed_f == 8'hac; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_172; // @[Reg.scala 27:20]
  wire [1:0] _T_23153 = _T_22813 ? bht_bank_rd_data_out_1_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23408 = _T_23407 | _T_23153; // @[Mux.scala 27:72]
  wire  _T_22815 = bht_rd_addr_hashed_f == 8'had; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_173; // @[Reg.scala 27:20]
  wire [1:0] _T_23154 = _T_22815 ? bht_bank_rd_data_out_1_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23409 = _T_23408 | _T_23154; // @[Mux.scala 27:72]
  wire  _T_22817 = bht_rd_addr_hashed_f == 8'hae; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_174; // @[Reg.scala 27:20]
  wire [1:0] _T_23155 = _T_22817 ? bht_bank_rd_data_out_1_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23410 = _T_23409 | _T_23155; // @[Mux.scala 27:72]
  wire  _T_22819 = bht_rd_addr_hashed_f == 8'haf; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_175; // @[Reg.scala 27:20]
  wire [1:0] _T_23156 = _T_22819 ? bht_bank_rd_data_out_1_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23411 = _T_23410 | _T_23156; // @[Mux.scala 27:72]
  wire  _T_22821 = bht_rd_addr_hashed_f == 8'hb0; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_176; // @[Reg.scala 27:20]
  wire [1:0] _T_23157 = _T_22821 ? bht_bank_rd_data_out_1_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23412 = _T_23411 | _T_23157; // @[Mux.scala 27:72]
  wire  _T_22823 = bht_rd_addr_hashed_f == 8'hb1; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_177; // @[Reg.scala 27:20]
  wire [1:0] _T_23158 = _T_22823 ? bht_bank_rd_data_out_1_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23413 = _T_23412 | _T_23158; // @[Mux.scala 27:72]
  wire  _T_22825 = bht_rd_addr_hashed_f == 8'hb2; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_178; // @[Reg.scala 27:20]
  wire [1:0] _T_23159 = _T_22825 ? bht_bank_rd_data_out_1_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23414 = _T_23413 | _T_23159; // @[Mux.scala 27:72]
  wire  _T_22827 = bht_rd_addr_hashed_f == 8'hb3; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_179; // @[Reg.scala 27:20]
  wire [1:0] _T_23160 = _T_22827 ? bht_bank_rd_data_out_1_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23415 = _T_23414 | _T_23160; // @[Mux.scala 27:72]
  wire  _T_22829 = bht_rd_addr_hashed_f == 8'hb4; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_180; // @[Reg.scala 27:20]
  wire [1:0] _T_23161 = _T_22829 ? bht_bank_rd_data_out_1_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23416 = _T_23415 | _T_23161; // @[Mux.scala 27:72]
  wire  _T_22831 = bht_rd_addr_hashed_f == 8'hb5; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_181; // @[Reg.scala 27:20]
  wire [1:0] _T_23162 = _T_22831 ? bht_bank_rd_data_out_1_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23417 = _T_23416 | _T_23162; // @[Mux.scala 27:72]
  wire  _T_22833 = bht_rd_addr_hashed_f == 8'hb6; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_182; // @[Reg.scala 27:20]
  wire [1:0] _T_23163 = _T_22833 ? bht_bank_rd_data_out_1_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23418 = _T_23417 | _T_23163; // @[Mux.scala 27:72]
  wire  _T_22835 = bht_rd_addr_hashed_f == 8'hb7; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_183; // @[Reg.scala 27:20]
  wire [1:0] _T_23164 = _T_22835 ? bht_bank_rd_data_out_1_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23419 = _T_23418 | _T_23164; // @[Mux.scala 27:72]
  wire  _T_22837 = bht_rd_addr_hashed_f == 8'hb8; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_184; // @[Reg.scala 27:20]
  wire [1:0] _T_23165 = _T_22837 ? bht_bank_rd_data_out_1_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23420 = _T_23419 | _T_23165; // @[Mux.scala 27:72]
  wire  _T_22839 = bht_rd_addr_hashed_f == 8'hb9; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_185; // @[Reg.scala 27:20]
  wire [1:0] _T_23166 = _T_22839 ? bht_bank_rd_data_out_1_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23421 = _T_23420 | _T_23166; // @[Mux.scala 27:72]
  wire  _T_22841 = bht_rd_addr_hashed_f == 8'hba; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_186; // @[Reg.scala 27:20]
  wire [1:0] _T_23167 = _T_22841 ? bht_bank_rd_data_out_1_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23422 = _T_23421 | _T_23167; // @[Mux.scala 27:72]
  wire  _T_22843 = bht_rd_addr_hashed_f == 8'hbb; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_187; // @[Reg.scala 27:20]
  wire [1:0] _T_23168 = _T_22843 ? bht_bank_rd_data_out_1_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23423 = _T_23422 | _T_23168; // @[Mux.scala 27:72]
  wire  _T_22845 = bht_rd_addr_hashed_f == 8'hbc; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_188; // @[Reg.scala 27:20]
  wire [1:0] _T_23169 = _T_22845 ? bht_bank_rd_data_out_1_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23424 = _T_23423 | _T_23169; // @[Mux.scala 27:72]
  wire  _T_22847 = bht_rd_addr_hashed_f == 8'hbd; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_189; // @[Reg.scala 27:20]
  wire [1:0] _T_23170 = _T_22847 ? bht_bank_rd_data_out_1_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23425 = _T_23424 | _T_23170; // @[Mux.scala 27:72]
  wire  _T_22849 = bht_rd_addr_hashed_f == 8'hbe; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_190; // @[Reg.scala 27:20]
  wire [1:0] _T_23171 = _T_22849 ? bht_bank_rd_data_out_1_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23426 = _T_23425 | _T_23171; // @[Mux.scala 27:72]
  wire  _T_22851 = bht_rd_addr_hashed_f == 8'hbf; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_191; // @[Reg.scala 27:20]
  wire [1:0] _T_23172 = _T_22851 ? bht_bank_rd_data_out_1_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23427 = _T_23426 | _T_23172; // @[Mux.scala 27:72]
  wire  _T_22853 = bht_rd_addr_hashed_f == 8'hc0; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_192; // @[Reg.scala 27:20]
  wire [1:0] _T_23173 = _T_22853 ? bht_bank_rd_data_out_1_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23428 = _T_23427 | _T_23173; // @[Mux.scala 27:72]
  wire  _T_22855 = bht_rd_addr_hashed_f == 8'hc1; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_193; // @[Reg.scala 27:20]
  wire [1:0] _T_23174 = _T_22855 ? bht_bank_rd_data_out_1_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23429 = _T_23428 | _T_23174; // @[Mux.scala 27:72]
  wire  _T_22857 = bht_rd_addr_hashed_f == 8'hc2; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_194; // @[Reg.scala 27:20]
  wire [1:0] _T_23175 = _T_22857 ? bht_bank_rd_data_out_1_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23430 = _T_23429 | _T_23175; // @[Mux.scala 27:72]
  wire  _T_22859 = bht_rd_addr_hashed_f == 8'hc3; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_195; // @[Reg.scala 27:20]
  wire [1:0] _T_23176 = _T_22859 ? bht_bank_rd_data_out_1_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23431 = _T_23430 | _T_23176; // @[Mux.scala 27:72]
  wire  _T_22861 = bht_rd_addr_hashed_f == 8'hc4; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_196; // @[Reg.scala 27:20]
  wire [1:0] _T_23177 = _T_22861 ? bht_bank_rd_data_out_1_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23432 = _T_23431 | _T_23177; // @[Mux.scala 27:72]
  wire  _T_22863 = bht_rd_addr_hashed_f == 8'hc5; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_197; // @[Reg.scala 27:20]
  wire [1:0] _T_23178 = _T_22863 ? bht_bank_rd_data_out_1_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23433 = _T_23432 | _T_23178; // @[Mux.scala 27:72]
  wire  _T_22865 = bht_rd_addr_hashed_f == 8'hc6; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_198; // @[Reg.scala 27:20]
  wire [1:0] _T_23179 = _T_22865 ? bht_bank_rd_data_out_1_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23434 = _T_23433 | _T_23179; // @[Mux.scala 27:72]
  wire  _T_22867 = bht_rd_addr_hashed_f == 8'hc7; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_199; // @[Reg.scala 27:20]
  wire [1:0] _T_23180 = _T_22867 ? bht_bank_rd_data_out_1_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23435 = _T_23434 | _T_23180; // @[Mux.scala 27:72]
  wire  _T_22869 = bht_rd_addr_hashed_f == 8'hc8; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_200; // @[Reg.scala 27:20]
  wire [1:0] _T_23181 = _T_22869 ? bht_bank_rd_data_out_1_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23436 = _T_23435 | _T_23181; // @[Mux.scala 27:72]
  wire  _T_22871 = bht_rd_addr_hashed_f == 8'hc9; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_201; // @[Reg.scala 27:20]
  wire [1:0] _T_23182 = _T_22871 ? bht_bank_rd_data_out_1_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23437 = _T_23436 | _T_23182; // @[Mux.scala 27:72]
  wire  _T_22873 = bht_rd_addr_hashed_f == 8'hca; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_202; // @[Reg.scala 27:20]
  wire [1:0] _T_23183 = _T_22873 ? bht_bank_rd_data_out_1_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23438 = _T_23437 | _T_23183; // @[Mux.scala 27:72]
  wire  _T_22875 = bht_rd_addr_hashed_f == 8'hcb; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_203; // @[Reg.scala 27:20]
  wire [1:0] _T_23184 = _T_22875 ? bht_bank_rd_data_out_1_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23439 = _T_23438 | _T_23184; // @[Mux.scala 27:72]
  wire  _T_22877 = bht_rd_addr_hashed_f == 8'hcc; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_204; // @[Reg.scala 27:20]
  wire [1:0] _T_23185 = _T_22877 ? bht_bank_rd_data_out_1_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23440 = _T_23439 | _T_23185; // @[Mux.scala 27:72]
  wire  _T_22879 = bht_rd_addr_hashed_f == 8'hcd; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_205; // @[Reg.scala 27:20]
  wire [1:0] _T_23186 = _T_22879 ? bht_bank_rd_data_out_1_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23441 = _T_23440 | _T_23186; // @[Mux.scala 27:72]
  wire  _T_22881 = bht_rd_addr_hashed_f == 8'hce; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_206; // @[Reg.scala 27:20]
  wire [1:0] _T_23187 = _T_22881 ? bht_bank_rd_data_out_1_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23442 = _T_23441 | _T_23187; // @[Mux.scala 27:72]
  wire  _T_22883 = bht_rd_addr_hashed_f == 8'hcf; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_207; // @[Reg.scala 27:20]
  wire [1:0] _T_23188 = _T_22883 ? bht_bank_rd_data_out_1_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23443 = _T_23442 | _T_23188; // @[Mux.scala 27:72]
  wire  _T_22885 = bht_rd_addr_hashed_f == 8'hd0; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_208; // @[Reg.scala 27:20]
  wire [1:0] _T_23189 = _T_22885 ? bht_bank_rd_data_out_1_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23444 = _T_23443 | _T_23189; // @[Mux.scala 27:72]
  wire  _T_22887 = bht_rd_addr_hashed_f == 8'hd1; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_209; // @[Reg.scala 27:20]
  wire [1:0] _T_23190 = _T_22887 ? bht_bank_rd_data_out_1_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23445 = _T_23444 | _T_23190; // @[Mux.scala 27:72]
  wire  _T_22889 = bht_rd_addr_hashed_f == 8'hd2; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_210; // @[Reg.scala 27:20]
  wire [1:0] _T_23191 = _T_22889 ? bht_bank_rd_data_out_1_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23446 = _T_23445 | _T_23191; // @[Mux.scala 27:72]
  wire  _T_22891 = bht_rd_addr_hashed_f == 8'hd3; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_211; // @[Reg.scala 27:20]
  wire [1:0] _T_23192 = _T_22891 ? bht_bank_rd_data_out_1_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23447 = _T_23446 | _T_23192; // @[Mux.scala 27:72]
  wire  _T_22893 = bht_rd_addr_hashed_f == 8'hd4; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_212; // @[Reg.scala 27:20]
  wire [1:0] _T_23193 = _T_22893 ? bht_bank_rd_data_out_1_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23448 = _T_23447 | _T_23193; // @[Mux.scala 27:72]
  wire  _T_22895 = bht_rd_addr_hashed_f == 8'hd5; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_213; // @[Reg.scala 27:20]
  wire [1:0] _T_23194 = _T_22895 ? bht_bank_rd_data_out_1_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23449 = _T_23448 | _T_23194; // @[Mux.scala 27:72]
  wire  _T_22897 = bht_rd_addr_hashed_f == 8'hd6; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_214; // @[Reg.scala 27:20]
  wire [1:0] _T_23195 = _T_22897 ? bht_bank_rd_data_out_1_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23450 = _T_23449 | _T_23195; // @[Mux.scala 27:72]
  wire  _T_22899 = bht_rd_addr_hashed_f == 8'hd7; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_215; // @[Reg.scala 27:20]
  wire [1:0] _T_23196 = _T_22899 ? bht_bank_rd_data_out_1_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23451 = _T_23450 | _T_23196; // @[Mux.scala 27:72]
  wire  _T_22901 = bht_rd_addr_hashed_f == 8'hd8; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_216; // @[Reg.scala 27:20]
  wire [1:0] _T_23197 = _T_22901 ? bht_bank_rd_data_out_1_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23452 = _T_23451 | _T_23197; // @[Mux.scala 27:72]
  wire  _T_22903 = bht_rd_addr_hashed_f == 8'hd9; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_217; // @[Reg.scala 27:20]
  wire [1:0] _T_23198 = _T_22903 ? bht_bank_rd_data_out_1_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23453 = _T_23452 | _T_23198; // @[Mux.scala 27:72]
  wire  _T_22905 = bht_rd_addr_hashed_f == 8'hda; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_218; // @[Reg.scala 27:20]
  wire [1:0] _T_23199 = _T_22905 ? bht_bank_rd_data_out_1_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23454 = _T_23453 | _T_23199; // @[Mux.scala 27:72]
  wire  _T_22907 = bht_rd_addr_hashed_f == 8'hdb; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_219; // @[Reg.scala 27:20]
  wire [1:0] _T_23200 = _T_22907 ? bht_bank_rd_data_out_1_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23455 = _T_23454 | _T_23200; // @[Mux.scala 27:72]
  wire  _T_22909 = bht_rd_addr_hashed_f == 8'hdc; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_220; // @[Reg.scala 27:20]
  wire [1:0] _T_23201 = _T_22909 ? bht_bank_rd_data_out_1_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23456 = _T_23455 | _T_23201; // @[Mux.scala 27:72]
  wire  _T_22911 = bht_rd_addr_hashed_f == 8'hdd; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_221; // @[Reg.scala 27:20]
  wire [1:0] _T_23202 = _T_22911 ? bht_bank_rd_data_out_1_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23457 = _T_23456 | _T_23202; // @[Mux.scala 27:72]
  wire  _T_22913 = bht_rd_addr_hashed_f == 8'hde; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_222; // @[Reg.scala 27:20]
  wire [1:0] _T_23203 = _T_22913 ? bht_bank_rd_data_out_1_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23458 = _T_23457 | _T_23203; // @[Mux.scala 27:72]
  wire  _T_22915 = bht_rd_addr_hashed_f == 8'hdf; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_223; // @[Reg.scala 27:20]
  wire [1:0] _T_23204 = _T_22915 ? bht_bank_rd_data_out_1_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23459 = _T_23458 | _T_23204; // @[Mux.scala 27:72]
  wire  _T_22917 = bht_rd_addr_hashed_f == 8'he0; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_224; // @[Reg.scala 27:20]
  wire [1:0] _T_23205 = _T_22917 ? bht_bank_rd_data_out_1_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23460 = _T_23459 | _T_23205; // @[Mux.scala 27:72]
  wire  _T_22919 = bht_rd_addr_hashed_f == 8'he1; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_225; // @[Reg.scala 27:20]
  wire [1:0] _T_23206 = _T_22919 ? bht_bank_rd_data_out_1_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23461 = _T_23460 | _T_23206; // @[Mux.scala 27:72]
  wire  _T_22921 = bht_rd_addr_hashed_f == 8'he2; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_226; // @[Reg.scala 27:20]
  wire [1:0] _T_23207 = _T_22921 ? bht_bank_rd_data_out_1_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23462 = _T_23461 | _T_23207; // @[Mux.scala 27:72]
  wire  _T_22923 = bht_rd_addr_hashed_f == 8'he3; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_227; // @[Reg.scala 27:20]
  wire [1:0] _T_23208 = _T_22923 ? bht_bank_rd_data_out_1_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23463 = _T_23462 | _T_23208; // @[Mux.scala 27:72]
  wire  _T_22925 = bht_rd_addr_hashed_f == 8'he4; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_228; // @[Reg.scala 27:20]
  wire [1:0] _T_23209 = _T_22925 ? bht_bank_rd_data_out_1_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23464 = _T_23463 | _T_23209; // @[Mux.scala 27:72]
  wire  _T_22927 = bht_rd_addr_hashed_f == 8'he5; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_229; // @[Reg.scala 27:20]
  wire [1:0] _T_23210 = _T_22927 ? bht_bank_rd_data_out_1_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23465 = _T_23464 | _T_23210; // @[Mux.scala 27:72]
  wire  _T_22929 = bht_rd_addr_hashed_f == 8'he6; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_230; // @[Reg.scala 27:20]
  wire [1:0] _T_23211 = _T_22929 ? bht_bank_rd_data_out_1_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23466 = _T_23465 | _T_23211; // @[Mux.scala 27:72]
  wire  _T_22931 = bht_rd_addr_hashed_f == 8'he7; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_231; // @[Reg.scala 27:20]
  wire [1:0] _T_23212 = _T_22931 ? bht_bank_rd_data_out_1_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23467 = _T_23466 | _T_23212; // @[Mux.scala 27:72]
  wire  _T_22933 = bht_rd_addr_hashed_f == 8'he8; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_232; // @[Reg.scala 27:20]
  wire [1:0] _T_23213 = _T_22933 ? bht_bank_rd_data_out_1_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23468 = _T_23467 | _T_23213; // @[Mux.scala 27:72]
  wire  _T_22935 = bht_rd_addr_hashed_f == 8'he9; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_233; // @[Reg.scala 27:20]
  wire [1:0] _T_23214 = _T_22935 ? bht_bank_rd_data_out_1_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23469 = _T_23468 | _T_23214; // @[Mux.scala 27:72]
  wire  _T_22937 = bht_rd_addr_hashed_f == 8'hea; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_234; // @[Reg.scala 27:20]
  wire [1:0] _T_23215 = _T_22937 ? bht_bank_rd_data_out_1_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23470 = _T_23469 | _T_23215; // @[Mux.scala 27:72]
  wire  _T_22939 = bht_rd_addr_hashed_f == 8'heb; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_235; // @[Reg.scala 27:20]
  wire [1:0] _T_23216 = _T_22939 ? bht_bank_rd_data_out_1_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23471 = _T_23470 | _T_23216; // @[Mux.scala 27:72]
  wire  _T_22941 = bht_rd_addr_hashed_f == 8'hec; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_236; // @[Reg.scala 27:20]
  wire [1:0] _T_23217 = _T_22941 ? bht_bank_rd_data_out_1_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23472 = _T_23471 | _T_23217; // @[Mux.scala 27:72]
  wire  _T_22943 = bht_rd_addr_hashed_f == 8'hed; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_237; // @[Reg.scala 27:20]
  wire [1:0] _T_23218 = _T_22943 ? bht_bank_rd_data_out_1_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23473 = _T_23472 | _T_23218; // @[Mux.scala 27:72]
  wire  _T_22945 = bht_rd_addr_hashed_f == 8'hee; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_238; // @[Reg.scala 27:20]
  wire [1:0] _T_23219 = _T_22945 ? bht_bank_rd_data_out_1_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23474 = _T_23473 | _T_23219; // @[Mux.scala 27:72]
  wire  _T_22947 = bht_rd_addr_hashed_f == 8'hef; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_239; // @[Reg.scala 27:20]
  wire [1:0] _T_23220 = _T_22947 ? bht_bank_rd_data_out_1_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23475 = _T_23474 | _T_23220; // @[Mux.scala 27:72]
  wire  _T_22949 = bht_rd_addr_hashed_f == 8'hf0; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_240; // @[Reg.scala 27:20]
  wire [1:0] _T_23221 = _T_22949 ? bht_bank_rd_data_out_1_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23476 = _T_23475 | _T_23221; // @[Mux.scala 27:72]
  wire  _T_22951 = bht_rd_addr_hashed_f == 8'hf1; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_241; // @[Reg.scala 27:20]
  wire [1:0] _T_23222 = _T_22951 ? bht_bank_rd_data_out_1_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23477 = _T_23476 | _T_23222; // @[Mux.scala 27:72]
  wire  _T_22953 = bht_rd_addr_hashed_f == 8'hf2; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_242; // @[Reg.scala 27:20]
  wire [1:0] _T_23223 = _T_22953 ? bht_bank_rd_data_out_1_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23478 = _T_23477 | _T_23223; // @[Mux.scala 27:72]
  wire  _T_22955 = bht_rd_addr_hashed_f == 8'hf3; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_243; // @[Reg.scala 27:20]
  wire [1:0] _T_23224 = _T_22955 ? bht_bank_rd_data_out_1_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23479 = _T_23478 | _T_23224; // @[Mux.scala 27:72]
  wire  _T_22957 = bht_rd_addr_hashed_f == 8'hf4; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_244; // @[Reg.scala 27:20]
  wire [1:0] _T_23225 = _T_22957 ? bht_bank_rd_data_out_1_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23480 = _T_23479 | _T_23225; // @[Mux.scala 27:72]
  wire  _T_22959 = bht_rd_addr_hashed_f == 8'hf5; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_245; // @[Reg.scala 27:20]
  wire [1:0] _T_23226 = _T_22959 ? bht_bank_rd_data_out_1_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23481 = _T_23480 | _T_23226; // @[Mux.scala 27:72]
  wire  _T_22961 = bht_rd_addr_hashed_f == 8'hf6; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_246; // @[Reg.scala 27:20]
  wire [1:0] _T_23227 = _T_22961 ? bht_bank_rd_data_out_1_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23482 = _T_23481 | _T_23227; // @[Mux.scala 27:72]
  wire  _T_22963 = bht_rd_addr_hashed_f == 8'hf7; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_247; // @[Reg.scala 27:20]
  wire [1:0] _T_23228 = _T_22963 ? bht_bank_rd_data_out_1_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23483 = _T_23482 | _T_23228; // @[Mux.scala 27:72]
  wire  _T_22965 = bht_rd_addr_hashed_f == 8'hf8; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_248; // @[Reg.scala 27:20]
  wire [1:0] _T_23229 = _T_22965 ? bht_bank_rd_data_out_1_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23484 = _T_23483 | _T_23229; // @[Mux.scala 27:72]
  wire  _T_22967 = bht_rd_addr_hashed_f == 8'hf9; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_249; // @[Reg.scala 27:20]
  wire [1:0] _T_23230 = _T_22967 ? bht_bank_rd_data_out_1_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23485 = _T_23484 | _T_23230; // @[Mux.scala 27:72]
  wire  _T_22969 = bht_rd_addr_hashed_f == 8'hfa; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_250; // @[Reg.scala 27:20]
  wire [1:0] _T_23231 = _T_22969 ? bht_bank_rd_data_out_1_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23486 = _T_23485 | _T_23231; // @[Mux.scala 27:72]
  wire  _T_22971 = bht_rd_addr_hashed_f == 8'hfb; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_251; // @[Reg.scala 27:20]
  wire [1:0] _T_23232 = _T_22971 ? bht_bank_rd_data_out_1_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23487 = _T_23486 | _T_23232; // @[Mux.scala 27:72]
  wire  _T_22973 = bht_rd_addr_hashed_f == 8'hfc; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_252; // @[Reg.scala 27:20]
  wire [1:0] _T_23233 = _T_22973 ? bht_bank_rd_data_out_1_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23488 = _T_23487 | _T_23233; // @[Mux.scala 27:72]
  wire  _T_22975 = bht_rd_addr_hashed_f == 8'hfd; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_253; // @[Reg.scala 27:20]
  wire [1:0] _T_23234 = _T_22975 ? bht_bank_rd_data_out_1_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23489 = _T_23488 | _T_23234; // @[Mux.scala 27:72]
  wire  _T_22977 = bht_rd_addr_hashed_f == 8'hfe; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_254; // @[Reg.scala 27:20]
  wire [1:0] _T_23235 = _T_22977 ? bht_bank_rd_data_out_1_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_23490 = _T_23489 | _T_23235; // @[Mux.scala 27:72]
  wire  _T_22979 = bht_rd_addr_hashed_f == 8'hff; // @[ifu_bp_ctl.scala 531:79]
  reg [1:0] bht_bank_rd_data_out_1_255; // @[Reg.scala 27:20]
  wire [1:0] _T_23236 = _T_22979 ? bht_bank_rd_data_out_1_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank1_rd_data_f = _T_23490 | _T_23236; // @[Mux.scala 27:72]
  wire [1:0] _T_253 = _T_147 ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [9:0] _T_585 = {btb_rd_addr_p1_f,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] bht_rd_addr_hashed_p1_f = _T_585[9:2] ^ fghr; // @[lib.scala 56:35]
  wire  _T_23493 = bht_rd_addr_hashed_p1_f == 8'h0; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_0; // @[Reg.scala 27:20]
  wire [1:0] _T_24005 = _T_23493 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire  _T_23495 = bht_rd_addr_hashed_p1_f == 8'h1; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_1; // @[Reg.scala 27:20]
  wire [1:0] _T_24006 = _T_23495 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24261 = _T_24005 | _T_24006; // @[Mux.scala 27:72]
  wire  _T_23497 = bht_rd_addr_hashed_p1_f == 8'h2; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_2; // @[Reg.scala 27:20]
  wire [1:0] _T_24007 = _T_23497 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24262 = _T_24261 | _T_24007; // @[Mux.scala 27:72]
  wire  _T_23499 = bht_rd_addr_hashed_p1_f == 8'h3; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_3; // @[Reg.scala 27:20]
  wire [1:0] _T_24008 = _T_23499 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24263 = _T_24262 | _T_24008; // @[Mux.scala 27:72]
  wire  _T_23501 = bht_rd_addr_hashed_p1_f == 8'h4; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_4; // @[Reg.scala 27:20]
  wire [1:0] _T_24009 = _T_23501 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24264 = _T_24263 | _T_24009; // @[Mux.scala 27:72]
  wire  _T_23503 = bht_rd_addr_hashed_p1_f == 8'h5; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_5; // @[Reg.scala 27:20]
  wire [1:0] _T_24010 = _T_23503 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24265 = _T_24264 | _T_24010; // @[Mux.scala 27:72]
  wire  _T_23505 = bht_rd_addr_hashed_p1_f == 8'h6; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_6; // @[Reg.scala 27:20]
  wire [1:0] _T_24011 = _T_23505 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24266 = _T_24265 | _T_24011; // @[Mux.scala 27:72]
  wire  _T_23507 = bht_rd_addr_hashed_p1_f == 8'h7; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_7; // @[Reg.scala 27:20]
  wire [1:0] _T_24012 = _T_23507 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24267 = _T_24266 | _T_24012; // @[Mux.scala 27:72]
  wire  _T_23509 = bht_rd_addr_hashed_p1_f == 8'h8; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_8; // @[Reg.scala 27:20]
  wire [1:0] _T_24013 = _T_23509 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24268 = _T_24267 | _T_24013; // @[Mux.scala 27:72]
  wire  _T_23511 = bht_rd_addr_hashed_p1_f == 8'h9; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_9; // @[Reg.scala 27:20]
  wire [1:0] _T_24014 = _T_23511 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24269 = _T_24268 | _T_24014; // @[Mux.scala 27:72]
  wire  _T_23513 = bht_rd_addr_hashed_p1_f == 8'ha; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_10; // @[Reg.scala 27:20]
  wire [1:0] _T_24015 = _T_23513 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24270 = _T_24269 | _T_24015; // @[Mux.scala 27:72]
  wire  _T_23515 = bht_rd_addr_hashed_p1_f == 8'hb; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_11; // @[Reg.scala 27:20]
  wire [1:0] _T_24016 = _T_23515 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24271 = _T_24270 | _T_24016; // @[Mux.scala 27:72]
  wire  _T_23517 = bht_rd_addr_hashed_p1_f == 8'hc; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_12; // @[Reg.scala 27:20]
  wire [1:0] _T_24017 = _T_23517 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24272 = _T_24271 | _T_24017; // @[Mux.scala 27:72]
  wire  _T_23519 = bht_rd_addr_hashed_p1_f == 8'hd; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_13; // @[Reg.scala 27:20]
  wire [1:0] _T_24018 = _T_23519 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24273 = _T_24272 | _T_24018; // @[Mux.scala 27:72]
  wire  _T_23521 = bht_rd_addr_hashed_p1_f == 8'he; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_14; // @[Reg.scala 27:20]
  wire [1:0] _T_24019 = _T_23521 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24274 = _T_24273 | _T_24019; // @[Mux.scala 27:72]
  wire  _T_23523 = bht_rd_addr_hashed_p1_f == 8'hf; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_15; // @[Reg.scala 27:20]
  wire [1:0] _T_24020 = _T_23523 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24275 = _T_24274 | _T_24020; // @[Mux.scala 27:72]
  wire  _T_23525 = bht_rd_addr_hashed_p1_f == 8'h10; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_16; // @[Reg.scala 27:20]
  wire [1:0] _T_24021 = _T_23525 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24276 = _T_24275 | _T_24021; // @[Mux.scala 27:72]
  wire  _T_23527 = bht_rd_addr_hashed_p1_f == 8'h11; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_17; // @[Reg.scala 27:20]
  wire [1:0] _T_24022 = _T_23527 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24277 = _T_24276 | _T_24022; // @[Mux.scala 27:72]
  wire  _T_23529 = bht_rd_addr_hashed_p1_f == 8'h12; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_18; // @[Reg.scala 27:20]
  wire [1:0] _T_24023 = _T_23529 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24278 = _T_24277 | _T_24023; // @[Mux.scala 27:72]
  wire  _T_23531 = bht_rd_addr_hashed_p1_f == 8'h13; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_19; // @[Reg.scala 27:20]
  wire [1:0] _T_24024 = _T_23531 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24279 = _T_24278 | _T_24024; // @[Mux.scala 27:72]
  wire  _T_23533 = bht_rd_addr_hashed_p1_f == 8'h14; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_20; // @[Reg.scala 27:20]
  wire [1:0] _T_24025 = _T_23533 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24280 = _T_24279 | _T_24025; // @[Mux.scala 27:72]
  wire  _T_23535 = bht_rd_addr_hashed_p1_f == 8'h15; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_21; // @[Reg.scala 27:20]
  wire [1:0] _T_24026 = _T_23535 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24281 = _T_24280 | _T_24026; // @[Mux.scala 27:72]
  wire  _T_23537 = bht_rd_addr_hashed_p1_f == 8'h16; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_22; // @[Reg.scala 27:20]
  wire [1:0] _T_24027 = _T_23537 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24282 = _T_24281 | _T_24027; // @[Mux.scala 27:72]
  wire  _T_23539 = bht_rd_addr_hashed_p1_f == 8'h17; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_23; // @[Reg.scala 27:20]
  wire [1:0] _T_24028 = _T_23539 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24283 = _T_24282 | _T_24028; // @[Mux.scala 27:72]
  wire  _T_23541 = bht_rd_addr_hashed_p1_f == 8'h18; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_24; // @[Reg.scala 27:20]
  wire [1:0] _T_24029 = _T_23541 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24284 = _T_24283 | _T_24029; // @[Mux.scala 27:72]
  wire  _T_23543 = bht_rd_addr_hashed_p1_f == 8'h19; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_25; // @[Reg.scala 27:20]
  wire [1:0] _T_24030 = _T_23543 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24285 = _T_24284 | _T_24030; // @[Mux.scala 27:72]
  wire  _T_23545 = bht_rd_addr_hashed_p1_f == 8'h1a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_26; // @[Reg.scala 27:20]
  wire [1:0] _T_24031 = _T_23545 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24286 = _T_24285 | _T_24031; // @[Mux.scala 27:72]
  wire  _T_23547 = bht_rd_addr_hashed_p1_f == 8'h1b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_27; // @[Reg.scala 27:20]
  wire [1:0] _T_24032 = _T_23547 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24287 = _T_24286 | _T_24032; // @[Mux.scala 27:72]
  wire  _T_23549 = bht_rd_addr_hashed_p1_f == 8'h1c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_28; // @[Reg.scala 27:20]
  wire [1:0] _T_24033 = _T_23549 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24288 = _T_24287 | _T_24033; // @[Mux.scala 27:72]
  wire  _T_23551 = bht_rd_addr_hashed_p1_f == 8'h1d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_29; // @[Reg.scala 27:20]
  wire [1:0] _T_24034 = _T_23551 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24289 = _T_24288 | _T_24034; // @[Mux.scala 27:72]
  wire  _T_23553 = bht_rd_addr_hashed_p1_f == 8'h1e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_30; // @[Reg.scala 27:20]
  wire [1:0] _T_24035 = _T_23553 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24290 = _T_24289 | _T_24035; // @[Mux.scala 27:72]
  wire  _T_23555 = bht_rd_addr_hashed_p1_f == 8'h1f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_31; // @[Reg.scala 27:20]
  wire [1:0] _T_24036 = _T_23555 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24291 = _T_24290 | _T_24036; // @[Mux.scala 27:72]
  wire  _T_23557 = bht_rd_addr_hashed_p1_f == 8'h20; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_32; // @[Reg.scala 27:20]
  wire [1:0] _T_24037 = _T_23557 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24292 = _T_24291 | _T_24037; // @[Mux.scala 27:72]
  wire  _T_23559 = bht_rd_addr_hashed_p1_f == 8'h21; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_33; // @[Reg.scala 27:20]
  wire [1:0] _T_24038 = _T_23559 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24293 = _T_24292 | _T_24038; // @[Mux.scala 27:72]
  wire  _T_23561 = bht_rd_addr_hashed_p1_f == 8'h22; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_34; // @[Reg.scala 27:20]
  wire [1:0] _T_24039 = _T_23561 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24294 = _T_24293 | _T_24039; // @[Mux.scala 27:72]
  wire  _T_23563 = bht_rd_addr_hashed_p1_f == 8'h23; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_35; // @[Reg.scala 27:20]
  wire [1:0] _T_24040 = _T_23563 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24295 = _T_24294 | _T_24040; // @[Mux.scala 27:72]
  wire  _T_23565 = bht_rd_addr_hashed_p1_f == 8'h24; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_36; // @[Reg.scala 27:20]
  wire [1:0] _T_24041 = _T_23565 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24296 = _T_24295 | _T_24041; // @[Mux.scala 27:72]
  wire  _T_23567 = bht_rd_addr_hashed_p1_f == 8'h25; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_37; // @[Reg.scala 27:20]
  wire [1:0] _T_24042 = _T_23567 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24297 = _T_24296 | _T_24042; // @[Mux.scala 27:72]
  wire  _T_23569 = bht_rd_addr_hashed_p1_f == 8'h26; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_38; // @[Reg.scala 27:20]
  wire [1:0] _T_24043 = _T_23569 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24298 = _T_24297 | _T_24043; // @[Mux.scala 27:72]
  wire  _T_23571 = bht_rd_addr_hashed_p1_f == 8'h27; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_39; // @[Reg.scala 27:20]
  wire [1:0] _T_24044 = _T_23571 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24299 = _T_24298 | _T_24044; // @[Mux.scala 27:72]
  wire  _T_23573 = bht_rd_addr_hashed_p1_f == 8'h28; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_40; // @[Reg.scala 27:20]
  wire [1:0] _T_24045 = _T_23573 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24300 = _T_24299 | _T_24045; // @[Mux.scala 27:72]
  wire  _T_23575 = bht_rd_addr_hashed_p1_f == 8'h29; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_41; // @[Reg.scala 27:20]
  wire [1:0] _T_24046 = _T_23575 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24301 = _T_24300 | _T_24046; // @[Mux.scala 27:72]
  wire  _T_23577 = bht_rd_addr_hashed_p1_f == 8'h2a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_42; // @[Reg.scala 27:20]
  wire [1:0] _T_24047 = _T_23577 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24302 = _T_24301 | _T_24047; // @[Mux.scala 27:72]
  wire  _T_23579 = bht_rd_addr_hashed_p1_f == 8'h2b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_43; // @[Reg.scala 27:20]
  wire [1:0] _T_24048 = _T_23579 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24303 = _T_24302 | _T_24048; // @[Mux.scala 27:72]
  wire  _T_23581 = bht_rd_addr_hashed_p1_f == 8'h2c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_44; // @[Reg.scala 27:20]
  wire [1:0] _T_24049 = _T_23581 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24304 = _T_24303 | _T_24049; // @[Mux.scala 27:72]
  wire  _T_23583 = bht_rd_addr_hashed_p1_f == 8'h2d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_45; // @[Reg.scala 27:20]
  wire [1:0] _T_24050 = _T_23583 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24305 = _T_24304 | _T_24050; // @[Mux.scala 27:72]
  wire  _T_23585 = bht_rd_addr_hashed_p1_f == 8'h2e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_46; // @[Reg.scala 27:20]
  wire [1:0] _T_24051 = _T_23585 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24306 = _T_24305 | _T_24051; // @[Mux.scala 27:72]
  wire  _T_23587 = bht_rd_addr_hashed_p1_f == 8'h2f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_47; // @[Reg.scala 27:20]
  wire [1:0] _T_24052 = _T_23587 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24307 = _T_24306 | _T_24052; // @[Mux.scala 27:72]
  wire  _T_23589 = bht_rd_addr_hashed_p1_f == 8'h30; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_48; // @[Reg.scala 27:20]
  wire [1:0] _T_24053 = _T_23589 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24308 = _T_24307 | _T_24053; // @[Mux.scala 27:72]
  wire  _T_23591 = bht_rd_addr_hashed_p1_f == 8'h31; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_49; // @[Reg.scala 27:20]
  wire [1:0] _T_24054 = _T_23591 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24309 = _T_24308 | _T_24054; // @[Mux.scala 27:72]
  wire  _T_23593 = bht_rd_addr_hashed_p1_f == 8'h32; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_50; // @[Reg.scala 27:20]
  wire [1:0] _T_24055 = _T_23593 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24310 = _T_24309 | _T_24055; // @[Mux.scala 27:72]
  wire  _T_23595 = bht_rd_addr_hashed_p1_f == 8'h33; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_51; // @[Reg.scala 27:20]
  wire [1:0] _T_24056 = _T_23595 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24311 = _T_24310 | _T_24056; // @[Mux.scala 27:72]
  wire  _T_23597 = bht_rd_addr_hashed_p1_f == 8'h34; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_52; // @[Reg.scala 27:20]
  wire [1:0] _T_24057 = _T_23597 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24312 = _T_24311 | _T_24057; // @[Mux.scala 27:72]
  wire  _T_23599 = bht_rd_addr_hashed_p1_f == 8'h35; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_53; // @[Reg.scala 27:20]
  wire [1:0] _T_24058 = _T_23599 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24313 = _T_24312 | _T_24058; // @[Mux.scala 27:72]
  wire  _T_23601 = bht_rd_addr_hashed_p1_f == 8'h36; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_54; // @[Reg.scala 27:20]
  wire [1:0] _T_24059 = _T_23601 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24314 = _T_24313 | _T_24059; // @[Mux.scala 27:72]
  wire  _T_23603 = bht_rd_addr_hashed_p1_f == 8'h37; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_55; // @[Reg.scala 27:20]
  wire [1:0] _T_24060 = _T_23603 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24315 = _T_24314 | _T_24060; // @[Mux.scala 27:72]
  wire  _T_23605 = bht_rd_addr_hashed_p1_f == 8'h38; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_56; // @[Reg.scala 27:20]
  wire [1:0] _T_24061 = _T_23605 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24316 = _T_24315 | _T_24061; // @[Mux.scala 27:72]
  wire  _T_23607 = bht_rd_addr_hashed_p1_f == 8'h39; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_57; // @[Reg.scala 27:20]
  wire [1:0] _T_24062 = _T_23607 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24317 = _T_24316 | _T_24062; // @[Mux.scala 27:72]
  wire  _T_23609 = bht_rd_addr_hashed_p1_f == 8'h3a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_58; // @[Reg.scala 27:20]
  wire [1:0] _T_24063 = _T_23609 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24318 = _T_24317 | _T_24063; // @[Mux.scala 27:72]
  wire  _T_23611 = bht_rd_addr_hashed_p1_f == 8'h3b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_59; // @[Reg.scala 27:20]
  wire [1:0] _T_24064 = _T_23611 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24319 = _T_24318 | _T_24064; // @[Mux.scala 27:72]
  wire  _T_23613 = bht_rd_addr_hashed_p1_f == 8'h3c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_60; // @[Reg.scala 27:20]
  wire [1:0] _T_24065 = _T_23613 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24320 = _T_24319 | _T_24065; // @[Mux.scala 27:72]
  wire  _T_23615 = bht_rd_addr_hashed_p1_f == 8'h3d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_61; // @[Reg.scala 27:20]
  wire [1:0] _T_24066 = _T_23615 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24321 = _T_24320 | _T_24066; // @[Mux.scala 27:72]
  wire  _T_23617 = bht_rd_addr_hashed_p1_f == 8'h3e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_62; // @[Reg.scala 27:20]
  wire [1:0] _T_24067 = _T_23617 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24322 = _T_24321 | _T_24067; // @[Mux.scala 27:72]
  wire  _T_23619 = bht_rd_addr_hashed_p1_f == 8'h3f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_63; // @[Reg.scala 27:20]
  wire [1:0] _T_24068 = _T_23619 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24323 = _T_24322 | _T_24068; // @[Mux.scala 27:72]
  wire  _T_23621 = bht_rd_addr_hashed_p1_f == 8'h40; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_64; // @[Reg.scala 27:20]
  wire [1:0] _T_24069 = _T_23621 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24324 = _T_24323 | _T_24069; // @[Mux.scala 27:72]
  wire  _T_23623 = bht_rd_addr_hashed_p1_f == 8'h41; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_65; // @[Reg.scala 27:20]
  wire [1:0] _T_24070 = _T_23623 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24325 = _T_24324 | _T_24070; // @[Mux.scala 27:72]
  wire  _T_23625 = bht_rd_addr_hashed_p1_f == 8'h42; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_66; // @[Reg.scala 27:20]
  wire [1:0] _T_24071 = _T_23625 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24326 = _T_24325 | _T_24071; // @[Mux.scala 27:72]
  wire  _T_23627 = bht_rd_addr_hashed_p1_f == 8'h43; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_67; // @[Reg.scala 27:20]
  wire [1:0] _T_24072 = _T_23627 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24327 = _T_24326 | _T_24072; // @[Mux.scala 27:72]
  wire  _T_23629 = bht_rd_addr_hashed_p1_f == 8'h44; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_68; // @[Reg.scala 27:20]
  wire [1:0] _T_24073 = _T_23629 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24328 = _T_24327 | _T_24073; // @[Mux.scala 27:72]
  wire  _T_23631 = bht_rd_addr_hashed_p1_f == 8'h45; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_69; // @[Reg.scala 27:20]
  wire [1:0] _T_24074 = _T_23631 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24329 = _T_24328 | _T_24074; // @[Mux.scala 27:72]
  wire  _T_23633 = bht_rd_addr_hashed_p1_f == 8'h46; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_70; // @[Reg.scala 27:20]
  wire [1:0] _T_24075 = _T_23633 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24330 = _T_24329 | _T_24075; // @[Mux.scala 27:72]
  wire  _T_23635 = bht_rd_addr_hashed_p1_f == 8'h47; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_71; // @[Reg.scala 27:20]
  wire [1:0] _T_24076 = _T_23635 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24331 = _T_24330 | _T_24076; // @[Mux.scala 27:72]
  wire  _T_23637 = bht_rd_addr_hashed_p1_f == 8'h48; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_72; // @[Reg.scala 27:20]
  wire [1:0] _T_24077 = _T_23637 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24332 = _T_24331 | _T_24077; // @[Mux.scala 27:72]
  wire  _T_23639 = bht_rd_addr_hashed_p1_f == 8'h49; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_73; // @[Reg.scala 27:20]
  wire [1:0] _T_24078 = _T_23639 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24333 = _T_24332 | _T_24078; // @[Mux.scala 27:72]
  wire  _T_23641 = bht_rd_addr_hashed_p1_f == 8'h4a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_74; // @[Reg.scala 27:20]
  wire [1:0] _T_24079 = _T_23641 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24334 = _T_24333 | _T_24079; // @[Mux.scala 27:72]
  wire  _T_23643 = bht_rd_addr_hashed_p1_f == 8'h4b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_75; // @[Reg.scala 27:20]
  wire [1:0] _T_24080 = _T_23643 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24335 = _T_24334 | _T_24080; // @[Mux.scala 27:72]
  wire  _T_23645 = bht_rd_addr_hashed_p1_f == 8'h4c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_76; // @[Reg.scala 27:20]
  wire [1:0] _T_24081 = _T_23645 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24336 = _T_24335 | _T_24081; // @[Mux.scala 27:72]
  wire  _T_23647 = bht_rd_addr_hashed_p1_f == 8'h4d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_77; // @[Reg.scala 27:20]
  wire [1:0] _T_24082 = _T_23647 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24337 = _T_24336 | _T_24082; // @[Mux.scala 27:72]
  wire  _T_23649 = bht_rd_addr_hashed_p1_f == 8'h4e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_78; // @[Reg.scala 27:20]
  wire [1:0] _T_24083 = _T_23649 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24338 = _T_24337 | _T_24083; // @[Mux.scala 27:72]
  wire  _T_23651 = bht_rd_addr_hashed_p1_f == 8'h4f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_79; // @[Reg.scala 27:20]
  wire [1:0] _T_24084 = _T_23651 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24339 = _T_24338 | _T_24084; // @[Mux.scala 27:72]
  wire  _T_23653 = bht_rd_addr_hashed_p1_f == 8'h50; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_80; // @[Reg.scala 27:20]
  wire [1:0] _T_24085 = _T_23653 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24340 = _T_24339 | _T_24085; // @[Mux.scala 27:72]
  wire  _T_23655 = bht_rd_addr_hashed_p1_f == 8'h51; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_81; // @[Reg.scala 27:20]
  wire [1:0] _T_24086 = _T_23655 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24341 = _T_24340 | _T_24086; // @[Mux.scala 27:72]
  wire  _T_23657 = bht_rd_addr_hashed_p1_f == 8'h52; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_82; // @[Reg.scala 27:20]
  wire [1:0] _T_24087 = _T_23657 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24342 = _T_24341 | _T_24087; // @[Mux.scala 27:72]
  wire  _T_23659 = bht_rd_addr_hashed_p1_f == 8'h53; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_83; // @[Reg.scala 27:20]
  wire [1:0] _T_24088 = _T_23659 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24343 = _T_24342 | _T_24088; // @[Mux.scala 27:72]
  wire  _T_23661 = bht_rd_addr_hashed_p1_f == 8'h54; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_84; // @[Reg.scala 27:20]
  wire [1:0] _T_24089 = _T_23661 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24344 = _T_24343 | _T_24089; // @[Mux.scala 27:72]
  wire  _T_23663 = bht_rd_addr_hashed_p1_f == 8'h55; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_85; // @[Reg.scala 27:20]
  wire [1:0] _T_24090 = _T_23663 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24345 = _T_24344 | _T_24090; // @[Mux.scala 27:72]
  wire  _T_23665 = bht_rd_addr_hashed_p1_f == 8'h56; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_86; // @[Reg.scala 27:20]
  wire [1:0] _T_24091 = _T_23665 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24346 = _T_24345 | _T_24091; // @[Mux.scala 27:72]
  wire  _T_23667 = bht_rd_addr_hashed_p1_f == 8'h57; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_87; // @[Reg.scala 27:20]
  wire [1:0] _T_24092 = _T_23667 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24347 = _T_24346 | _T_24092; // @[Mux.scala 27:72]
  wire  _T_23669 = bht_rd_addr_hashed_p1_f == 8'h58; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_88; // @[Reg.scala 27:20]
  wire [1:0] _T_24093 = _T_23669 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24348 = _T_24347 | _T_24093; // @[Mux.scala 27:72]
  wire  _T_23671 = bht_rd_addr_hashed_p1_f == 8'h59; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_89; // @[Reg.scala 27:20]
  wire [1:0] _T_24094 = _T_23671 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24349 = _T_24348 | _T_24094; // @[Mux.scala 27:72]
  wire  _T_23673 = bht_rd_addr_hashed_p1_f == 8'h5a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_90; // @[Reg.scala 27:20]
  wire [1:0] _T_24095 = _T_23673 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24350 = _T_24349 | _T_24095; // @[Mux.scala 27:72]
  wire  _T_23675 = bht_rd_addr_hashed_p1_f == 8'h5b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_91; // @[Reg.scala 27:20]
  wire [1:0] _T_24096 = _T_23675 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24351 = _T_24350 | _T_24096; // @[Mux.scala 27:72]
  wire  _T_23677 = bht_rd_addr_hashed_p1_f == 8'h5c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_92; // @[Reg.scala 27:20]
  wire [1:0] _T_24097 = _T_23677 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24352 = _T_24351 | _T_24097; // @[Mux.scala 27:72]
  wire  _T_23679 = bht_rd_addr_hashed_p1_f == 8'h5d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_93; // @[Reg.scala 27:20]
  wire [1:0] _T_24098 = _T_23679 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24353 = _T_24352 | _T_24098; // @[Mux.scala 27:72]
  wire  _T_23681 = bht_rd_addr_hashed_p1_f == 8'h5e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_94; // @[Reg.scala 27:20]
  wire [1:0] _T_24099 = _T_23681 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24354 = _T_24353 | _T_24099; // @[Mux.scala 27:72]
  wire  _T_23683 = bht_rd_addr_hashed_p1_f == 8'h5f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_95; // @[Reg.scala 27:20]
  wire [1:0] _T_24100 = _T_23683 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24355 = _T_24354 | _T_24100; // @[Mux.scala 27:72]
  wire  _T_23685 = bht_rd_addr_hashed_p1_f == 8'h60; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_96; // @[Reg.scala 27:20]
  wire [1:0] _T_24101 = _T_23685 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24356 = _T_24355 | _T_24101; // @[Mux.scala 27:72]
  wire  _T_23687 = bht_rd_addr_hashed_p1_f == 8'h61; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_97; // @[Reg.scala 27:20]
  wire [1:0] _T_24102 = _T_23687 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24357 = _T_24356 | _T_24102; // @[Mux.scala 27:72]
  wire  _T_23689 = bht_rd_addr_hashed_p1_f == 8'h62; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_98; // @[Reg.scala 27:20]
  wire [1:0] _T_24103 = _T_23689 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24358 = _T_24357 | _T_24103; // @[Mux.scala 27:72]
  wire  _T_23691 = bht_rd_addr_hashed_p1_f == 8'h63; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_99; // @[Reg.scala 27:20]
  wire [1:0] _T_24104 = _T_23691 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24359 = _T_24358 | _T_24104; // @[Mux.scala 27:72]
  wire  _T_23693 = bht_rd_addr_hashed_p1_f == 8'h64; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_100; // @[Reg.scala 27:20]
  wire [1:0] _T_24105 = _T_23693 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24360 = _T_24359 | _T_24105; // @[Mux.scala 27:72]
  wire  _T_23695 = bht_rd_addr_hashed_p1_f == 8'h65; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_101; // @[Reg.scala 27:20]
  wire [1:0] _T_24106 = _T_23695 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24361 = _T_24360 | _T_24106; // @[Mux.scala 27:72]
  wire  _T_23697 = bht_rd_addr_hashed_p1_f == 8'h66; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_102; // @[Reg.scala 27:20]
  wire [1:0] _T_24107 = _T_23697 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24362 = _T_24361 | _T_24107; // @[Mux.scala 27:72]
  wire  _T_23699 = bht_rd_addr_hashed_p1_f == 8'h67; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_103; // @[Reg.scala 27:20]
  wire [1:0] _T_24108 = _T_23699 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24363 = _T_24362 | _T_24108; // @[Mux.scala 27:72]
  wire  _T_23701 = bht_rd_addr_hashed_p1_f == 8'h68; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_104; // @[Reg.scala 27:20]
  wire [1:0] _T_24109 = _T_23701 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24364 = _T_24363 | _T_24109; // @[Mux.scala 27:72]
  wire  _T_23703 = bht_rd_addr_hashed_p1_f == 8'h69; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_105; // @[Reg.scala 27:20]
  wire [1:0] _T_24110 = _T_23703 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24365 = _T_24364 | _T_24110; // @[Mux.scala 27:72]
  wire  _T_23705 = bht_rd_addr_hashed_p1_f == 8'h6a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_106; // @[Reg.scala 27:20]
  wire [1:0] _T_24111 = _T_23705 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24366 = _T_24365 | _T_24111; // @[Mux.scala 27:72]
  wire  _T_23707 = bht_rd_addr_hashed_p1_f == 8'h6b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_107; // @[Reg.scala 27:20]
  wire [1:0] _T_24112 = _T_23707 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24367 = _T_24366 | _T_24112; // @[Mux.scala 27:72]
  wire  _T_23709 = bht_rd_addr_hashed_p1_f == 8'h6c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_108; // @[Reg.scala 27:20]
  wire [1:0] _T_24113 = _T_23709 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24368 = _T_24367 | _T_24113; // @[Mux.scala 27:72]
  wire  _T_23711 = bht_rd_addr_hashed_p1_f == 8'h6d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_109; // @[Reg.scala 27:20]
  wire [1:0] _T_24114 = _T_23711 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24369 = _T_24368 | _T_24114; // @[Mux.scala 27:72]
  wire  _T_23713 = bht_rd_addr_hashed_p1_f == 8'h6e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_110; // @[Reg.scala 27:20]
  wire [1:0] _T_24115 = _T_23713 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24370 = _T_24369 | _T_24115; // @[Mux.scala 27:72]
  wire  _T_23715 = bht_rd_addr_hashed_p1_f == 8'h6f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_111; // @[Reg.scala 27:20]
  wire [1:0] _T_24116 = _T_23715 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24371 = _T_24370 | _T_24116; // @[Mux.scala 27:72]
  wire  _T_23717 = bht_rd_addr_hashed_p1_f == 8'h70; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_112; // @[Reg.scala 27:20]
  wire [1:0] _T_24117 = _T_23717 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24372 = _T_24371 | _T_24117; // @[Mux.scala 27:72]
  wire  _T_23719 = bht_rd_addr_hashed_p1_f == 8'h71; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_113; // @[Reg.scala 27:20]
  wire [1:0] _T_24118 = _T_23719 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24373 = _T_24372 | _T_24118; // @[Mux.scala 27:72]
  wire  _T_23721 = bht_rd_addr_hashed_p1_f == 8'h72; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_114; // @[Reg.scala 27:20]
  wire [1:0] _T_24119 = _T_23721 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24374 = _T_24373 | _T_24119; // @[Mux.scala 27:72]
  wire  _T_23723 = bht_rd_addr_hashed_p1_f == 8'h73; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_115; // @[Reg.scala 27:20]
  wire [1:0] _T_24120 = _T_23723 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24375 = _T_24374 | _T_24120; // @[Mux.scala 27:72]
  wire  _T_23725 = bht_rd_addr_hashed_p1_f == 8'h74; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_116; // @[Reg.scala 27:20]
  wire [1:0] _T_24121 = _T_23725 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24376 = _T_24375 | _T_24121; // @[Mux.scala 27:72]
  wire  _T_23727 = bht_rd_addr_hashed_p1_f == 8'h75; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_117; // @[Reg.scala 27:20]
  wire [1:0] _T_24122 = _T_23727 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24377 = _T_24376 | _T_24122; // @[Mux.scala 27:72]
  wire  _T_23729 = bht_rd_addr_hashed_p1_f == 8'h76; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_118; // @[Reg.scala 27:20]
  wire [1:0] _T_24123 = _T_23729 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24378 = _T_24377 | _T_24123; // @[Mux.scala 27:72]
  wire  _T_23731 = bht_rd_addr_hashed_p1_f == 8'h77; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_119; // @[Reg.scala 27:20]
  wire [1:0] _T_24124 = _T_23731 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24379 = _T_24378 | _T_24124; // @[Mux.scala 27:72]
  wire  _T_23733 = bht_rd_addr_hashed_p1_f == 8'h78; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_120; // @[Reg.scala 27:20]
  wire [1:0] _T_24125 = _T_23733 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24380 = _T_24379 | _T_24125; // @[Mux.scala 27:72]
  wire  _T_23735 = bht_rd_addr_hashed_p1_f == 8'h79; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_121; // @[Reg.scala 27:20]
  wire [1:0] _T_24126 = _T_23735 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24381 = _T_24380 | _T_24126; // @[Mux.scala 27:72]
  wire  _T_23737 = bht_rd_addr_hashed_p1_f == 8'h7a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_122; // @[Reg.scala 27:20]
  wire [1:0] _T_24127 = _T_23737 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24382 = _T_24381 | _T_24127; // @[Mux.scala 27:72]
  wire  _T_23739 = bht_rd_addr_hashed_p1_f == 8'h7b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_123; // @[Reg.scala 27:20]
  wire [1:0] _T_24128 = _T_23739 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24383 = _T_24382 | _T_24128; // @[Mux.scala 27:72]
  wire  _T_23741 = bht_rd_addr_hashed_p1_f == 8'h7c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_124; // @[Reg.scala 27:20]
  wire [1:0] _T_24129 = _T_23741 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24384 = _T_24383 | _T_24129; // @[Mux.scala 27:72]
  wire  _T_23743 = bht_rd_addr_hashed_p1_f == 8'h7d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_125; // @[Reg.scala 27:20]
  wire [1:0] _T_24130 = _T_23743 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24385 = _T_24384 | _T_24130; // @[Mux.scala 27:72]
  wire  _T_23745 = bht_rd_addr_hashed_p1_f == 8'h7e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_126; // @[Reg.scala 27:20]
  wire [1:0] _T_24131 = _T_23745 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24386 = _T_24385 | _T_24131; // @[Mux.scala 27:72]
  wire  _T_23747 = bht_rd_addr_hashed_p1_f == 8'h7f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_127; // @[Reg.scala 27:20]
  wire [1:0] _T_24132 = _T_23747 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24387 = _T_24386 | _T_24132; // @[Mux.scala 27:72]
  wire  _T_23749 = bht_rd_addr_hashed_p1_f == 8'h80; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_128; // @[Reg.scala 27:20]
  wire [1:0] _T_24133 = _T_23749 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24388 = _T_24387 | _T_24133; // @[Mux.scala 27:72]
  wire  _T_23751 = bht_rd_addr_hashed_p1_f == 8'h81; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_129; // @[Reg.scala 27:20]
  wire [1:0] _T_24134 = _T_23751 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24389 = _T_24388 | _T_24134; // @[Mux.scala 27:72]
  wire  _T_23753 = bht_rd_addr_hashed_p1_f == 8'h82; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_130; // @[Reg.scala 27:20]
  wire [1:0] _T_24135 = _T_23753 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24390 = _T_24389 | _T_24135; // @[Mux.scala 27:72]
  wire  _T_23755 = bht_rd_addr_hashed_p1_f == 8'h83; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_131; // @[Reg.scala 27:20]
  wire [1:0] _T_24136 = _T_23755 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24391 = _T_24390 | _T_24136; // @[Mux.scala 27:72]
  wire  _T_23757 = bht_rd_addr_hashed_p1_f == 8'h84; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_132; // @[Reg.scala 27:20]
  wire [1:0] _T_24137 = _T_23757 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24392 = _T_24391 | _T_24137; // @[Mux.scala 27:72]
  wire  _T_23759 = bht_rd_addr_hashed_p1_f == 8'h85; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_133; // @[Reg.scala 27:20]
  wire [1:0] _T_24138 = _T_23759 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24393 = _T_24392 | _T_24138; // @[Mux.scala 27:72]
  wire  _T_23761 = bht_rd_addr_hashed_p1_f == 8'h86; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_134; // @[Reg.scala 27:20]
  wire [1:0] _T_24139 = _T_23761 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24394 = _T_24393 | _T_24139; // @[Mux.scala 27:72]
  wire  _T_23763 = bht_rd_addr_hashed_p1_f == 8'h87; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_135; // @[Reg.scala 27:20]
  wire [1:0] _T_24140 = _T_23763 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24395 = _T_24394 | _T_24140; // @[Mux.scala 27:72]
  wire  _T_23765 = bht_rd_addr_hashed_p1_f == 8'h88; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_136; // @[Reg.scala 27:20]
  wire [1:0] _T_24141 = _T_23765 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24396 = _T_24395 | _T_24141; // @[Mux.scala 27:72]
  wire  _T_23767 = bht_rd_addr_hashed_p1_f == 8'h89; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_137; // @[Reg.scala 27:20]
  wire [1:0] _T_24142 = _T_23767 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24397 = _T_24396 | _T_24142; // @[Mux.scala 27:72]
  wire  _T_23769 = bht_rd_addr_hashed_p1_f == 8'h8a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_138; // @[Reg.scala 27:20]
  wire [1:0] _T_24143 = _T_23769 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24398 = _T_24397 | _T_24143; // @[Mux.scala 27:72]
  wire  _T_23771 = bht_rd_addr_hashed_p1_f == 8'h8b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_139; // @[Reg.scala 27:20]
  wire [1:0] _T_24144 = _T_23771 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24399 = _T_24398 | _T_24144; // @[Mux.scala 27:72]
  wire  _T_23773 = bht_rd_addr_hashed_p1_f == 8'h8c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_140; // @[Reg.scala 27:20]
  wire [1:0] _T_24145 = _T_23773 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24400 = _T_24399 | _T_24145; // @[Mux.scala 27:72]
  wire  _T_23775 = bht_rd_addr_hashed_p1_f == 8'h8d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_141; // @[Reg.scala 27:20]
  wire [1:0] _T_24146 = _T_23775 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24401 = _T_24400 | _T_24146; // @[Mux.scala 27:72]
  wire  _T_23777 = bht_rd_addr_hashed_p1_f == 8'h8e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_142; // @[Reg.scala 27:20]
  wire [1:0] _T_24147 = _T_23777 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24402 = _T_24401 | _T_24147; // @[Mux.scala 27:72]
  wire  _T_23779 = bht_rd_addr_hashed_p1_f == 8'h8f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_143; // @[Reg.scala 27:20]
  wire [1:0] _T_24148 = _T_23779 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24403 = _T_24402 | _T_24148; // @[Mux.scala 27:72]
  wire  _T_23781 = bht_rd_addr_hashed_p1_f == 8'h90; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_144; // @[Reg.scala 27:20]
  wire [1:0] _T_24149 = _T_23781 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24404 = _T_24403 | _T_24149; // @[Mux.scala 27:72]
  wire  _T_23783 = bht_rd_addr_hashed_p1_f == 8'h91; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_145; // @[Reg.scala 27:20]
  wire [1:0] _T_24150 = _T_23783 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24405 = _T_24404 | _T_24150; // @[Mux.scala 27:72]
  wire  _T_23785 = bht_rd_addr_hashed_p1_f == 8'h92; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_146; // @[Reg.scala 27:20]
  wire [1:0] _T_24151 = _T_23785 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24406 = _T_24405 | _T_24151; // @[Mux.scala 27:72]
  wire  _T_23787 = bht_rd_addr_hashed_p1_f == 8'h93; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_147; // @[Reg.scala 27:20]
  wire [1:0] _T_24152 = _T_23787 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24407 = _T_24406 | _T_24152; // @[Mux.scala 27:72]
  wire  _T_23789 = bht_rd_addr_hashed_p1_f == 8'h94; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_148; // @[Reg.scala 27:20]
  wire [1:0] _T_24153 = _T_23789 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24408 = _T_24407 | _T_24153; // @[Mux.scala 27:72]
  wire  _T_23791 = bht_rd_addr_hashed_p1_f == 8'h95; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_149; // @[Reg.scala 27:20]
  wire [1:0] _T_24154 = _T_23791 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24409 = _T_24408 | _T_24154; // @[Mux.scala 27:72]
  wire  _T_23793 = bht_rd_addr_hashed_p1_f == 8'h96; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_150; // @[Reg.scala 27:20]
  wire [1:0] _T_24155 = _T_23793 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24410 = _T_24409 | _T_24155; // @[Mux.scala 27:72]
  wire  _T_23795 = bht_rd_addr_hashed_p1_f == 8'h97; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_151; // @[Reg.scala 27:20]
  wire [1:0] _T_24156 = _T_23795 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24411 = _T_24410 | _T_24156; // @[Mux.scala 27:72]
  wire  _T_23797 = bht_rd_addr_hashed_p1_f == 8'h98; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_152; // @[Reg.scala 27:20]
  wire [1:0] _T_24157 = _T_23797 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24412 = _T_24411 | _T_24157; // @[Mux.scala 27:72]
  wire  _T_23799 = bht_rd_addr_hashed_p1_f == 8'h99; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_153; // @[Reg.scala 27:20]
  wire [1:0] _T_24158 = _T_23799 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24413 = _T_24412 | _T_24158; // @[Mux.scala 27:72]
  wire  _T_23801 = bht_rd_addr_hashed_p1_f == 8'h9a; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_154; // @[Reg.scala 27:20]
  wire [1:0] _T_24159 = _T_23801 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24414 = _T_24413 | _T_24159; // @[Mux.scala 27:72]
  wire  _T_23803 = bht_rd_addr_hashed_p1_f == 8'h9b; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_155; // @[Reg.scala 27:20]
  wire [1:0] _T_24160 = _T_23803 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24415 = _T_24414 | _T_24160; // @[Mux.scala 27:72]
  wire  _T_23805 = bht_rd_addr_hashed_p1_f == 8'h9c; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_156; // @[Reg.scala 27:20]
  wire [1:0] _T_24161 = _T_23805 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24416 = _T_24415 | _T_24161; // @[Mux.scala 27:72]
  wire  _T_23807 = bht_rd_addr_hashed_p1_f == 8'h9d; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_157; // @[Reg.scala 27:20]
  wire [1:0] _T_24162 = _T_23807 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24417 = _T_24416 | _T_24162; // @[Mux.scala 27:72]
  wire  _T_23809 = bht_rd_addr_hashed_p1_f == 8'h9e; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_158; // @[Reg.scala 27:20]
  wire [1:0] _T_24163 = _T_23809 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24418 = _T_24417 | _T_24163; // @[Mux.scala 27:72]
  wire  _T_23811 = bht_rd_addr_hashed_p1_f == 8'h9f; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_159; // @[Reg.scala 27:20]
  wire [1:0] _T_24164 = _T_23811 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24419 = _T_24418 | _T_24164; // @[Mux.scala 27:72]
  wire  _T_23813 = bht_rd_addr_hashed_p1_f == 8'ha0; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_160; // @[Reg.scala 27:20]
  wire [1:0] _T_24165 = _T_23813 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24420 = _T_24419 | _T_24165; // @[Mux.scala 27:72]
  wire  _T_23815 = bht_rd_addr_hashed_p1_f == 8'ha1; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_161; // @[Reg.scala 27:20]
  wire [1:0] _T_24166 = _T_23815 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24421 = _T_24420 | _T_24166; // @[Mux.scala 27:72]
  wire  _T_23817 = bht_rd_addr_hashed_p1_f == 8'ha2; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_162; // @[Reg.scala 27:20]
  wire [1:0] _T_24167 = _T_23817 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24422 = _T_24421 | _T_24167; // @[Mux.scala 27:72]
  wire  _T_23819 = bht_rd_addr_hashed_p1_f == 8'ha3; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_163; // @[Reg.scala 27:20]
  wire [1:0] _T_24168 = _T_23819 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24423 = _T_24422 | _T_24168; // @[Mux.scala 27:72]
  wire  _T_23821 = bht_rd_addr_hashed_p1_f == 8'ha4; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_164; // @[Reg.scala 27:20]
  wire [1:0] _T_24169 = _T_23821 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24424 = _T_24423 | _T_24169; // @[Mux.scala 27:72]
  wire  _T_23823 = bht_rd_addr_hashed_p1_f == 8'ha5; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_165; // @[Reg.scala 27:20]
  wire [1:0] _T_24170 = _T_23823 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24425 = _T_24424 | _T_24170; // @[Mux.scala 27:72]
  wire  _T_23825 = bht_rd_addr_hashed_p1_f == 8'ha6; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_166; // @[Reg.scala 27:20]
  wire [1:0] _T_24171 = _T_23825 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24426 = _T_24425 | _T_24171; // @[Mux.scala 27:72]
  wire  _T_23827 = bht_rd_addr_hashed_p1_f == 8'ha7; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_167; // @[Reg.scala 27:20]
  wire [1:0] _T_24172 = _T_23827 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24427 = _T_24426 | _T_24172; // @[Mux.scala 27:72]
  wire  _T_23829 = bht_rd_addr_hashed_p1_f == 8'ha8; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_168; // @[Reg.scala 27:20]
  wire [1:0] _T_24173 = _T_23829 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24428 = _T_24427 | _T_24173; // @[Mux.scala 27:72]
  wire  _T_23831 = bht_rd_addr_hashed_p1_f == 8'ha9; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_169; // @[Reg.scala 27:20]
  wire [1:0] _T_24174 = _T_23831 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24429 = _T_24428 | _T_24174; // @[Mux.scala 27:72]
  wire  _T_23833 = bht_rd_addr_hashed_p1_f == 8'haa; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_170; // @[Reg.scala 27:20]
  wire [1:0] _T_24175 = _T_23833 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24430 = _T_24429 | _T_24175; // @[Mux.scala 27:72]
  wire  _T_23835 = bht_rd_addr_hashed_p1_f == 8'hab; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_171; // @[Reg.scala 27:20]
  wire [1:0] _T_24176 = _T_23835 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24431 = _T_24430 | _T_24176; // @[Mux.scala 27:72]
  wire  _T_23837 = bht_rd_addr_hashed_p1_f == 8'hac; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_172; // @[Reg.scala 27:20]
  wire [1:0] _T_24177 = _T_23837 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24432 = _T_24431 | _T_24177; // @[Mux.scala 27:72]
  wire  _T_23839 = bht_rd_addr_hashed_p1_f == 8'had; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_173; // @[Reg.scala 27:20]
  wire [1:0] _T_24178 = _T_23839 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24433 = _T_24432 | _T_24178; // @[Mux.scala 27:72]
  wire  _T_23841 = bht_rd_addr_hashed_p1_f == 8'hae; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_174; // @[Reg.scala 27:20]
  wire [1:0] _T_24179 = _T_23841 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24434 = _T_24433 | _T_24179; // @[Mux.scala 27:72]
  wire  _T_23843 = bht_rd_addr_hashed_p1_f == 8'haf; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_175; // @[Reg.scala 27:20]
  wire [1:0] _T_24180 = _T_23843 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24435 = _T_24434 | _T_24180; // @[Mux.scala 27:72]
  wire  _T_23845 = bht_rd_addr_hashed_p1_f == 8'hb0; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_176; // @[Reg.scala 27:20]
  wire [1:0] _T_24181 = _T_23845 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24436 = _T_24435 | _T_24181; // @[Mux.scala 27:72]
  wire  _T_23847 = bht_rd_addr_hashed_p1_f == 8'hb1; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_177; // @[Reg.scala 27:20]
  wire [1:0] _T_24182 = _T_23847 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24437 = _T_24436 | _T_24182; // @[Mux.scala 27:72]
  wire  _T_23849 = bht_rd_addr_hashed_p1_f == 8'hb2; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_178; // @[Reg.scala 27:20]
  wire [1:0] _T_24183 = _T_23849 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24438 = _T_24437 | _T_24183; // @[Mux.scala 27:72]
  wire  _T_23851 = bht_rd_addr_hashed_p1_f == 8'hb3; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_179; // @[Reg.scala 27:20]
  wire [1:0] _T_24184 = _T_23851 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24439 = _T_24438 | _T_24184; // @[Mux.scala 27:72]
  wire  _T_23853 = bht_rd_addr_hashed_p1_f == 8'hb4; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_180; // @[Reg.scala 27:20]
  wire [1:0] _T_24185 = _T_23853 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24440 = _T_24439 | _T_24185; // @[Mux.scala 27:72]
  wire  _T_23855 = bht_rd_addr_hashed_p1_f == 8'hb5; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_181; // @[Reg.scala 27:20]
  wire [1:0] _T_24186 = _T_23855 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24441 = _T_24440 | _T_24186; // @[Mux.scala 27:72]
  wire  _T_23857 = bht_rd_addr_hashed_p1_f == 8'hb6; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_182; // @[Reg.scala 27:20]
  wire [1:0] _T_24187 = _T_23857 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24442 = _T_24441 | _T_24187; // @[Mux.scala 27:72]
  wire  _T_23859 = bht_rd_addr_hashed_p1_f == 8'hb7; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_183; // @[Reg.scala 27:20]
  wire [1:0] _T_24188 = _T_23859 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24443 = _T_24442 | _T_24188; // @[Mux.scala 27:72]
  wire  _T_23861 = bht_rd_addr_hashed_p1_f == 8'hb8; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_184; // @[Reg.scala 27:20]
  wire [1:0] _T_24189 = _T_23861 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24444 = _T_24443 | _T_24189; // @[Mux.scala 27:72]
  wire  _T_23863 = bht_rd_addr_hashed_p1_f == 8'hb9; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_185; // @[Reg.scala 27:20]
  wire [1:0] _T_24190 = _T_23863 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24445 = _T_24444 | _T_24190; // @[Mux.scala 27:72]
  wire  _T_23865 = bht_rd_addr_hashed_p1_f == 8'hba; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_186; // @[Reg.scala 27:20]
  wire [1:0] _T_24191 = _T_23865 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24446 = _T_24445 | _T_24191; // @[Mux.scala 27:72]
  wire  _T_23867 = bht_rd_addr_hashed_p1_f == 8'hbb; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_187; // @[Reg.scala 27:20]
  wire [1:0] _T_24192 = _T_23867 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24447 = _T_24446 | _T_24192; // @[Mux.scala 27:72]
  wire  _T_23869 = bht_rd_addr_hashed_p1_f == 8'hbc; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_188; // @[Reg.scala 27:20]
  wire [1:0] _T_24193 = _T_23869 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24448 = _T_24447 | _T_24193; // @[Mux.scala 27:72]
  wire  _T_23871 = bht_rd_addr_hashed_p1_f == 8'hbd; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_189; // @[Reg.scala 27:20]
  wire [1:0] _T_24194 = _T_23871 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24449 = _T_24448 | _T_24194; // @[Mux.scala 27:72]
  wire  _T_23873 = bht_rd_addr_hashed_p1_f == 8'hbe; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_190; // @[Reg.scala 27:20]
  wire [1:0] _T_24195 = _T_23873 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24450 = _T_24449 | _T_24195; // @[Mux.scala 27:72]
  wire  _T_23875 = bht_rd_addr_hashed_p1_f == 8'hbf; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_191; // @[Reg.scala 27:20]
  wire [1:0] _T_24196 = _T_23875 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24451 = _T_24450 | _T_24196; // @[Mux.scala 27:72]
  wire  _T_23877 = bht_rd_addr_hashed_p1_f == 8'hc0; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_192; // @[Reg.scala 27:20]
  wire [1:0] _T_24197 = _T_23877 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24452 = _T_24451 | _T_24197; // @[Mux.scala 27:72]
  wire  _T_23879 = bht_rd_addr_hashed_p1_f == 8'hc1; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_193; // @[Reg.scala 27:20]
  wire [1:0] _T_24198 = _T_23879 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24453 = _T_24452 | _T_24198; // @[Mux.scala 27:72]
  wire  _T_23881 = bht_rd_addr_hashed_p1_f == 8'hc2; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_194; // @[Reg.scala 27:20]
  wire [1:0] _T_24199 = _T_23881 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24454 = _T_24453 | _T_24199; // @[Mux.scala 27:72]
  wire  _T_23883 = bht_rd_addr_hashed_p1_f == 8'hc3; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_195; // @[Reg.scala 27:20]
  wire [1:0] _T_24200 = _T_23883 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24455 = _T_24454 | _T_24200; // @[Mux.scala 27:72]
  wire  _T_23885 = bht_rd_addr_hashed_p1_f == 8'hc4; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_196; // @[Reg.scala 27:20]
  wire [1:0] _T_24201 = _T_23885 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24456 = _T_24455 | _T_24201; // @[Mux.scala 27:72]
  wire  _T_23887 = bht_rd_addr_hashed_p1_f == 8'hc5; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_197; // @[Reg.scala 27:20]
  wire [1:0] _T_24202 = _T_23887 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24457 = _T_24456 | _T_24202; // @[Mux.scala 27:72]
  wire  _T_23889 = bht_rd_addr_hashed_p1_f == 8'hc6; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_198; // @[Reg.scala 27:20]
  wire [1:0] _T_24203 = _T_23889 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24458 = _T_24457 | _T_24203; // @[Mux.scala 27:72]
  wire  _T_23891 = bht_rd_addr_hashed_p1_f == 8'hc7; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_199; // @[Reg.scala 27:20]
  wire [1:0] _T_24204 = _T_23891 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24459 = _T_24458 | _T_24204; // @[Mux.scala 27:72]
  wire  _T_23893 = bht_rd_addr_hashed_p1_f == 8'hc8; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_200; // @[Reg.scala 27:20]
  wire [1:0] _T_24205 = _T_23893 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24460 = _T_24459 | _T_24205; // @[Mux.scala 27:72]
  wire  _T_23895 = bht_rd_addr_hashed_p1_f == 8'hc9; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_201; // @[Reg.scala 27:20]
  wire [1:0] _T_24206 = _T_23895 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24461 = _T_24460 | _T_24206; // @[Mux.scala 27:72]
  wire  _T_23897 = bht_rd_addr_hashed_p1_f == 8'hca; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_202; // @[Reg.scala 27:20]
  wire [1:0] _T_24207 = _T_23897 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24462 = _T_24461 | _T_24207; // @[Mux.scala 27:72]
  wire  _T_23899 = bht_rd_addr_hashed_p1_f == 8'hcb; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_203; // @[Reg.scala 27:20]
  wire [1:0] _T_24208 = _T_23899 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24463 = _T_24462 | _T_24208; // @[Mux.scala 27:72]
  wire  _T_23901 = bht_rd_addr_hashed_p1_f == 8'hcc; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_204; // @[Reg.scala 27:20]
  wire [1:0] _T_24209 = _T_23901 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24464 = _T_24463 | _T_24209; // @[Mux.scala 27:72]
  wire  _T_23903 = bht_rd_addr_hashed_p1_f == 8'hcd; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_205; // @[Reg.scala 27:20]
  wire [1:0] _T_24210 = _T_23903 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24465 = _T_24464 | _T_24210; // @[Mux.scala 27:72]
  wire  _T_23905 = bht_rd_addr_hashed_p1_f == 8'hce; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_206; // @[Reg.scala 27:20]
  wire [1:0] _T_24211 = _T_23905 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24466 = _T_24465 | _T_24211; // @[Mux.scala 27:72]
  wire  _T_23907 = bht_rd_addr_hashed_p1_f == 8'hcf; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_207; // @[Reg.scala 27:20]
  wire [1:0] _T_24212 = _T_23907 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24467 = _T_24466 | _T_24212; // @[Mux.scala 27:72]
  wire  _T_23909 = bht_rd_addr_hashed_p1_f == 8'hd0; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_208; // @[Reg.scala 27:20]
  wire [1:0] _T_24213 = _T_23909 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24468 = _T_24467 | _T_24213; // @[Mux.scala 27:72]
  wire  _T_23911 = bht_rd_addr_hashed_p1_f == 8'hd1; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_209; // @[Reg.scala 27:20]
  wire [1:0] _T_24214 = _T_23911 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24469 = _T_24468 | _T_24214; // @[Mux.scala 27:72]
  wire  _T_23913 = bht_rd_addr_hashed_p1_f == 8'hd2; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_210; // @[Reg.scala 27:20]
  wire [1:0] _T_24215 = _T_23913 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24470 = _T_24469 | _T_24215; // @[Mux.scala 27:72]
  wire  _T_23915 = bht_rd_addr_hashed_p1_f == 8'hd3; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_211; // @[Reg.scala 27:20]
  wire [1:0] _T_24216 = _T_23915 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24471 = _T_24470 | _T_24216; // @[Mux.scala 27:72]
  wire  _T_23917 = bht_rd_addr_hashed_p1_f == 8'hd4; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_212; // @[Reg.scala 27:20]
  wire [1:0] _T_24217 = _T_23917 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24472 = _T_24471 | _T_24217; // @[Mux.scala 27:72]
  wire  _T_23919 = bht_rd_addr_hashed_p1_f == 8'hd5; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_213; // @[Reg.scala 27:20]
  wire [1:0] _T_24218 = _T_23919 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24473 = _T_24472 | _T_24218; // @[Mux.scala 27:72]
  wire  _T_23921 = bht_rd_addr_hashed_p1_f == 8'hd6; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_214; // @[Reg.scala 27:20]
  wire [1:0] _T_24219 = _T_23921 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24474 = _T_24473 | _T_24219; // @[Mux.scala 27:72]
  wire  _T_23923 = bht_rd_addr_hashed_p1_f == 8'hd7; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_215; // @[Reg.scala 27:20]
  wire [1:0] _T_24220 = _T_23923 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24475 = _T_24474 | _T_24220; // @[Mux.scala 27:72]
  wire  _T_23925 = bht_rd_addr_hashed_p1_f == 8'hd8; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_216; // @[Reg.scala 27:20]
  wire [1:0] _T_24221 = _T_23925 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24476 = _T_24475 | _T_24221; // @[Mux.scala 27:72]
  wire  _T_23927 = bht_rd_addr_hashed_p1_f == 8'hd9; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_217; // @[Reg.scala 27:20]
  wire [1:0] _T_24222 = _T_23927 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24477 = _T_24476 | _T_24222; // @[Mux.scala 27:72]
  wire  _T_23929 = bht_rd_addr_hashed_p1_f == 8'hda; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_218; // @[Reg.scala 27:20]
  wire [1:0] _T_24223 = _T_23929 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24478 = _T_24477 | _T_24223; // @[Mux.scala 27:72]
  wire  _T_23931 = bht_rd_addr_hashed_p1_f == 8'hdb; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_219; // @[Reg.scala 27:20]
  wire [1:0] _T_24224 = _T_23931 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24479 = _T_24478 | _T_24224; // @[Mux.scala 27:72]
  wire  _T_23933 = bht_rd_addr_hashed_p1_f == 8'hdc; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_220; // @[Reg.scala 27:20]
  wire [1:0] _T_24225 = _T_23933 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24480 = _T_24479 | _T_24225; // @[Mux.scala 27:72]
  wire  _T_23935 = bht_rd_addr_hashed_p1_f == 8'hdd; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_221; // @[Reg.scala 27:20]
  wire [1:0] _T_24226 = _T_23935 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24481 = _T_24480 | _T_24226; // @[Mux.scala 27:72]
  wire  _T_23937 = bht_rd_addr_hashed_p1_f == 8'hde; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_222; // @[Reg.scala 27:20]
  wire [1:0] _T_24227 = _T_23937 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24482 = _T_24481 | _T_24227; // @[Mux.scala 27:72]
  wire  _T_23939 = bht_rd_addr_hashed_p1_f == 8'hdf; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_223; // @[Reg.scala 27:20]
  wire [1:0] _T_24228 = _T_23939 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24483 = _T_24482 | _T_24228; // @[Mux.scala 27:72]
  wire  _T_23941 = bht_rd_addr_hashed_p1_f == 8'he0; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_224; // @[Reg.scala 27:20]
  wire [1:0] _T_24229 = _T_23941 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24484 = _T_24483 | _T_24229; // @[Mux.scala 27:72]
  wire  _T_23943 = bht_rd_addr_hashed_p1_f == 8'he1; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_225; // @[Reg.scala 27:20]
  wire [1:0] _T_24230 = _T_23943 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24485 = _T_24484 | _T_24230; // @[Mux.scala 27:72]
  wire  _T_23945 = bht_rd_addr_hashed_p1_f == 8'he2; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_226; // @[Reg.scala 27:20]
  wire [1:0] _T_24231 = _T_23945 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24486 = _T_24485 | _T_24231; // @[Mux.scala 27:72]
  wire  _T_23947 = bht_rd_addr_hashed_p1_f == 8'he3; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_227; // @[Reg.scala 27:20]
  wire [1:0] _T_24232 = _T_23947 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24487 = _T_24486 | _T_24232; // @[Mux.scala 27:72]
  wire  _T_23949 = bht_rd_addr_hashed_p1_f == 8'he4; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_228; // @[Reg.scala 27:20]
  wire [1:0] _T_24233 = _T_23949 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24488 = _T_24487 | _T_24233; // @[Mux.scala 27:72]
  wire  _T_23951 = bht_rd_addr_hashed_p1_f == 8'he5; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_229; // @[Reg.scala 27:20]
  wire [1:0] _T_24234 = _T_23951 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24489 = _T_24488 | _T_24234; // @[Mux.scala 27:72]
  wire  _T_23953 = bht_rd_addr_hashed_p1_f == 8'he6; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_230; // @[Reg.scala 27:20]
  wire [1:0] _T_24235 = _T_23953 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24490 = _T_24489 | _T_24235; // @[Mux.scala 27:72]
  wire  _T_23955 = bht_rd_addr_hashed_p1_f == 8'he7; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_231; // @[Reg.scala 27:20]
  wire [1:0] _T_24236 = _T_23955 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24491 = _T_24490 | _T_24236; // @[Mux.scala 27:72]
  wire  _T_23957 = bht_rd_addr_hashed_p1_f == 8'he8; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_232; // @[Reg.scala 27:20]
  wire [1:0] _T_24237 = _T_23957 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24492 = _T_24491 | _T_24237; // @[Mux.scala 27:72]
  wire  _T_23959 = bht_rd_addr_hashed_p1_f == 8'he9; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_233; // @[Reg.scala 27:20]
  wire [1:0] _T_24238 = _T_23959 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24493 = _T_24492 | _T_24238; // @[Mux.scala 27:72]
  wire  _T_23961 = bht_rd_addr_hashed_p1_f == 8'hea; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_234; // @[Reg.scala 27:20]
  wire [1:0] _T_24239 = _T_23961 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24494 = _T_24493 | _T_24239; // @[Mux.scala 27:72]
  wire  _T_23963 = bht_rd_addr_hashed_p1_f == 8'heb; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_235; // @[Reg.scala 27:20]
  wire [1:0] _T_24240 = _T_23963 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24495 = _T_24494 | _T_24240; // @[Mux.scala 27:72]
  wire  _T_23965 = bht_rd_addr_hashed_p1_f == 8'hec; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_236; // @[Reg.scala 27:20]
  wire [1:0] _T_24241 = _T_23965 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24496 = _T_24495 | _T_24241; // @[Mux.scala 27:72]
  wire  _T_23967 = bht_rd_addr_hashed_p1_f == 8'hed; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_237; // @[Reg.scala 27:20]
  wire [1:0] _T_24242 = _T_23967 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24497 = _T_24496 | _T_24242; // @[Mux.scala 27:72]
  wire  _T_23969 = bht_rd_addr_hashed_p1_f == 8'hee; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_238; // @[Reg.scala 27:20]
  wire [1:0] _T_24243 = _T_23969 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24498 = _T_24497 | _T_24243; // @[Mux.scala 27:72]
  wire  _T_23971 = bht_rd_addr_hashed_p1_f == 8'hef; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_239; // @[Reg.scala 27:20]
  wire [1:0] _T_24244 = _T_23971 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24499 = _T_24498 | _T_24244; // @[Mux.scala 27:72]
  wire  _T_23973 = bht_rd_addr_hashed_p1_f == 8'hf0; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_240; // @[Reg.scala 27:20]
  wire [1:0] _T_24245 = _T_23973 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24500 = _T_24499 | _T_24245; // @[Mux.scala 27:72]
  wire  _T_23975 = bht_rd_addr_hashed_p1_f == 8'hf1; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_241; // @[Reg.scala 27:20]
  wire [1:0] _T_24246 = _T_23975 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24501 = _T_24500 | _T_24246; // @[Mux.scala 27:72]
  wire  _T_23977 = bht_rd_addr_hashed_p1_f == 8'hf2; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_242; // @[Reg.scala 27:20]
  wire [1:0] _T_24247 = _T_23977 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24502 = _T_24501 | _T_24247; // @[Mux.scala 27:72]
  wire  _T_23979 = bht_rd_addr_hashed_p1_f == 8'hf3; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_243; // @[Reg.scala 27:20]
  wire [1:0] _T_24248 = _T_23979 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24503 = _T_24502 | _T_24248; // @[Mux.scala 27:72]
  wire  _T_23981 = bht_rd_addr_hashed_p1_f == 8'hf4; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_244; // @[Reg.scala 27:20]
  wire [1:0] _T_24249 = _T_23981 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24504 = _T_24503 | _T_24249; // @[Mux.scala 27:72]
  wire  _T_23983 = bht_rd_addr_hashed_p1_f == 8'hf5; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_245; // @[Reg.scala 27:20]
  wire [1:0] _T_24250 = _T_23983 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24505 = _T_24504 | _T_24250; // @[Mux.scala 27:72]
  wire  _T_23985 = bht_rd_addr_hashed_p1_f == 8'hf6; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_246; // @[Reg.scala 27:20]
  wire [1:0] _T_24251 = _T_23985 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24506 = _T_24505 | _T_24251; // @[Mux.scala 27:72]
  wire  _T_23987 = bht_rd_addr_hashed_p1_f == 8'hf7; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_247; // @[Reg.scala 27:20]
  wire [1:0] _T_24252 = _T_23987 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24507 = _T_24506 | _T_24252; // @[Mux.scala 27:72]
  wire  _T_23989 = bht_rd_addr_hashed_p1_f == 8'hf8; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_248; // @[Reg.scala 27:20]
  wire [1:0] _T_24253 = _T_23989 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24508 = _T_24507 | _T_24253; // @[Mux.scala 27:72]
  wire  _T_23991 = bht_rd_addr_hashed_p1_f == 8'hf9; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_249; // @[Reg.scala 27:20]
  wire [1:0] _T_24254 = _T_23991 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24509 = _T_24508 | _T_24254; // @[Mux.scala 27:72]
  wire  _T_23993 = bht_rd_addr_hashed_p1_f == 8'hfa; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_250; // @[Reg.scala 27:20]
  wire [1:0] _T_24255 = _T_23993 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24510 = _T_24509 | _T_24255; // @[Mux.scala 27:72]
  wire  _T_23995 = bht_rd_addr_hashed_p1_f == 8'hfb; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_251; // @[Reg.scala 27:20]
  wire [1:0] _T_24256 = _T_23995 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24511 = _T_24510 | _T_24256; // @[Mux.scala 27:72]
  wire  _T_23997 = bht_rd_addr_hashed_p1_f == 8'hfc; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_252; // @[Reg.scala 27:20]
  wire [1:0] _T_24257 = _T_23997 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24512 = _T_24511 | _T_24257; // @[Mux.scala 27:72]
  wire  _T_23999 = bht_rd_addr_hashed_p1_f == 8'hfd; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_253; // @[Reg.scala 27:20]
  wire [1:0] _T_24258 = _T_23999 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24513 = _T_24512 | _T_24258; // @[Mux.scala 27:72]
  wire  _T_24001 = bht_rd_addr_hashed_p1_f == 8'hfe; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_254; // @[Reg.scala 27:20]
  wire [1:0] _T_24259 = _T_24001 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_24514 = _T_24513 | _T_24259; // @[Mux.scala 27:72]
  wire  _T_24003 = bht_rd_addr_hashed_p1_f == 8'hff; // @[ifu_bp_ctl.scala 532:85]
  reg [1:0] bht_bank_rd_data_out_0_255; // @[Reg.scala 27:20]
  wire [1:0] _T_24260 = _T_24003 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_p1_f = _T_24514 | _T_24260; // @[Mux.scala 27:72]
  wire [1:0] _T_254 = io_ifc_fetch_addr_f[0] ? bht_bank0_rd_data_p1_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank1_rd_data_f = _T_253 | _T_254; // @[Mux.scala 27:72]
  wire  _T_258 = bht_force_taken_f[1] | bht_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 298:42]
  wire [1:0] wayhit_f = tag_match_way0_expanded_f | tag_match_way1_expanded_f; // @[ifu_bp_ctl.scala 172:41]
  wire [1:0] _T_607 = _T_147 ? wayhit_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] wayhit_p1_f = tag_match_way0_expanded_p1_f | tag_match_way1_expanded_p1_f; // @[ifu_bp_ctl.scala 174:47]
  wire [1:0] _T_606 = {wayhit_p1_f[0],wayhit_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_608 = io_ifc_fetch_addr_f[0] ? _T_606 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_609 = _T_607 | _T_608; // @[Mux.scala 27:72]
  wire  eoc_near = &io_ifc_fetch_addr_f[4:2]; // @[ifu_bp_ctl.scala 258:64]
  wire  _T_212 = ~eoc_near; // @[ifu_bp_ctl.scala 260:15]
  wire [1:0] _T_214 = ~io_ifc_fetch_addr_f[1:0]; // @[ifu_bp_ctl.scala 260:28]
  wire  _T_215 = |_T_214; // @[ifu_bp_ctl.scala 260:58]
  wire  eoc_mask = _T_212 | _T_215; // @[ifu_bp_ctl.scala 260:25]
  wire [1:0] _T_611 = {eoc_mask,1'h1}; // @[Cat.scala 29:58]
  wire [1:0] vwayhit_f = _T_609 & _T_611; // @[ifu_bp_ctl.scala 432:71]
  wire  _T_260 = _T_258 & vwayhit_f[1]; // @[ifu_bp_ctl.scala 298:69]
  wire [1:0] _T_21957 = _T_22469 ? bht_bank_rd_data_out_0_0 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_21958 = _T_22471 ? bht_bank_rd_data_out_0_1 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22213 = _T_21957 | _T_21958; // @[Mux.scala 27:72]
  wire [1:0] _T_21959 = _T_22473 ? bht_bank_rd_data_out_0_2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22214 = _T_22213 | _T_21959; // @[Mux.scala 27:72]
  wire [1:0] _T_21960 = _T_22475 ? bht_bank_rd_data_out_0_3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22215 = _T_22214 | _T_21960; // @[Mux.scala 27:72]
  wire [1:0] _T_21961 = _T_22477 ? bht_bank_rd_data_out_0_4 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22216 = _T_22215 | _T_21961; // @[Mux.scala 27:72]
  wire [1:0] _T_21962 = _T_22479 ? bht_bank_rd_data_out_0_5 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22217 = _T_22216 | _T_21962; // @[Mux.scala 27:72]
  wire [1:0] _T_21963 = _T_22481 ? bht_bank_rd_data_out_0_6 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22218 = _T_22217 | _T_21963; // @[Mux.scala 27:72]
  wire [1:0] _T_21964 = _T_22483 ? bht_bank_rd_data_out_0_7 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22219 = _T_22218 | _T_21964; // @[Mux.scala 27:72]
  wire [1:0] _T_21965 = _T_22485 ? bht_bank_rd_data_out_0_8 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22220 = _T_22219 | _T_21965; // @[Mux.scala 27:72]
  wire [1:0] _T_21966 = _T_22487 ? bht_bank_rd_data_out_0_9 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22221 = _T_22220 | _T_21966; // @[Mux.scala 27:72]
  wire [1:0] _T_21967 = _T_22489 ? bht_bank_rd_data_out_0_10 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22222 = _T_22221 | _T_21967; // @[Mux.scala 27:72]
  wire [1:0] _T_21968 = _T_22491 ? bht_bank_rd_data_out_0_11 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22223 = _T_22222 | _T_21968; // @[Mux.scala 27:72]
  wire [1:0] _T_21969 = _T_22493 ? bht_bank_rd_data_out_0_12 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22224 = _T_22223 | _T_21969; // @[Mux.scala 27:72]
  wire [1:0] _T_21970 = _T_22495 ? bht_bank_rd_data_out_0_13 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22225 = _T_22224 | _T_21970; // @[Mux.scala 27:72]
  wire [1:0] _T_21971 = _T_22497 ? bht_bank_rd_data_out_0_14 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22226 = _T_22225 | _T_21971; // @[Mux.scala 27:72]
  wire [1:0] _T_21972 = _T_22499 ? bht_bank_rd_data_out_0_15 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22227 = _T_22226 | _T_21972; // @[Mux.scala 27:72]
  wire [1:0] _T_21973 = _T_22501 ? bht_bank_rd_data_out_0_16 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22228 = _T_22227 | _T_21973; // @[Mux.scala 27:72]
  wire [1:0] _T_21974 = _T_22503 ? bht_bank_rd_data_out_0_17 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22229 = _T_22228 | _T_21974; // @[Mux.scala 27:72]
  wire [1:0] _T_21975 = _T_22505 ? bht_bank_rd_data_out_0_18 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22230 = _T_22229 | _T_21975; // @[Mux.scala 27:72]
  wire [1:0] _T_21976 = _T_22507 ? bht_bank_rd_data_out_0_19 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22231 = _T_22230 | _T_21976; // @[Mux.scala 27:72]
  wire [1:0] _T_21977 = _T_22509 ? bht_bank_rd_data_out_0_20 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22232 = _T_22231 | _T_21977; // @[Mux.scala 27:72]
  wire [1:0] _T_21978 = _T_22511 ? bht_bank_rd_data_out_0_21 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22233 = _T_22232 | _T_21978; // @[Mux.scala 27:72]
  wire [1:0] _T_21979 = _T_22513 ? bht_bank_rd_data_out_0_22 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22234 = _T_22233 | _T_21979; // @[Mux.scala 27:72]
  wire [1:0] _T_21980 = _T_22515 ? bht_bank_rd_data_out_0_23 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22235 = _T_22234 | _T_21980; // @[Mux.scala 27:72]
  wire [1:0] _T_21981 = _T_22517 ? bht_bank_rd_data_out_0_24 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22236 = _T_22235 | _T_21981; // @[Mux.scala 27:72]
  wire [1:0] _T_21982 = _T_22519 ? bht_bank_rd_data_out_0_25 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22237 = _T_22236 | _T_21982; // @[Mux.scala 27:72]
  wire [1:0] _T_21983 = _T_22521 ? bht_bank_rd_data_out_0_26 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22238 = _T_22237 | _T_21983; // @[Mux.scala 27:72]
  wire [1:0] _T_21984 = _T_22523 ? bht_bank_rd_data_out_0_27 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22239 = _T_22238 | _T_21984; // @[Mux.scala 27:72]
  wire [1:0] _T_21985 = _T_22525 ? bht_bank_rd_data_out_0_28 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22240 = _T_22239 | _T_21985; // @[Mux.scala 27:72]
  wire [1:0] _T_21986 = _T_22527 ? bht_bank_rd_data_out_0_29 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22241 = _T_22240 | _T_21986; // @[Mux.scala 27:72]
  wire [1:0] _T_21987 = _T_22529 ? bht_bank_rd_data_out_0_30 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22242 = _T_22241 | _T_21987; // @[Mux.scala 27:72]
  wire [1:0] _T_21988 = _T_22531 ? bht_bank_rd_data_out_0_31 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22243 = _T_22242 | _T_21988; // @[Mux.scala 27:72]
  wire [1:0] _T_21989 = _T_22533 ? bht_bank_rd_data_out_0_32 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22244 = _T_22243 | _T_21989; // @[Mux.scala 27:72]
  wire [1:0] _T_21990 = _T_22535 ? bht_bank_rd_data_out_0_33 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22245 = _T_22244 | _T_21990; // @[Mux.scala 27:72]
  wire [1:0] _T_21991 = _T_22537 ? bht_bank_rd_data_out_0_34 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22246 = _T_22245 | _T_21991; // @[Mux.scala 27:72]
  wire [1:0] _T_21992 = _T_22539 ? bht_bank_rd_data_out_0_35 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22247 = _T_22246 | _T_21992; // @[Mux.scala 27:72]
  wire [1:0] _T_21993 = _T_22541 ? bht_bank_rd_data_out_0_36 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22248 = _T_22247 | _T_21993; // @[Mux.scala 27:72]
  wire [1:0] _T_21994 = _T_22543 ? bht_bank_rd_data_out_0_37 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22249 = _T_22248 | _T_21994; // @[Mux.scala 27:72]
  wire [1:0] _T_21995 = _T_22545 ? bht_bank_rd_data_out_0_38 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22250 = _T_22249 | _T_21995; // @[Mux.scala 27:72]
  wire [1:0] _T_21996 = _T_22547 ? bht_bank_rd_data_out_0_39 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22251 = _T_22250 | _T_21996; // @[Mux.scala 27:72]
  wire [1:0] _T_21997 = _T_22549 ? bht_bank_rd_data_out_0_40 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22252 = _T_22251 | _T_21997; // @[Mux.scala 27:72]
  wire [1:0] _T_21998 = _T_22551 ? bht_bank_rd_data_out_0_41 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22253 = _T_22252 | _T_21998; // @[Mux.scala 27:72]
  wire [1:0] _T_21999 = _T_22553 ? bht_bank_rd_data_out_0_42 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22254 = _T_22253 | _T_21999; // @[Mux.scala 27:72]
  wire [1:0] _T_22000 = _T_22555 ? bht_bank_rd_data_out_0_43 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22255 = _T_22254 | _T_22000; // @[Mux.scala 27:72]
  wire [1:0] _T_22001 = _T_22557 ? bht_bank_rd_data_out_0_44 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22256 = _T_22255 | _T_22001; // @[Mux.scala 27:72]
  wire [1:0] _T_22002 = _T_22559 ? bht_bank_rd_data_out_0_45 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22257 = _T_22256 | _T_22002; // @[Mux.scala 27:72]
  wire [1:0] _T_22003 = _T_22561 ? bht_bank_rd_data_out_0_46 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22258 = _T_22257 | _T_22003; // @[Mux.scala 27:72]
  wire [1:0] _T_22004 = _T_22563 ? bht_bank_rd_data_out_0_47 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22259 = _T_22258 | _T_22004; // @[Mux.scala 27:72]
  wire [1:0] _T_22005 = _T_22565 ? bht_bank_rd_data_out_0_48 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22260 = _T_22259 | _T_22005; // @[Mux.scala 27:72]
  wire [1:0] _T_22006 = _T_22567 ? bht_bank_rd_data_out_0_49 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22261 = _T_22260 | _T_22006; // @[Mux.scala 27:72]
  wire [1:0] _T_22007 = _T_22569 ? bht_bank_rd_data_out_0_50 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22262 = _T_22261 | _T_22007; // @[Mux.scala 27:72]
  wire [1:0] _T_22008 = _T_22571 ? bht_bank_rd_data_out_0_51 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22263 = _T_22262 | _T_22008; // @[Mux.scala 27:72]
  wire [1:0] _T_22009 = _T_22573 ? bht_bank_rd_data_out_0_52 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22264 = _T_22263 | _T_22009; // @[Mux.scala 27:72]
  wire [1:0] _T_22010 = _T_22575 ? bht_bank_rd_data_out_0_53 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22265 = _T_22264 | _T_22010; // @[Mux.scala 27:72]
  wire [1:0] _T_22011 = _T_22577 ? bht_bank_rd_data_out_0_54 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22266 = _T_22265 | _T_22011; // @[Mux.scala 27:72]
  wire [1:0] _T_22012 = _T_22579 ? bht_bank_rd_data_out_0_55 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22267 = _T_22266 | _T_22012; // @[Mux.scala 27:72]
  wire [1:0] _T_22013 = _T_22581 ? bht_bank_rd_data_out_0_56 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22268 = _T_22267 | _T_22013; // @[Mux.scala 27:72]
  wire [1:0] _T_22014 = _T_22583 ? bht_bank_rd_data_out_0_57 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22269 = _T_22268 | _T_22014; // @[Mux.scala 27:72]
  wire [1:0] _T_22015 = _T_22585 ? bht_bank_rd_data_out_0_58 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22270 = _T_22269 | _T_22015; // @[Mux.scala 27:72]
  wire [1:0] _T_22016 = _T_22587 ? bht_bank_rd_data_out_0_59 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22271 = _T_22270 | _T_22016; // @[Mux.scala 27:72]
  wire [1:0] _T_22017 = _T_22589 ? bht_bank_rd_data_out_0_60 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22272 = _T_22271 | _T_22017; // @[Mux.scala 27:72]
  wire [1:0] _T_22018 = _T_22591 ? bht_bank_rd_data_out_0_61 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22273 = _T_22272 | _T_22018; // @[Mux.scala 27:72]
  wire [1:0] _T_22019 = _T_22593 ? bht_bank_rd_data_out_0_62 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22274 = _T_22273 | _T_22019; // @[Mux.scala 27:72]
  wire [1:0] _T_22020 = _T_22595 ? bht_bank_rd_data_out_0_63 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22275 = _T_22274 | _T_22020; // @[Mux.scala 27:72]
  wire [1:0] _T_22021 = _T_22597 ? bht_bank_rd_data_out_0_64 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22276 = _T_22275 | _T_22021; // @[Mux.scala 27:72]
  wire [1:0] _T_22022 = _T_22599 ? bht_bank_rd_data_out_0_65 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22277 = _T_22276 | _T_22022; // @[Mux.scala 27:72]
  wire [1:0] _T_22023 = _T_22601 ? bht_bank_rd_data_out_0_66 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22278 = _T_22277 | _T_22023; // @[Mux.scala 27:72]
  wire [1:0] _T_22024 = _T_22603 ? bht_bank_rd_data_out_0_67 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22279 = _T_22278 | _T_22024; // @[Mux.scala 27:72]
  wire [1:0] _T_22025 = _T_22605 ? bht_bank_rd_data_out_0_68 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22280 = _T_22279 | _T_22025; // @[Mux.scala 27:72]
  wire [1:0] _T_22026 = _T_22607 ? bht_bank_rd_data_out_0_69 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22281 = _T_22280 | _T_22026; // @[Mux.scala 27:72]
  wire [1:0] _T_22027 = _T_22609 ? bht_bank_rd_data_out_0_70 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22282 = _T_22281 | _T_22027; // @[Mux.scala 27:72]
  wire [1:0] _T_22028 = _T_22611 ? bht_bank_rd_data_out_0_71 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22283 = _T_22282 | _T_22028; // @[Mux.scala 27:72]
  wire [1:0] _T_22029 = _T_22613 ? bht_bank_rd_data_out_0_72 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22284 = _T_22283 | _T_22029; // @[Mux.scala 27:72]
  wire [1:0] _T_22030 = _T_22615 ? bht_bank_rd_data_out_0_73 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22285 = _T_22284 | _T_22030; // @[Mux.scala 27:72]
  wire [1:0] _T_22031 = _T_22617 ? bht_bank_rd_data_out_0_74 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22286 = _T_22285 | _T_22031; // @[Mux.scala 27:72]
  wire [1:0] _T_22032 = _T_22619 ? bht_bank_rd_data_out_0_75 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22287 = _T_22286 | _T_22032; // @[Mux.scala 27:72]
  wire [1:0] _T_22033 = _T_22621 ? bht_bank_rd_data_out_0_76 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22288 = _T_22287 | _T_22033; // @[Mux.scala 27:72]
  wire [1:0] _T_22034 = _T_22623 ? bht_bank_rd_data_out_0_77 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22289 = _T_22288 | _T_22034; // @[Mux.scala 27:72]
  wire [1:0] _T_22035 = _T_22625 ? bht_bank_rd_data_out_0_78 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22290 = _T_22289 | _T_22035; // @[Mux.scala 27:72]
  wire [1:0] _T_22036 = _T_22627 ? bht_bank_rd_data_out_0_79 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22291 = _T_22290 | _T_22036; // @[Mux.scala 27:72]
  wire [1:0] _T_22037 = _T_22629 ? bht_bank_rd_data_out_0_80 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22292 = _T_22291 | _T_22037; // @[Mux.scala 27:72]
  wire [1:0] _T_22038 = _T_22631 ? bht_bank_rd_data_out_0_81 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22293 = _T_22292 | _T_22038; // @[Mux.scala 27:72]
  wire [1:0] _T_22039 = _T_22633 ? bht_bank_rd_data_out_0_82 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22294 = _T_22293 | _T_22039; // @[Mux.scala 27:72]
  wire [1:0] _T_22040 = _T_22635 ? bht_bank_rd_data_out_0_83 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22295 = _T_22294 | _T_22040; // @[Mux.scala 27:72]
  wire [1:0] _T_22041 = _T_22637 ? bht_bank_rd_data_out_0_84 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22296 = _T_22295 | _T_22041; // @[Mux.scala 27:72]
  wire [1:0] _T_22042 = _T_22639 ? bht_bank_rd_data_out_0_85 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22297 = _T_22296 | _T_22042; // @[Mux.scala 27:72]
  wire [1:0] _T_22043 = _T_22641 ? bht_bank_rd_data_out_0_86 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22298 = _T_22297 | _T_22043; // @[Mux.scala 27:72]
  wire [1:0] _T_22044 = _T_22643 ? bht_bank_rd_data_out_0_87 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22299 = _T_22298 | _T_22044; // @[Mux.scala 27:72]
  wire [1:0] _T_22045 = _T_22645 ? bht_bank_rd_data_out_0_88 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22300 = _T_22299 | _T_22045; // @[Mux.scala 27:72]
  wire [1:0] _T_22046 = _T_22647 ? bht_bank_rd_data_out_0_89 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22301 = _T_22300 | _T_22046; // @[Mux.scala 27:72]
  wire [1:0] _T_22047 = _T_22649 ? bht_bank_rd_data_out_0_90 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22302 = _T_22301 | _T_22047; // @[Mux.scala 27:72]
  wire [1:0] _T_22048 = _T_22651 ? bht_bank_rd_data_out_0_91 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22303 = _T_22302 | _T_22048; // @[Mux.scala 27:72]
  wire [1:0] _T_22049 = _T_22653 ? bht_bank_rd_data_out_0_92 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22304 = _T_22303 | _T_22049; // @[Mux.scala 27:72]
  wire [1:0] _T_22050 = _T_22655 ? bht_bank_rd_data_out_0_93 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22305 = _T_22304 | _T_22050; // @[Mux.scala 27:72]
  wire [1:0] _T_22051 = _T_22657 ? bht_bank_rd_data_out_0_94 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22306 = _T_22305 | _T_22051; // @[Mux.scala 27:72]
  wire [1:0] _T_22052 = _T_22659 ? bht_bank_rd_data_out_0_95 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22307 = _T_22306 | _T_22052; // @[Mux.scala 27:72]
  wire [1:0] _T_22053 = _T_22661 ? bht_bank_rd_data_out_0_96 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22308 = _T_22307 | _T_22053; // @[Mux.scala 27:72]
  wire [1:0] _T_22054 = _T_22663 ? bht_bank_rd_data_out_0_97 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22309 = _T_22308 | _T_22054; // @[Mux.scala 27:72]
  wire [1:0] _T_22055 = _T_22665 ? bht_bank_rd_data_out_0_98 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22310 = _T_22309 | _T_22055; // @[Mux.scala 27:72]
  wire [1:0] _T_22056 = _T_22667 ? bht_bank_rd_data_out_0_99 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22311 = _T_22310 | _T_22056; // @[Mux.scala 27:72]
  wire [1:0] _T_22057 = _T_22669 ? bht_bank_rd_data_out_0_100 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22312 = _T_22311 | _T_22057; // @[Mux.scala 27:72]
  wire [1:0] _T_22058 = _T_22671 ? bht_bank_rd_data_out_0_101 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22313 = _T_22312 | _T_22058; // @[Mux.scala 27:72]
  wire [1:0] _T_22059 = _T_22673 ? bht_bank_rd_data_out_0_102 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22314 = _T_22313 | _T_22059; // @[Mux.scala 27:72]
  wire [1:0] _T_22060 = _T_22675 ? bht_bank_rd_data_out_0_103 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22315 = _T_22314 | _T_22060; // @[Mux.scala 27:72]
  wire [1:0] _T_22061 = _T_22677 ? bht_bank_rd_data_out_0_104 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22316 = _T_22315 | _T_22061; // @[Mux.scala 27:72]
  wire [1:0] _T_22062 = _T_22679 ? bht_bank_rd_data_out_0_105 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22317 = _T_22316 | _T_22062; // @[Mux.scala 27:72]
  wire [1:0] _T_22063 = _T_22681 ? bht_bank_rd_data_out_0_106 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22318 = _T_22317 | _T_22063; // @[Mux.scala 27:72]
  wire [1:0] _T_22064 = _T_22683 ? bht_bank_rd_data_out_0_107 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22319 = _T_22318 | _T_22064; // @[Mux.scala 27:72]
  wire [1:0] _T_22065 = _T_22685 ? bht_bank_rd_data_out_0_108 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22320 = _T_22319 | _T_22065; // @[Mux.scala 27:72]
  wire [1:0] _T_22066 = _T_22687 ? bht_bank_rd_data_out_0_109 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22321 = _T_22320 | _T_22066; // @[Mux.scala 27:72]
  wire [1:0] _T_22067 = _T_22689 ? bht_bank_rd_data_out_0_110 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22322 = _T_22321 | _T_22067; // @[Mux.scala 27:72]
  wire [1:0] _T_22068 = _T_22691 ? bht_bank_rd_data_out_0_111 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22323 = _T_22322 | _T_22068; // @[Mux.scala 27:72]
  wire [1:0] _T_22069 = _T_22693 ? bht_bank_rd_data_out_0_112 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22324 = _T_22323 | _T_22069; // @[Mux.scala 27:72]
  wire [1:0] _T_22070 = _T_22695 ? bht_bank_rd_data_out_0_113 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22325 = _T_22324 | _T_22070; // @[Mux.scala 27:72]
  wire [1:0] _T_22071 = _T_22697 ? bht_bank_rd_data_out_0_114 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22326 = _T_22325 | _T_22071; // @[Mux.scala 27:72]
  wire [1:0] _T_22072 = _T_22699 ? bht_bank_rd_data_out_0_115 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22327 = _T_22326 | _T_22072; // @[Mux.scala 27:72]
  wire [1:0] _T_22073 = _T_22701 ? bht_bank_rd_data_out_0_116 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22328 = _T_22327 | _T_22073; // @[Mux.scala 27:72]
  wire [1:0] _T_22074 = _T_22703 ? bht_bank_rd_data_out_0_117 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22329 = _T_22328 | _T_22074; // @[Mux.scala 27:72]
  wire [1:0] _T_22075 = _T_22705 ? bht_bank_rd_data_out_0_118 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22330 = _T_22329 | _T_22075; // @[Mux.scala 27:72]
  wire [1:0] _T_22076 = _T_22707 ? bht_bank_rd_data_out_0_119 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22331 = _T_22330 | _T_22076; // @[Mux.scala 27:72]
  wire [1:0] _T_22077 = _T_22709 ? bht_bank_rd_data_out_0_120 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22332 = _T_22331 | _T_22077; // @[Mux.scala 27:72]
  wire [1:0] _T_22078 = _T_22711 ? bht_bank_rd_data_out_0_121 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22333 = _T_22332 | _T_22078; // @[Mux.scala 27:72]
  wire [1:0] _T_22079 = _T_22713 ? bht_bank_rd_data_out_0_122 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22334 = _T_22333 | _T_22079; // @[Mux.scala 27:72]
  wire [1:0] _T_22080 = _T_22715 ? bht_bank_rd_data_out_0_123 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22335 = _T_22334 | _T_22080; // @[Mux.scala 27:72]
  wire [1:0] _T_22081 = _T_22717 ? bht_bank_rd_data_out_0_124 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22336 = _T_22335 | _T_22081; // @[Mux.scala 27:72]
  wire [1:0] _T_22082 = _T_22719 ? bht_bank_rd_data_out_0_125 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22337 = _T_22336 | _T_22082; // @[Mux.scala 27:72]
  wire [1:0] _T_22083 = _T_22721 ? bht_bank_rd_data_out_0_126 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22338 = _T_22337 | _T_22083; // @[Mux.scala 27:72]
  wire [1:0] _T_22084 = _T_22723 ? bht_bank_rd_data_out_0_127 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22339 = _T_22338 | _T_22084; // @[Mux.scala 27:72]
  wire [1:0] _T_22085 = _T_22725 ? bht_bank_rd_data_out_0_128 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22340 = _T_22339 | _T_22085; // @[Mux.scala 27:72]
  wire [1:0] _T_22086 = _T_22727 ? bht_bank_rd_data_out_0_129 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22341 = _T_22340 | _T_22086; // @[Mux.scala 27:72]
  wire [1:0] _T_22087 = _T_22729 ? bht_bank_rd_data_out_0_130 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22342 = _T_22341 | _T_22087; // @[Mux.scala 27:72]
  wire [1:0] _T_22088 = _T_22731 ? bht_bank_rd_data_out_0_131 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22343 = _T_22342 | _T_22088; // @[Mux.scala 27:72]
  wire [1:0] _T_22089 = _T_22733 ? bht_bank_rd_data_out_0_132 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22344 = _T_22343 | _T_22089; // @[Mux.scala 27:72]
  wire [1:0] _T_22090 = _T_22735 ? bht_bank_rd_data_out_0_133 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22345 = _T_22344 | _T_22090; // @[Mux.scala 27:72]
  wire [1:0] _T_22091 = _T_22737 ? bht_bank_rd_data_out_0_134 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22346 = _T_22345 | _T_22091; // @[Mux.scala 27:72]
  wire [1:0] _T_22092 = _T_22739 ? bht_bank_rd_data_out_0_135 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22347 = _T_22346 | _T_22092; // @[Mux.scala 27:72]
  wire [1:0] _T_22093 = _T_22741 ? bht_bank_rd_data_out_0_136 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22348 = _T_22347 | _T_22093; // @[Mux.scala 27:72]
  wire [1:0] _T_22094 = _T_22743 ? bht_bank_rd_data_out_0_137 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22349 = _T_22348 | _T_22094; // @[Mux.scala 27:72]
  wire [1:0] _T_22095 = _T_22745 ? bht_bank_rd_data_out_0_138 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22350 = _T_22349 | _T_22095; // @[Mux.scala 27:72]
  wire [1:0] _T_22096 = _T_22747 ? bht_bank_rd_data_out_0_139 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22351 = _T_22350 | _T_22096; // @[Mux.scala 27:72]
  wire [1:0] _T_22097 = _T_22749 ? bht_bank_rd_data_out_0_140 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22352 = _T_22351 | _T_22097; // @[Mux.scala 27:72]
  wire [1:0] _T_22098 = _T_22751 ? bht_bank_rd_data_out_0_141 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22353 = _T_22352 | _T_22098; // @[Mux.scala 27:72]
  wire [1:0] _T_22099 = _T_22753 ? bht_bank_rd_data_out_0_142 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22354 = _T_22353 | _T_22099; // @[Mux.scala 27:72]
  wire [1:0] _T_22100 = _T_22755 ? bht_bank_rd_data_out_0_143 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22355 = _T_22354 | _T_22100; // @[Mux.scala 27:72]
  wire [1:0] _T_22101 = _T_22757 ? bht_bank_rd_data_out_0_144 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22356 = _T_22355 | _T_22101; // @[Mux.scala 27:72]
  wire [1:0] _T_22102 = _T_22759 ? bht_bank_rd_data_out_0_145 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22357 = _T_22356 | _T_22102; // @[Mux.scala 27:72]
  wire [1:0] _T_22103 = _T_22761 ? bht_bank_rd_data_out_0_146 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22358 = _T_22357 | _T_22103; // @[Mux.scala 27:72]
  wire [1:0] _T_22104 = _T_22763 ? bht_bank_rd_data_out_0_147 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22359 = _T_22358 | _T_22104; // @[Mux.scala 27:72]
  wire [1:0] _T_22105 = _T_22765 ? bht_bank_rd_data_out_0_148 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22360 = _T_22359 | _T_22105; // @[Mux.scala 27:72]
  wire [1:0] _T_22106 = _T_22767 ? bht_bank_rd_data_out_0_149 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22361 = _T_22360 | _T_22106; // @[Mux.scala 27:72]
  wire [1:0] _T_22107 = _T_22769 ? bht_bank_rd_data_out_0_150 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22362 = _T_22361 | _T_22107; // @[Mux.scala 27:72]
  wire [1:0] _T_22108 = _T_22771 ? bht_bank_rd_data_out_0_151 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22363 = _T_22362 | _T_22108; // @[Mux.scala 27:72]
  wire [1:0] _T_22109 = _T_22773 ? bht_bank_rd_data_out_0_152 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22364 = _T_22363 | _T_22109; // @[Mux.scala 27:72]
  wire [1:0] _T_22110 = _T_22775 ? bht_bank_rd_data_out_0_153 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22365 = _T_22364 | _T_22110; // @[Mux.scala 27:72]
  wire [1:0] _T_22111 = _T_22777 ? bht_bank_rd_data_out_0_154 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22366 = _T_22365 | _T_22111; // @[Mux.scala 27:72]
  wire [1:0] _T_22112 = _T_22779 ? bht_bank_rd_data_out_0_155 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22367 = _T_22366 | _T_22112; // @[Mux.scala 27:72]
  wire [1:0] _T_22113 = _T_22781 ? bht_bank_rd_data_out_0_156 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22368 = _T_22367 | _T_22113; // @[Mux.scala 27:72]
  wire [1:0] _T_22114 = _T_22783 ? bht_bank_rd_data_out_0_157 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22369 = _T_22368 | _T_22114; // @[Mux.scala 27:72]
  wire [1:0] _T_22115 = _T_22785 ? bht_bank_rd_data_out_0_158 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22370 = _T_22369 | _T_22115; // @[Mux.scala 27:72]
  wire [1:0] _T_22116 = _T_22787 ? bht_bank_rd_data_out_0_159 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22371 = _T_22370 | _T_22116; // @[Mux.scala 27:72]
  wire [1:0] _T_22117 = _T_22789 ? bht_bank_rd_data_out_0_160 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22372 = _T_22371 | _T_22117; // @[Mux.scala 27:72]
  wire [1:0] _T_22118 = _T_22791 ? bht_bank_rd_data_out_0_161 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22373 = _T_22372 | _T_22118; // @[Mux.scala 27:72]
  wire [1:0] _T_22119 = _T_22793 ? bht_bank_rd_data_out_0_162 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22374 = _T_22373 | _T_22119; // @[Mux.scala 27:72]
  wire [1:0] _T_22120 = _T_22795 ? bht_bank_rd_data_out_0_163 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22375 = _T_22374 | _T_22120; // @[Mux.scala 27:72]
  wire [1:0] _T_22121 = _T_22797 ? bht_bank_rd_data_out_0_164 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22376 = _T_22375 | _T_22121; // @[Mux.scala 27:72]
  wire [1:0] _T_22122 = _T_22799 ? bht_bank_rd_data_out_0_165 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22377 = _T_22376 | _T_22122; // @[Mux.scala 27:72]
  wire [1:0] _T_22123 = _T_22801 ? bht_bank_rd_data_out_0_166 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22378 = _T_22377 | _T_22123; // @[Mux.scala 27:72]
  wire [1:0] _T_22124 = _T_22803 ? bht_bank_rd_data_out_0_167 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22379 = _T_22378 | _T_22124; // @[Mux.scala 27:72]
  wire [1:0] _T_22125 = _T_22805 ? bht_bank_rd_data_out_0_168 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22380 = _T_22379 | _T_22125; // @[Mux.scala 27:72]
  wire [1:0] _T_22126 = _T_22807 ? bht_bank_rd_data_out_0_169 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22381 = _T_22380 | _T_22126; // @[Mux.scala 27:72]
  wire [1:0] _T_22127 = _T_22809 ? bht_bank_rd_data_out_0_170 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22382 = _T_22381 | _T_22127; // @[Mux.scala 27:72]
  wire [1:0] _T_22128 = _T_22811 ? bht_bank_rd_data_out_0_171 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22383 = _T_22382 | _T_22128; // @[Mux.scala 27:72]
  wire [1:0] _T_22129 = _T_22813 ? bht_bank_rd_data_out_0_172 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22384 = _T_22383 | _T_22129; // @[Mux.scala 27:72]
  wire [1:0] _T_22130 = _T_22815 ? bht_bank_rd_data_out_0_173 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22385 = _T_22384 | _T_22130; // @[Mux.scala 27:72]
  wire [1:0] _T_22131 = _T_22817 ? bht_bank_rd_data_out_0_174 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22386 = _T_22385 | _T_22131; // @[Mux.scala 27:72]
  wire [1:0] _T_22132 = _T_22819 ? bht_bank_rd_data_out_0_175 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22387 = _T_22386 | _T_22132; // @[Mux.scala 27:72]
  wire [1:0] _T_22133 = _T_22821 ? bht_bank_rd_data_out_0_176 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22388 = _T_22387 | _T_22133; // @[Mux.scala 27:72]
  wire [1:0] _T_22134 = _T_22823 ? bht_bank_rd_data_out_0_177 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22389 = _T_22388 | _T_22134; // @[Mux.scala 27:72]
  wire [1:0] _T_22135 = _T_22825 ? bht_bank_rd_data_out_0_178 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22390 = _T_22389 | _T_22135; // @[Mux.scala 27:72]
  wire [1:0] _T_22136 = _T_22827 ? bht_bank_rd_data_out_0_179 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22391 = _T_22390 | _T_22136; // @[Mux.scala 27:72]
  wire [1:0] _T_22137 = _T_22829 ? bht_bank_rd_data_out_0_180 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22392 = _T_22391 | _T_22137; // @[Mux.scala 27:72]
  wire [1:0] _T_22138 = _T_22831 ? bht_bank_rd_data_out_0_181 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22393 = _T_22392 | _T_22138; // @[Mux.scala 27:72]
  wire [1:0] _T_22139 = _T_22833 ? bht_bank_rd_data_out_0_182 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22394 = _T_22393 | _T_22139; // @[Mux.scala 27:72]
  wire [1:0] _T_22140 = _T_22835 ? bht_bank_rd_data_out_0_183 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22395 = _T_22394 | _T_22140; // @[Mux.scala 27:72]
  wire [1:0] _T_22141 = _T_22837 ? bht_bank_rd_data_out_0_184 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22396 = _T_22395 | _T_22141; // @[Mux.scala 27:72]
  wire [1:0] _T_22142 = _T_22839 ? bht_bank_rd_data_out_0_185 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22397 = _T_22396 | _T_22142; // @[Mux.scala 27:72]
  wire [1:0] _T_22143 = _T_22841 ? bht_bank_rd_data_out_0_186 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22398 = _T_22397 | _T_22143; // @[Mux.scala 27:72]
  wire [1:0] _T_22144 = _T_22843 ? bht_bank_rd_data_out_0_187 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22399 = _T_22398 | _T_22144; // @[Mux.scala 27:72]
  wire [1:0] _T_22145 = _T_22845 ? bht_bank_rd_data_out_0_188 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22400 = _T_22399 | _T_22145; // @[Mux.scala 27:72]
  wire [1:0] _T_22146 = _T_22847 ? bht_bank_rd_data_out_0_189 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22401 = _T_22400 | _T_22146; // @[Mux.scala 27:72]
  wire [1:0] _T_22147 = _T_22849 ? bht_bank_rd_data_out_0_190 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22402 = _T_22401 | _T_22147; // @[Mux.scala 27:72]
  wire [1:0] _T_22148 = _T_22851 ? bht_bank_rd_data_out_0_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22403 = _T_22402 | _T_22148; // @[Mux.scala 27:72]
  wire [1:0] _T_22149 = _T_22853 ? bht_bank_rd_data_out_0_192 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22404 = _T_22403 | _T_22149; // @[Mux.scala 27:72]
  wire [1:0] _T_22150 = _T_22855 ? bht_bank_rd_data_out_0_193 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22405 = _T_22404 | _T_22150; // @[Mux.scala 27:72]
  wire [1:0] _T_22151 = _T_22857 ? bht_bank_rd_data_out_0_194 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22406 = _T_22405 | _T_22151; // @[Mux.scala 27:72]
  wire [1:0] _T_22152 = _T_22859 ? bht_bank_rd_data_out_0_195 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22407 = _T_22406 | _T_22152; // @[Mux.scala 27:72]
  wire [1:0] _T_22153 = _T_22861 ? bht_bank_rd_data_out_0_196 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22408 = _T_22407 | _T_22153; // @[Mux.scala 27:72]
  wire [1:0] _T_22154 = _T_22863 ? bht_bank_rd_data_out_0_197 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22409 = _T_22408 | _T_22154; // @[Mux.scala 27:72]
  wire [1:0] _T_22155 = _T_22865 ? bht_bank_rd_data_out_0_198 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22410 = _T_22409 | _T_22155; // @[Mux.scala 27:72]
  wire [1:0] _T_22156 = _T_22867 ? bht_bank_rd_data_out_0_199 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22411 = _T_22410 | _T_22156; // @[Mux.scala 27:72]
  wire [1:0] _T_22157 = _T_22869 ? bht_bank_rd_data_out_0_200 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22412 = _T_22411 | _T_22157; // @[Mux.scala 27:72]
  wire [1:0] _T_22158 = _T_22871 ? bht_bank_rd_data_out_0_201 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22413 = _T_22412 | _T_22158; // @[Mux.scala 27:72]
  wire [1:0] _T_22159 = _T_22873 ? bht_bank_rd_data_out_0_202 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22414 = _T_22413 | _T_22159; // @[Mux.scala 27:72]
  wire [1:0] _T_22160 = _T_22875 ? bht_bank_rd_data_out_0_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22415 = _T_22414 | _T_22160; // @[Mux.scala 27:72]
  wire [1:0] _T_22161 = _T_22877 ? bht_bank_rd_data_out_0_204 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22416 = _T_22415 | _T_22161; // @[Mux.scala 27:72]
  wire [1:0] _T_22162 = _T_22879 ? bht_bank_rd_data_out_0_205 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22417 = _T_22416 | _T_22162; // @[Mux.scala 27:72]
  wire [1:0] _T_22163 = _T_22881 ? bht_bank_rd_data_out_0_206 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22418 = _T_22417 | _T_22163; // @[Mux.scala 27:72]
  wire [1:0] _T_22164 = _T_22883 ? bht_bank_rd_data_out_0_207 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22419 = _T_22418 | _T_22164; // @[Mux.scala 27:72]
  wire [1:0] _T_22165 = _T_22885 ? bht_bank_rd_data_out_0_208 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22420 = _T_22419 | _T_22165; // @[Mux.scala 27:72]
  wire [1:0] _T_22166 = _T_22887 ? bht_bank_rd_data_out_0_209 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22421 = _T_22420 | _T_22166; // @[Mux.scala 27:72]
  wire [1:0] _T_22167 = _T_22889 ? bht_bank_rd_data_out_0_210 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22422 = _T_22421 | _T_22167; // @[Mux.scala 27:72]
  wire [1:0] _T_22168 = _T_22891 ? bht_bank_rd_data_out_0_211 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22423 = _T_22422 | _T_22168; // @[Mux.scala 27:72]
  wire [1:0] _T_22169 = _T_22893 ? bht_bank_rd_data_out_0_212 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22424 = _T_22423 | _T_22169; // @[Mux.scala 27:72]
  wire [1:0] _T_22170 = _T_22895 ? bht_bank_rd_data_out_0_213 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22425 = _T_22424 | _T_22170; // @[Mux.scala 27:72]
  wire [1:0] _T_22171 = _T_22897 ? bht_bank_rd_data_out_0_214 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22426 = _T_22425 | _T_22171; // @[Mux.scala 27:72]
  wire [1:0] _T_22172 = _T_22899 ? bht_bank_rd_data_out_0_215 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22427 = _T_22426 | _T_22172; // @[Mux.scala 27:72]
  wire [1:0] _T_22173 = _T_22901 ? bht_bank_rd_data_out_0_216 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22428 = _T_22427 | _T_22173; // @[Mux.scala 27:72]
  wire [1:0] _T_22174 = _T_22903 ? bht_bank_rd_data_out_0_217 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22429 = _T_22428 | _T_22174; // @[Mux.scala 27:72]
  wire [1:0] _T_22175 = _T_22905 ? bht_bank_rd_data_out_0_218 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22430 = _T_22429 | _T_22175; // @[Mux.scala 27:72]
  wire [1:0] _T_22176 = _T_22907 ? bht_bank_rd_data_out_0_219 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22431 = _T_22430 | _T_22176; // @[Mux.scala 27:72]
  wire [1:0] _T_22177 = _T_22909 ? bht_bank_rd_data_out_0_220 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22432 = _T_22431 | _T_22177; // @[Mux.scala 27:72]
  wire [1:0] _T_22178 = _T_22911 ? bht_bank_rd_data_out_0_221 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22433 = _T_22432 | _T_22178; // @[Mux.scala 27:72]
  wire [1:0] _T_22179 = _T_22913 ? bht_bank_rd_data_out_0_222 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22434 = _T_22433 | _T_22179; // @[Mux.scala 27:72]
  wire [1:0] _T_22180 = _T_22915 ? bht_bank_rd_data_out_0_223 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22435 = _T_22434 | _T_22180; // @[Mux.scala 27:72]
  wire [1:0] _T_22181 = _T_22917 ? bht_bank_rd_data_out_0_224 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22436 = _T_22435 | _T_22181; // @[Mux.scala 27:72]
  wire [1:0] _T_22182 = _T_22919 ? bht_bank_rd_data_out_0_225 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22437 = _T_22436 | _T_22182; // @[Mux.scala 27:72]
  wire [1:0] _T_22183 = _T_22921 ? bht_bank_rd_data_out_0_226 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22438 = _T_22437 | _T_22183; // @[Mux.scala 27:72]
  wire [1:0] _T_22184 = _T_22923 ? bht_bank_rd_data_out_0_227 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22439 = _T_22438 | _T_22184; // @[Mux.scala 27:72]
  wire [1:0] _T_22185 = _T_22925 ? bht_bank_rd_data_out_0_228 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22440 = _T_22439 | _T_22185; // @[Mux.scala 27:72]
  wire [1:0] _T_22186 = _T_22927 ? bht_bank_rd_data_out_0_229 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22441 = _T_22440 | _T_22186; // @[Mux.scala 27:72]
  wire [1:0] _T_22187 = _T_22929 ? bht_bank_rd_data_out_0_230 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22442 = _T_22441 | _T_22187; // @[Mux.scala 27:72]
  wire [1:0] _T_22188 = _T_22931 ? bht_bank_rd_data_out_0_231 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22443 = _T_22442 | _T_22188; // @[Mux.scala 27:72]
  wire [1:0] _T_22189 = _T_22933 ? bht_bank_rd_data_out_0_232 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22444 = _T_22443 | _T_22189; // @[Mux.scala 27:72]
  wire [1:0] _T_22190 = _T_22935 ? bht_bank_rd_data_out_0_233 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22445 = _T_22444 | _T_22190; // @[Mux.scala 27:72]
  wire [1:0] _T_22191 = _T_22937 ? bht_bank_rd_data_out_0_234 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22446 = _T_22445 | _T_22191; // @[Mux.scala 27:72]
  wire [1:0] _T_22192 = _T_22939 ? bht_bank_rd_data_out_0_235 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22447 = _T_22446 | _T_22192; // @[Mux.scala 27:72]
  wire [1:0] _T_22193 = _T_22941 ? bht_bank_rd_data_out_0_236 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22448 = _T_22447 | _T_22193; // @[Mux.scala 27:72]
  wire [1:0] _T_22194 = _T_22943 ? bht_bank_rd_data_out_0_237 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22449 = _T_22448 | _T_22194; // @[Mux.scala 27:72]
  wire [1:0] _T_22195 = _T_22945 ? bht_bank_rd_data_out_0_238 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22450 = _T_22449 | _T_22195; // @[Mux.scala 27:72]
  wire [1:0] _T_22196 = _T_22947 ? bht_bank_rd_data_out_0_239 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22451 = _T_22450 | _T_22196; // @[Mux.scala 27:72]
  wire [1:0] _T_22197 = _T_22949 ? bht_bank_rd_data_out_0_240 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22452 = _T_22451 | _T_22197; // @[Mux.scala 27:72]
  wire [1:0] _T_22198 = _T_22951 ? bht_bank_rd_data_out_0_241 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22453 = _T_22452 | _T_22198; // @[Mux.scala 27:72]
  wire [1:0] _T_22199 = _T_22953 ? bht_bank_rd_data_out_0_242 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22454 = _T_22453 | _T_22199; // @[Mux.scala 27:72]
  wire [1:0] _T_22200 = _T_22955 ? bht_bank_rd_data_out_0_243 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22455 = _T_22454 | _T_22200; // @[Mux.scala 27:72]
  wire [1:0] _T_22201 = _T_22957 ? bht_bank_rd_data_out_0_244 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22456 = _T_22455 | _T_22201; // @[Mux.scala 27:72]
  wire [1:0] _T_22202 = _T_22959 ? bht_bank_rd_data_out_0_245 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22457 = _T_22456 | _T_22202; // @[Mux.scala 27:72]
  wire [1:0] _T_22203 = _T_22961 ? bht_bank_rd_data_out_0_246 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22458 = _T_22457 | _T_22203; // @[Mux.scala 27:72]
  wire [1:0] _T_22204 = _T_22963 ? bht_bank_rd_data_out_0_247 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22459 = _T_22458 | _T_22204; // @[Mux.scala 27:72]
  wire [1:0] _T_22205 = _T_22965 ? bht_bank_rd_data_out_0_248 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22460 = _T_22459 | _T_22205; // @[Mux.scala 27:72]
  wire [1:0] _T_22206 = _T_22967 ? bht_bank_rd_data_out_0_249 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22461 = _T_22460 | _T_22206; // @[Mux.scala 27:72]
  wire [1:0] _T_22207 = _T_22969 ? bht_bank_rd_data_out_0_250 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22462 = _T_22461 | _T_22207; // @[Mux.scala 27:72]
  wire [1:0] _T_22208 = _T_22971 ? bht_bank_rd_data_out_0_251 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22463 = _T_22462 | _T_22208; // @[Mux.scala 27:72]
  wire [1:0] _T_22209 = _T_22973 ? bht_bank_rd_data_out_0_252 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22464 = _T_22463 | _T_22209; // @[Mux.scala 27:72]
  wire [1:0] _T_22210 = _T_22975 ? bht_bank_rd_data_out_0_253 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22465 = _T_22464 | _T_22210; // @[Mux.scala 27:72]
  wire [1:0] _T_22211 = _T_22977 ? bht_bank_rd_data_out_0_254 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_22466 = _T_22465 | _T_22211; // @[Mux.scala 27:72]
  wire [1:0] _T_22212 = _T_22979 ? bht_bank_rd_data_out_0_255 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_bank0_rd_data_f = _T_22466 | _T_22212; // @[Mux.scala 27:72]
  wire [1:0] _T_245 = _T_147 ? bht_bank0_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_246 = io_ifc_fetch_addr_f[0] ? bht_bank1_rd_data_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] bht_vbank0_rd_data_f = _T_245 | _T_246; // @[Mux.scala 27:72]
  wire  _T_263 = bht_force_taken_f[0] | bht_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 299:45]
  wire  _T_265 = _T_263 & vwayhit_f[0]; // @[ifu_bp_ctl.scala 299:72]
  wire [1:0] bht_dir_f = {_T_260,_T_265}; // @[Cat.scala 29:58]
  wire  _T_14 = ~bht_dir_f[0]; // @[ifu_bp_ctl.scala 119:23]
  wire [1:0] btb_sel_f = {_T_14,bht_dir_f[0]}; // @[Cat.scala 29:58]
  wire [1:0] fetch_start_f = {io_ifc_fetch_addr_f[0],_T_147}; // @[Cat.scala 29:58]
  wire  _T_36 = io_exu_bp_exu_mp_btag == fetch_rd_tag_f; // @[ifu_bp_ctl.scala 140:53]
  wire  _T_37 = _T_36 & exu_mp_valid; // @[ifu_bp_ctl.scala 140:73]
  wire  _T_38 = _T_37 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 140:88]
  wire  _T_39 = io_exu_bp_exu_mp_index == btb_rd_addr_f; // @[ifu_bp_ctl.scala 140:124]
  wire  fetch_mp_collision_f = _T_38 & _T_39; // @[ifu_bp_ctl.scala 140:109]
  wire  _T_40 = io_exu_bp_exu_mp_btag == fetch_rd_tag_p1_f; // @[ifu_bp_ctl.scala 141:56]
  wire  _T_41 = _T_40 & exu_mp_valid; // @[ifu_bp_ctl.scala 141:79]
  wire  _T_42 = _T_41 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 141:94]
  wire  _T_43 = io_exu_bp_exu_mp_index == btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 141:130]
  wire  fetch_mp_collision_p1_f = _T_42 & _T_43; // @[ifu_bp_ctl.scala 141:115]
  wire [1:0] _T_153 = ~vwayhit_f; // @[ifu_bp_ctl.scala 194:44]
  reg  exu_mp_way_f; // @[Reg.scala 27:20]
  wire [255:0] fetch_wrindex_dec = 256'h1 << btb_rd_addr_f; // @[ifu_bp_ctl.scala 213:31]
  reg [255:0] btb_lru_b0_f; // @[Reg.scala 27:20]
  wire [255:0] _T_181 = fetch_wrindex_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 239:78]
  wire  _T_182 = |_T_181; // @[ifu_bp_ctl.scala 239:94]
  wire  btb_lru_rd_f = fetch_mp_collision_f ? exu_mp_way_f : _T_182; // @[ifu_bp_ctl.scala 239:25]
  wire [1:0] _T_188 = {btb_lru_rd_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_192 = _T_147 ? _T_188 : 2'h0; // @[Mux.scala 27:72]
  wire [255:0] fetch_wrindex_p1_dec = 256'h1 << btb_rd_addr_p1_f; // @[ifu_bp_ctl.scala 216:34]
  wire [255:0] _T_184 = fetch_wrindex_p1_dec & btb_lru_b0_f; // @[ifu_bp_ctl.scala 241:87]
  wire  _T_185 = |_T_184; // @[ifu_bp_ctl.scala 241:103]
  wire  btb_lru_rd_p1_f = fetch_mp_collision_p1_f ? exu_mp_way_f : _T_185; // @[ifu_bp_ctl.scala 241:28]
  wire [1:0] _T_191 = {btb_lru_rd_p1_f,btb_lru_rd_f}; // @[Cat.scala 29:58]
  wire [1:0] _T_193 = io_ifc_fetch_addr_f[0] ? _T_191 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] btb_vlru_rd_f = _T_192 | _T_193; // @[Mux.scala 27:72]
  wire [1:0] _T_154 = _T_153 & btb_vlru_rd_f; // @[ifu_bp_ctl.scala 194:55]
  wire [1:0] _T_204 = _T_147 ? tag_match_way1_expanded_f : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_203 = {tag_match_way1_expanded_p1_f[0],tag_match_way1_expanded_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] _T_205 = io_ifc_fetch_addr_f[0] ? _T_203 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] tag_match_vway1_expanded_f = _T_204 | _T_205; // @[Mux.scala 27:72]
  wire [255:0] mp_wrindex_dec = 256'h1 << io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 210:28]
  wire [255:0] _T_157 = exu_mp_valid ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] mp_wrlru_b0 = mp_wrindex_dec & _T_157; // @[ifu_bp_ctl.scala 219:36]
  wire  _T_160 = vwayhit_f[0] | vwayhit_f[1]; // @[ifu_bp_ctl.scala 222:42]
  wire  _T_161 = _T_160 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 222:58]
  wire  lru_update_valid_f = _T_161 & _T; // @[ifu_bp_ctl.scala 222:79]
  wire [255:0] _T_164 = lru_update_valid_f ? 256'hffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffffff : 256'h0; // @[Bitwise.scala 72:12]
  wire [255:0] fetch_wrlru_b0 = fetch_wrindex_dec & _T_164; // @[ifu_bp_ctl.scala 224:42]
  wire [255:0] fetch_wrlru_p1_b0 = fetch_wrindex_p1_dec & _T_164; // @[ifu_bp_ctl.scala 225:48]
  wire [255:0] _T_167 = ~mp_wrlru_b0; // @[ifu_bp_ctl.scala 227:25]
  wire [255:0] _T_168 = ~fetch_wrlru_b0; // @[ifu_bp_ctl.scala 227:40]
  wire [255:0] btb_lru_b0_hold = _T_167 & _T_168; // @[ifu_bp_ctl.scala 227:38]
  wire  _T_170 = ~io_exu_bp_exu_mp_pkt_bits_way; // @[ifu_bp_ctl.scala 234:39]
  wire [255:0] _T_173 = _T_170 ? mp_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_174 = tag_match_way0_f ? fetch_wrlru_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_175 = tag_match_way0_p1_f ? fetch_wrlru_p1_b0 : 256'h0; // @[Mux.scala 27:72]
  wire [255:0] _T_176 = _T_173 | _T_174; // @[Mux.scala 27:72]
  wire [255:0] _T_177 = _T_176 | _T_175; // @[Mux.scala 27:72]
  wire [255:0] _T_179 = btb_lru_b0_hold & btb_lru_b0_f; // @[ifu_bp_ctl.scala 236:73]
  wire [255:0] btb_lru_b0_ns = _T_177 | _T_179; // @[ifu_bp_ctl.scala 236:55]
  wire  _T_208 = io_ifc_fetch_req_f | exu_mp_valid; // @[ifu_bp_ctl.scala 251:60]
  wire [15:0] _T_223 = btb_sel_f[1] ? btb_vbank1_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_224 = btb_sel_f[0] ? btb_vbank0_rd_data_f[16:1] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] btb_sel_data_f = _T_223 | _T_224; // @[Mux.scala 27:72]
  wire [11:0] btb_rd_tgt_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 267:36]
  wire  btb_rd_pc4_f = btb_sel_data_f[3]; // @[ifu_bp_ctl.scala 268:36]
  wire  btb_rd_call_f = btb_sel_data_f[1]; // @[ifu_bp_ctl.scala 269:37]
  wire  btb_rd_ret_f = btb_sel_data_f[0]; // @[ifu_bp_ctl.scala 270:36]
  wire [1:0] _T_273 = {bht_vbank1_rd_data_f[1],bht_vbank0_rd_data_f[1]}; // @[Cat.scala 29:58]
  wire [1:0] hist1_raw = bht_force_taken_f | _T_273; // @[ifu_bp_ctl.scala 305:34]
  wire [1:0] _T_227 = vwayhit_f & hist1_raw; // @[ifu_bp_ctl.scala 277:39]
  wire  _T_228 = |_T_227; // @[ifu_bp_ctl.scala 277:52]
  wire  _T_229 = _T_228 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 277:56]
  wire  _T_230 = ~leak_one_f_d1; // @[ifu_bp_ctl.scala 277:79]
  wire  _T_231 = _T_229 & _T_230; // @[ifu_bp_ctl.scala 277:77]
  wire  _T_232 = ~io_dec_bp_dec_tlu_bpred_disable; // @[ifu_bp_ctl.scala 277:96]
  wire  _T_268 = io_ifu_bp_hit_taken_f & btb_sel_f[1]; // @[ifu_bp_ctl.scala 302:51]
  wire  _T_269 = ~io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 302:69]
  wire  _T_279 = vwayhit_f[1] & btb_vbank1_rd_data_f[4]; // @[ifu_bp_ctl.scala 311:34]
  wire  _T_282 = vwayhit_f[0] & btb_vbank0_rd_data_f[4]; // @[ifu_bp_ctl.scala 312:34]
  wire  _T_285 = ~btb_vbank1_rd_data_f[2]; // @[ifu_bp_ctl.scala 315:37]
  wire  _T_286 = vwayhit_f[1] & _T_285; // @[ifu_bp_ctl.scala 315:35]
  wire  _T_288 = _T_286 & btb_vbank1_rd_data_f[1]; // @[ifu_bp_ctl.scala 315:65]
  wire  _T_291 = ~btb_vbank0_rd_data_f[2]; // @[ifu_bp_ctl.scala 316:37]
  wire  _T_292 = vwayhit_f[0] & _T_291; // @[ifu_bp_ctl.scala 316:35]
  wire  _T_294 = _T_292 & btb_vbank0_rd_data_f[1]; // @[ifu_bp_ctl.scala 316:65]
  wire [1:0] num_valids = vwayhit_f[1] + vwayhit_f[0]; // @[ifu_bp_ctl.scala 319:35]
  wire [1:0] _T_297 = btb_sel_f & bht_dir_f; // @[ifu_bp_ctl.scala 322:28]
  wire  final_h = |_T_297; // @[ifu_bp_ctl.scala 322:41]
  wire  _T_298 = num_valids == 2'h2; // @[ifu_bp_ctl.scala 326:41]
  wire [7:0] _T_302 = {fghr[5:0],1'h0,final_h}; // @[Cat.scala 29:58]
  wire  _T_303 = num_valids == 2'h1; // @[ifu_bp_ctl.scala 327:41]
  wire [7:0] _T_306 = {fghr[6:0],final_h}; // @[Cat.scala 29:58]
  wire  _T_307 = num_valids == 2'h0; // @[ifu_bp_ctl.scala 328:41]
  wire [7:0] _T_310 = _T_298 ? _T_302 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_311 = _T_303 ? _T_306 : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_312 = _T_307 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_313 = _T_310 | _T_311; // @[Mux.scala 27:72]
  wire [7:0] merged_ghr = _T_313 | _T_312; // @[Mux.scala 27:72]
  reg  exu_flush_final_d1; // @[Reg.scala 27:20]
  wire  _T_316 = ~exu_flush_final_d1; // @[ifu_bp_ctl.scala 337:27]
  wire  _T_317 = _T_316 & io_ifc_fetch_req_f; // @[ifu_bp_ctl.scala 337:47]
  wire  _T_318 = _T_317 & io_ic_hit_f; // @[ifu_bp_ctl.scala 337:70]
  wire  _T_320 = _T_318 & _T_230; // @[ifu_bp_ctl.scala 337:84]
  wire  _T_323 = io_ifc_fetch_req_f & io_ic_hit_f; // @[ifu_bp_ctl.scala 338:70]
  wire  _T_325 = _T_323 & _T_230; // @[ifu_bp_ctl.scala 338:84]
  wire  _T_326 = ~_T_325; // @[ifu_bp_ctl.scala 338:49]
  wire  _T_327 = _T_316 & _T_326; // @[ifu_bp_ctl.scala 338:47]
  wire [7:0] _T_329 = exu_flush_final_d1 ? io_exu_bp_exu_mp_fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_330 = _T_320 ? merged_ghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_331 = _T_327 ? fghr : 8'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_332 = _T_329 | _T_330; // @[Mux.scala 27:72]
  wire [7:0] fghr_ns = _T_332 | _T_331; // @[Mux.scala 27:72]
  wire  _T_336 = leak_one_f ^ leak_one_f_d1; // @[lib.scala 453:21]
  wire  _T_337 = |_T_336; // @[lib.scala 453:29]
  wire  _T_340 = io_exu_bp_exu_mp_pkt_bits_way ^ exu_mp_way_f; // @[lib.scala 453:21]
  wire  _T_341 = |_T_340; // @[lib.scala 453:29]
  wire  _T_344 = io_exu_flush_final ^ exu_flush_final_d1; // @[lib.scala 475:21]
  wire  _T_345 = |_T_344; // @[lib.scala 475:29]
  wire [7:0] _T_348 = fghr_ns ^ fghr; // @[lib.scala 453:21]
  wire  _T_349 = |_T_348; // @[lib.scala 453:29]
  wire [1:0] _T_352 = io_dec_bp_dec_tlu_bpred_disable ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_353 = ~_T_352; // @[ifu_bp_ctl.scala 350:36]
  wire  _T_357 = ~fetch_start_f[0]; // @[ifu_bp_ctl.scala 354:36]
  wire  _T_358 = bht_dir_f[0] & _T_357; // @[ifu_bp_ctl.scala 354:34]
  wire  _T_362 = _T_14 & fetch_start_f[0]; // @[ifu_bp_ctl.scala 354:72]
  wire  _T_363 = _T_358 | _T_362; // @[ifu_bp_ctl.scala 354:55]
  wire  _T_366 = bht_dir_f[0] & fetch_start_f[0]; // @[ifu_bp_ctl.scala 355:34]
  wire  _T_371 = _T_14 & _T_357; // @[ifu_bp_ctl.scala 355:71]
  wire  _T_372 = _T_366 | _T_371; // @[ifu_bp_ctl.scala 355:54]
  wire [1:0] bloc_f = {_T_363,_T_372}; // @[Cat.scala 29:58]
  wire  _T_376 = _T_14 & io_ifc_fetch_addr_f[0]; // @[ifu_bp_ctl.scala 357:35]
  wire  _T_377 = ~btb_rd_pc4_f; // @[ifu_bp_ctl.scala 357:62]
  wire  use_fa_plus = _T_376 & _T_377; // @[ifu_bp_ctl.scala 357:60]
  wire  _T_380 = fetch_start_f[0] & btb_sel_f[0]; // @[ifu_bp_ctl.scala 359:44]
  wire  btb_fg_crossing_f = _T_380 & btb_rd_pc4_f; // @[ifu_bp_ctl.scala 359:59]
  wire  bp_total_branch_offset_f = bloc_f[1] ^ btb_rd_pc4_f; // @[ifu_bp_ctl.scala 360:43]
  wire  _T_384 = io_ifc_fetch_req_f & _T_269; // @[ifu_bp_ctl.scala 361:117]
  wire  _T_385 = _T_384 & io_ic_hit_f; // @[ifu_bp_ctl.scala 361:142]
  reg [29:0] ifc_fetch_adder_prior; // @[Reg.scala 27:20]
  wire  _T_390 = ~btb_fg_crossing_f; // @[ifu_bp_ctl.scala 366:32]
  wire  _T_391 = ~use_fa_plus; // @[ifu_bp_ctl.scala 366:53]
  wire  _T_392 = _T_390 & _T_391; // @[ifu_bp_ctl.scala 366:51]
  wire [29:0] _T_395 = use_fa_plus ? fetch_addr_p1_f : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_396 = btb_fg_crossing_f ? ifc_fetch_adder_prior : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_397 = _T_392 ? io_ifc_fetch_addr_f[30:1] : 30'h0; // @[Mux.scala 27:72]
  wire [29:0] _T_398 = _T_395 | _T_396; // @[Mux.scala 27:72]
  wire [29:0] adder_pc_in_f = _T_398 | _T_397; // @[Mux.scala 27:72]
  wire [31:0] _T_402 = {adder_pc_in_f,bp_total_branch_offset_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_403 = {btb_rd_tgt_f,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_406 = _T_402[12:1] + _T_403[12:1]; // @[lib.scala 68:31]
  wire [18:0] _T_409 = _T_402[31:13] + 19'h1; // @[lib.scala 69:27]
  wire [18:0] _T_412 = _T_402[31:13] - 19'h1; // @[lib.scala 70:27]
  wire  _T_415 = ~_T_406[12]; // @[lib.scala 72:28]
  wire  _T_416 = _T_403[12] ^ _T_415; // @[lib.scala 72:26]
  wire  _T_419 = ~_T_403[12]; // @[lib.scala 73:20]
  wire  _T_421 = _T_419 & _T_406[12]; // @[lib.scala 73:26]
  wire  _T_425 = _T_403[12] & _T_415; // @[lib.scala 74:26]
  wire [18:0] _T_427 = _T_416 ? _T_402[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_428 = _T_421 ? _T_409 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_429 = _T_425 ? _T_412 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_430 = _T_427 | _T_428; // @[Mux.scala 27:72]
  wire [18:0] _T_431 = _T_430 | _T_429; // @[Mux.scala 27:72]
  wire [31:0] bp_btb_target_adder_f = {_T_431,_T_406[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_435 = ~btb_rd_call_f; // @[ifu_bp_ctl.scala 374:55]
  wire  _T_436 = btb_rd_ret_f & _T_435; // @[ifu_bp_ctl.scala 374:53]
  reg [31:0] rets_out_0; // @[Reg.scala 27:20]
  wire  _T_438 = _T_436 & rets_out_0[0]; // @[ifu_bp_ctl.scala 374:70]
  wire  _T_439 = _T_438 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 374:87]
  wire [30:0] _T_441 = _T_439 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_443 = _T_441 & rets_out_0[31:1]; // @[ifu_bp_ctl.scala 374:113]
  wire  _T_448 = ~_T_438; // @[ifu_bp_ctl.scala 375:15]
  wire  _T_449 = _T_448 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 375:65]
  wire [30:0] _T_451 = _T_449 ? 31'h7fffffff : 31'h0; // @[Bitwise.scala 72:12]
  wire [30:0] _T_453 = _T_451 & bp_btb_target_adder_f[31:1]; // @[ifu_bp_ctl.scala 375:91]
  wire [12:0] _T_461 = {11'h0,_T_377,1'h0}; // @[Cat.scala 29:58]
  wire [12:0] _T_464 = _T_402[12:1] + _T_461[12:1]; // @[lib.scala 68:31]
  wire  _T_473 = ~_T_464[12]; // @[lib.scala 72:28]
  wire  _T_474 = _T_461[12] ^ _T_473; // @[lib.scala 72:26]
  wire  _T_477 = ~_T_461[12]; // @[lib.scala 73:20]
  wire  _T_479 = _T_477 & _T_464[12]; // @[lib.scala 73:26]
  wire  _T_483 = _T_461[12] & _T_473; // @[lib.scala 74:26]
  wire [18:0] _T_485 = _T_474 ? _T_402[31:13] : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_486 = _T_479 ? _T_409 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_487 = _T_483 ? _T_412 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_488 = _T_485 | _T_486; // @[Mux.scala 27:72]
  wire [18:0] _T_489 = _T_488 | _T_487; // @[Mux.scala 27:72]
  wire [31:0] bp_rs_call_target_f = {_T_489,_T_464[11:0],1'h0}; // @[Cat.scala 29:58]
  wire  _T_493 = ~btb_rd_ret_f; // @[ifu_bp_ctl.scala 379:33]
  wire  _T_494 = btb_rd_call_f & _T_493; // @[ifu_bp_ctl.scala 379:31]
  wire  rs_push = _T_494 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 379:47]
  wire  rs_pop = _T_436 & io_ifu_bp_hit_taken_f; // @[ifu_bp_ctl.scala 380:46]
  wire  _T_497 = ~rs_push; // @[ifu_bp_ctl.scala 381:17]
  wire  _T_498 = ~rs_pop; // @[ifu_bp_ctl.scala 381:28]
  wire  rs_hold = _T_497 & _T_498; // @[ifu_bp_ctl.scala 381:26]
  wire  rsenable_0 = ~rs_hold; // @[ifu_bp_ctl.scala 383:60]
  wire  rsenable_1 = rs_push | rs_pop; // @[ifu_bp_ctl.scala 383:119]
  wire [31:0] _T_501 = {bp_rs_call_target_f[31:1],1'h1}; // @[Cat.scala 29:58]
  wire [31:0] _T_503 = rs_push ? _T_501 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_1; // @[Reg.scala 27:20]
  wire [31:0] _T_504 = rs_pop ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_0 = _T_503 | _T_504; // @[Mux.scala 27:72]
  wire [31:0] _T_508 = rs_push ? rets_out_0 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_2; // @[Reg.scala 27:20]
  wire [31:0] _T_509 = rs_pop ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_1 = _T_508 | _T_509; // @[Mux.scala 27:72]
  wire [31:0] _T_513 = rs_push ? rets_out_1 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_3; // @[Reg.scala 27:20]
  wire [31:0] _T_514 = rs_pop ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_2 = _T_513 | _T_514; // @[Mux.scala 27:72]
  wire [31:0] _T_518 = rs_push ? rets_out_2 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_4; // @[Reg.scala 27:20]
  wire [31:0] _T_519 = rs_pop ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_3 = _T_518 | _T_519; // @[Mux.scala 27:72]
  wire [31:0] _T_523 = rs_push ? rets_out_3 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_5; // @[Reg.scala 27:20]
  wire [31:0] _T_524 = rs_pop ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_4 = _T_523 | _T_524; // @[Mux.scala 27:72]
  wire [31:0] _T_528 = rs_push ? rets_out_4 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_6; // @[Reg.scala 27:20]
  wire [31:0] _T_529 = rs_pop ? rets_out_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_5 = _T_528 | _T_529; // @[Mux.scala 27:72]
  wire [31:0] _T_533 = rs_push ? rets_out_5 : 32'h0; // @[Mux.scala 27:72]
  reg [31:0] rets_out_7; // @[Reg.scala 27:20]
  wire [31:0] _T_534 = rs_pop ? rets_out_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] rets_in_6 = _T_533 | _T_534; // @[Mux.scala 27:72]
  wire  _T_552 = ~dec_tlu_error_wb; // @[ifu_bp_ctl.scala 395:35]
  wire  btb_valid = exu_mp_valid & _T_552; // @[ifu_bp_ctl.scala 395:32]
  wire  _T_553 = io_exu_bp_exu_mp_pkt_bits_pcall | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 399:89]
  wire  _T_554 = io_exu_bp_exu_mp_pkt_bits_pret | io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 399:113]
  wire [21:0] btb_wr_data = {io_exu_bp_exu_mp_btag,io_exu_bp_exu_mp_pkt_bits_toffset,io_exu_bp_exu_mp_pkt_bits_pc4,io_exu_bp_exu_mp_pkt_bits_boffset,_T_553,_T_554,btb_valid}; // @[Cat.scala 29:58]
  wire  _T_560 = exu_mp_valid & io_exu_bp_exu_mp_pkt_bits_ataken; // @[ifu_bp_ctl.scala 400:41]
  wire  _T_561 = ~io_exu_bp_exu_mp_pkt_valid; // @[ifu_bp_ctl.scala 400:59]
  wire  exu_mp_valid_write = _T_560 & _T_561; // @[ifu_bp_ctl.scala 400:57]
  wire  middle_of_bank = io_exu_bp_exu_mp_pkt_bits_pc4 ^ io_exu_bp_exu_mp_pkt_bits_boffset; // @[ifu_bp_ctl.scala 401:35]
  wire  _T_562 = ~io_exu_bp_exu_mp_pkt_bits_pcall; // @[ifu_bp_ctl.scala 404:43]
  wire  _T_563 = exu_mp_valid & _T_562; // @[ifu_bp_ctl.scala 404:41]
  wire  _T_564 = ~io_exu_bp_exu_mp_pkt_bits_pret; // @[ifu_bp_ctl.scala 404:58]
  wire  _T_565 = _T_563 & _T_564; // @[ifu_bp_ctl.scala 404:56]
  wire  _T_566 = ~io_exu_bp_exu_mp_pkt_bits_pja; // @[ifu_bp_ctl.scala 404:72]
  wire  _T_567 = _T_565 & _T_566; // @[ifu_bp_ctl.scala 404:70]
  wire [1:0] _T_569 = _T_567 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_570 = ~middle_of_bank; // @[ifu_bp_ctl.scala 404:106]
  wire [1:0] _T_571 = {middle_of_bank,_T_570}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en0 = _T_569 & _T_571; // @[ifu_bp_ctl.scala 404:84]
  wire [1:0] _T_573 = io_dec_bp_dec_tlu_br0_r_pkt_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_574 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_middle; // @[ifu_bp_ctl.scala 405:75]
  wire [1:0] _T_575 = {io_dec_bp_dec_tlu_br0_r_pkt_bits_middle,_T_574}; // @[Cat.scala 29:58]
  wire [1:0] bht_wr_en2 = _T_573 & _T_575; // @[ifu_bp_ctl.scala 405:46]
  wire [9:0] _T_576 = {io_exu_bp_exu_mp_index,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] mp_hashed = _T_576[9:2] ^ io_exu_bp_exu_mp_eghr; // @[lib.scala 56:35]
  wire [9:0] _T_579 = {io_exu_bp_exu_i0_br_index_r,2'h0}; // @[Cat.scala 29:58]
  wire [7:0] br0_hashed_wb = _T_579[9:2] ^ io_exu_bp_exu_i0_br_fghr_r; // @[lib.scala 56:35]
  wire  _T_589 = _T_170 & exu_mp_valid_write; // @[ifu_bp_ctl.scala 425:39]
  wire  _T_591 = _T_589 & _T_552; // @[ifu_bp_ctl.scala 425:60]
  wire  _T_592 = ~io_dec_bp_dec_tlu_br0_r_pkt_bits_way; // @[ifu_bp_ctl.scala 425:87]
  wire  _T_593 = _T_592 & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 425:104]
  wire  btb_wr_en_way0 = _T_591 | _T_593; // @[ifu_bp_ctl.scala 425:83]
  wire  _T_594 = io_exu_bp_exu_mp_pkt_bits_way & exu_mp_valid_write; // @[ifu_bp_ctl.scala 426:36]
  wire  _T_596 = _T_594 & _T_552; // @[ifu_bp_ctl.scala 426:57]
  wire  _T_597 = io_dec_bp_dec_tlu_br0_r_pkt_bits_way & dec_tlu_error_wb; // @[ifu_bp_ctl.scala 426:98]
  wire  btb_wr_en_way1 = _T_596 | _T_597; // @[ifu_bp_ctl.scala 426:80]
  wire [7:0] btb_wr_addr = dec_tlu_error_wb ? io_exu_bp_exu_i0_br_index_r : io_exu_bp_exu_mp_index; // @[ifu_bp_ctl.scala 429:24]
  wire  _T_613 = btb_wr_addr == 8'h0; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_614 = _T_613 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_617 = btb_wr_addr == 8'h1; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_618 = _T_617 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_621 = btb_wr_addr == 8'h2; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_622 = _T_621 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_625 = btb_wr_addr == 8'h3; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_626 = _T_625 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_629 = btb_wr_addr == 8'h4; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_630 = _T_629 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_633 = btb_wr_addr == 8'h5; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_634 = _T_633 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_637 = btb_wr_addr == 8'h6; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_638 = _T_637 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_641 = btb_wr_addr == 8'h7; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_642 = _T_641 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_645 = btb_wr_addr == 8'h8; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_646 = _T_645 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_649 = btb_wr_addr == 8'h9; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_650 = _T_649 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_653 = btb_wr_addr == 8'ha; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_654 = _T_653 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_657 = btb_wr_addr == 8'hb; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_658 = _T_657 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_661 = btb_wr_addr == 8'hc; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_662 = _T_661 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_665 = btb_wr_addr == 8'hd; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_666 = _T_665 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_669 = btb_wr_addr == 8'he; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_670 = _T_669 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_673 = btb_wr_addr == 8'hf; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_674 = _T_673 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_677 = btb_wr_addr == 8'h10; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_678 = _T_677 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_681 = btb_wr_addr == 8'h11; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_682 = _T_681 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_685 = btb_wr_addr == 8'h12; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_686 = _T_685 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_689 = btb_wr_addr == 8'h13; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_690 = _T_689 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_693 = btb_wr_addr == 8'h14; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_694 = _T_693 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_697 = btb_wr_addr == 8'h15; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_698 = _T_697 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_701 = btb_wr_addr == 8'h16; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_702 = _T_701 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_705 = btb_wr_addr == 8'h17; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_706 = _T_705 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_709 = btb_wr_addr == 8'h18; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_710 = _T_709 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_713 = btb_wr_addr == 8'h19; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_714 = _T_713 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_717 = btb_wr_addr == 8'h1a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_718 = _T_717 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_721 = btb_wr_addr == 8'h1b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_722 = _T_721 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_725 = btb_wr_addr == 8'h1c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_726 = _T_725 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_729 = btb_wr_addr == 8'h1d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_730 = _T_729 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_733 = btb_wr_addr == 8'h1e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_734 = _T_733 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_737 = btb_wr_addr == 8'h1f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_738 = _T_737 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_741 = btb_wr_addr == 8'h20; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_742 = _T_741 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_745 = btb_wr_addr == 8'h21; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_746 = _T_745 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_749 = btb_wr_addr == 8'h22; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_750 = _T_749 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_753 = btb_wr_addr == 8'h23; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_754 = _T_753 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_757 = btb_wr_addr == 8'h24; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_758 = _T_757 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_761 = btb_wr_addr == 8'h25; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_762 = _T_761 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_765 = btb_wr_addr == 8'h26; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_766 = _T_765 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_769 = btb_wr_addr == 8'h27; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_770 = _T_769 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_773 = btb_wr_addr == 8'h28; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_774 = _T_773 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_777 = btb_wr_addr == 8'h29; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_778 = _T_777 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_781 = btb_wr_addr == 8'h2a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_782 = _T_781 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_785 = btb_wr_addr == 8'h2b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_786 = _T_785 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_789 = btb_wr_addr == 8'h2c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_790 = _T_789 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_793 = btb_wr_addr == 8'h2d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_794 = _T_793 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_797 = btb_wr_addr == 8'h2e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_798 = _T_797 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_801 = btb_wr_addr == 8'h2f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_802 = _T_801 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_805 = btb_wr_addr == 8'h30; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_806 = _T_805 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_809 = btb_wr_addr == 8'h31; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_810 = _T_809 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_813 = btb_wr_addr == 8'h32; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_814 = _T_813 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_817 = btb_wr_addr == 8'h33; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_818 = _T_817 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_821 = btb_wr_addr == 8'h34; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_822 = _T_821 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_825 = btb_wr_addr == 8'h35; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_826 = _T_825 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_829 = btb_wr_addr == 8'h36; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_830 = _T_829 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_833 = btb_wr_addr == 8'h37; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_834 = _T_833 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_837 = btb_wr_addr == 8'h38; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_838 = _T_837 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_841 = btb_wr_addr == 8'h39; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_842 = _T_841 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_845 = btb_wr_addr == 8'h3a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_846 = _T_845 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_849 = btb_wr_addr == 8'h3b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_850 = _T_849 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_853 = btb_wr_addr == 8'h3c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_854 = _T_853 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_857 = btb_wr_addr == 8'h3d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_858 = _T_857 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_861 = btb_wr_addr == 8'h3e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_862 = _T_861 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_865 = btb_wr_addr == 8'h3f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_866 = _T_865 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_869 = btb_wr_addr == 8'h40; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_870 = _T_869 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_873 = btb_wr_addr == 8'h41; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_874 = _T_873 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_877 = btb_wr_addr == 8'h42; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_878 = _T_877 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_881 = btb_wr_addr == 8'h43; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_882 = _T_881 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_885 = btb_wr_addr == 8'h44; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_886 = _T_885 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_889 = btb_wr_addr == 8'h45; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_890 = _T_889 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_893 = btb_wr_addr == 8'h46; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_894 = _T_893 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_897 = btb_wr_addr == 8'h47; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_898 = _T_897 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_901 = btb_wr_addr == 8'h48; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_902 = _T_901 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_905 = btb_wr_addr == 8'h49; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_906 = _T_905 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_909 = btb_wr_addr == 8'h4a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_910 = _T_909 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_913 = btb_wr_addr == 8'h4b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_914 = _T_913 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_917 = btb_wr_addr == 8'h4c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_918 = _T_917 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_921 = btb_wr_addr == 8'h4d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_922 = _T_921 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_925 = btb_wr_addr == 8'h4e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_926 = _T_925 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_929 = btb_wr_addr == 8'h4f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_930 = _T_929 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_933 = btb_wr_addr == 8'h50; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_934 = _T_933 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_937 = btb_wr_addr == 8'h51; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_938 = _T_937 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_941 = btb_wr_addr == 8'h52; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_942 = _T_941 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_945 = btb_wr_addr == 8'h53; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_946 = _T_945 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_949 = btb_wr_addr == 8'h54; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_950 = _T_949 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_953 = btb_wr_addr == 8'h55; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_954 = _T_953 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_957 = btb_wr_addr == 8'h56; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_958 = _T_957 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_961 = btb_wr_addr == 8'h57; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_962 = _T_961 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_965 = btb_wr_addr == 8'h58; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_966 = _T_965 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_969 = btb_wr_addr == 8'h59; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_970 = _T_969 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_973 = btb_wr_addr == 8'h5a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_974 = _T_973 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_977 = btb_wr_addr == 8'h5b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_978 = _T_977 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_981 = btb_wr_addr == 8'h5c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_982 = _T_981 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_985 = btb_wr_addr == 8'h5d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_986 = _T_985 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_989 = btb_wr_addr == 8'h5e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_990 = _T_989 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_993 = btb_wr_addr == 8'h5f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_994 = _T_993 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_997 = btb_wr_addr == 8'h60; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_998 = _T_997 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1001 = btb_wr_addr == 8'h61; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1002 = _T_1001 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1005 = btb_wr_addr == 8'h62; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1006 = _T_1005 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1009 = btb_wr_addr == 8'h63; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1010 = _T_1009 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1013 = btb_wr_addr == 8'h64; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1014 = _T_1013 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1017 = btb_wr_addr == 8'h65; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1018 = _T_1017 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1021 = btb_wr_addr == 8'h66; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1022 = _T_1021 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1025 = btb_wr_addr == 8'h67; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1026 = _T_1025 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1029 = btb_wr_addr == 8'h68; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1030 = _T_1029 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1033 = btb_wr_addr == 8'h69; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1034 = _T_1033 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1037 = btb_wr_addr == 8'h6a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1038 = _T_1037 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1041 = btb_wr_addr == 8'h6b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1042 = _T_1041 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1045 = btb_wr_addr == 8'h6c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1046 = _T_1045 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1049 = btb_wr_addr == 8'h6d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1050 = _T_1049 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1053 = btb_wr_addr == 8'h6e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1054 = _T_1053 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1057 = btb_wr_addr == 8'h6f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1058 = _T_1057 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1061 = btb_wr_addr == 8'h70; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1062 = _T_1061 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1065 = btb_wr_addr == 8'h71; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1066 = _T_1065 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1069 = btb_wr_addr == 8'h72; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1070 = _T_1069 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1073 = btb_wr_addr == 8'h73; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1074 = _T_1073 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1077 = btb_wr_addr == 8'h74; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1078 = _T_1077 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1081 = btb_wr_addr == 8'h75; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1082 = _T_1081 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1085 = btb_wr_addr == 8'h76; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1086 = _T_1085 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1089 = btb_wr_addr == 8'h77; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1090 = _T_1089 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1093 = btb_wr_addr == 8'h78; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1094 = _T_1093 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1097 = btb_wr_addr == 8'h79; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1098 = _T_1097 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1101 = btb_wr_addr == 8'h7a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1102 = _T_1101 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1105 = btb_wr_addr == 8'h7b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1106 = _T_1105 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1109 = btb_wr_addr == 8'h7c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1110 = _T_1109 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1113 = btb_wr_addr == 8'h7d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1114 = _T_1113 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1117 = btb_wr_addr == 8'h7e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1118 = _T_1117 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1121 = btb_wr_addr == 8'h7f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1122 = _T_1121 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1125 = btb_wr_addr == 8'h80; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1126 = _T_1125 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1129 = btb_wr_addr == 8'h81; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1130 = _T_1129 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1133 = btb_wr_addr == 8'h82; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1134 = _T_1133 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1137 = btb_wr_addr == 8'h83; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1138 = _T_1137 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1141 = btb_wr_addr == 8'h84; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1142 = _T_1141 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1145 = btb_wr_addr == 8'h85; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1146 = _T_1145 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1149 = btb_wr_addr == 8'h86; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1150 = _T_1149 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1153 = btb_wr_addr == 8'h87; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1154 = _T_1153 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1157 = btb_wr_addr == 8'h88; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1158 = _T_1157 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1161 = btb_wr_addr == 8'h89; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1162 = _T_1161 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1165 = btb_wr_addr == 8'h8a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1166 = _T_1165 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1169 = btb_wr_addr == 8'h8b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1170 = _T_1169 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1173 = btb_wr_addr == 8'h8c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1174 = _T_1173 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1177 = btb_wr_addr == 8'h8d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1178 = _T_1177 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1181 = btb_wr_addr == 8'h8e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1182 = _T_1181 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1185 = btb_wr_addr == 8'h8f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1186 = _T_1185 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1189 = btb_wr_addr == 8'h90; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1190 = _T_1189 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1193 = btb_wr_addr == 8'h91; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1194 = _T_1193 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1197 = btb_wr_addr == 8'h92; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1198 = _T_1197 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1201 = btb_wr_addr == 8'h93; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1202 = _T_1201 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1205 = btb_wr_addr == 8'h94; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1206 = _T_1205 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1209 = btb_wr_addr == 8'h95; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1210 = _T_1209 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1213 = btb_wr_addr == 8'h96; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1214 = _T_1213 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1217 = btb_wr_addr == 8'h97; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1218 = _T_1217 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1221 = btb_wr_addr == 8'h98; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1222 = _T_1221 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1225 = btb_wr_addr == 8'h99; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1226 = _T_1225 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1229 = btb_wr_addr == 8'h9a; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1230 = _T_1229 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1233 = btb_wr_addr == 8'h9b; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1234 = _T_1233 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1237 = btb_wr_addr == 8'h9c; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1238 = _T_1237 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1241 = btb_wr_addr == 8'h9d; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1242 = _T_1241 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1245 = btb_wr_addr == 8'h9e; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1246 = _T_1245 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1249 = btb_wr_addr == 8'h9f; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1250 = _T_1249 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1253 = btb_wr_addr == 8'ha0; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1254 = _T_1253 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1257 = btb_wr_addr == 8'ha1; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1258 = _T_1257 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1261 = btb_wr_addr == 8'ha2; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1262 = _T_1261 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1265 = btb_wr_addr == 8'ha3; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1266 = _T_1265 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1269 = btb_wr_addr == 8'ha4; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1270 = _T_1269 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1273 = btb_wr_addr == 8'ha5; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1274 = _T_1273 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1277 = btb_wr_addr == 8'ha6; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1278 = _T_1277 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1281 = btb_wr_addr == 8'ha7; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1282 = _T_1281 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1285 = btb_wr_addr == 8'ha8; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1286 = _T_1285 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1289 = btb_wr_addr == 8'ha9; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1290 = _T_1289 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1293 = btb_wr_addr == 8'haa; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1294 = _T_1293 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1297 = btb_wr_addr == 8'hab; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1298 = _T_1297 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1301 = btb_wr_addr == 8'hac; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1302 = _T_1301 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1305 = btb_wr_addr == 8'had; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1306 = _T_1305 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1309 = btb_wr_addr == 8'hae; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1310 = _T_1309 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1313 = btb_wr_addr == 8'haf; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1314 = _T_1313 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1317 = btb_wr_addr == 8'hb0; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1318 = _T_1317 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1321 = btb_wr_addr == 8'hb1; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1322 = _T_1321 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1325 = btb_wr_addr == 8'hb2; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1326 = _T_1325 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1329 = btb_wr_addr == 8'hb3; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1330 = _T_1329 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1333 = btb_wr_addr == 8'hb4; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1334 = _T_1333 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1337 = btb_wr_addr == 8'hb5; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1338 = _T_1337 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1341 = btb_wr_addr == 8'hb6; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1342 = _T_1341 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1345 = btb_wr_addr == 8'hb7; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1346 = _T_1345 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1349 = btb_wr_addr == 8'hb8; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1350 = _T_1349 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1353 = btb_wr_addr == 8'hb9; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1354 = _T_1353 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1357 = btb_wr_addr == 8'hba; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1358 = _T_1357 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1361 = btb_wr_addr == 8'hbb; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1362 = _T_1361 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1365 = btb_wr_addr == 8'hbc; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1366 = _T_1365 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1369 = btb_wr_addr == 8'hbd; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1370 = _T_1369 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1373 = btb_wr_addr == 8'hbe; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1374 = _T_1373 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1377 = btb_wr_addr == 8'hbf; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1378 = _T_1377 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1381 = btb_wr_addr == 8'hc0; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1382 = _T_1381 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1385 = btb_wr_addr == 8'hc1; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1386 = _T_1385 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1389 = btb_wr_addr == 8'hc2; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1390 = _T_1389 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1393 = btb_wr_addr == 8'hc3; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1394 = _T_1393 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1397 = btb_wr_addr == 8'hc4; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1398 = _T_1397 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1401 = btb_wr_addr == 8'hc5; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1402 = _T_1401 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1405 = btb_wr_addr == 8'hc6; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1406 = _T_1405 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1409 = btb_wr_addr == 8'hc7; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1410 = _T_1409 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1413 = btb_wr_addr == 8'hc8; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1414 = _T_1413 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1417 = btb_wr_addr == 8'hc9; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1418 = _T_1417 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1421 = btb_wr_addr == 8'hca; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1422 = _T_1421 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1425 = btb_wr_addr == 8'hcb; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1426 = _T_1425 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1429 = btb_wr_addr == 8'hcc; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1430 = _T_1429 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1433 = btb_wr_addr == 8'hcd; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1434 = _T_1433 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1437 = btb_wr_addr == 8'hce; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1438 = _T_1437 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1441 = btb_wr_addr == 8'hcf; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1442 = _T_1441 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1445 = btb_wr_addr == 8'hd0; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1446 = _T_1445 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1449 = btb_wr_addr == 8'hd1; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1450 = _T_1449 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1453 = btb_wr_addr == 8'hd2; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1454 = _T_1453 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1457 = btb_wr_addr == 8'hd3; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1458 = _T_1457 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1461 = btb_wr_addr == 8'hd4; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1462 = _T_1461 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1465 = btb_wr_addr == 8'hd5; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1466 = _T_1465 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1469 = btb_wr_addr == 8'hd6; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1470 = _T_1469 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1473 = btb_wr_addr == 8'hd7; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1474 = _T_1473 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1477 = btb_wr_addr == 8'hd8; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1478 = _T_1477 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1481 = btb_wr_addr == 8'hd9; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1482 = _T_1481 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1485 = btb_wr_addr == 8'hda; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1486 = _T_1485 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1489 = btb_wr_addr == 8'hdb; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1490 = _T_1489 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1493 = btb_wr_addr == 8'hdc; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1494 = _T_1493 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1497 = btb_wr_addr == 8'hdd; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1498 = _T_1497 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1501 = btb_wr_addr == 8'hde; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1502 = _T_1501 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1505 = btb_wr_addr == 8'hdf; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1506 = _T_1505 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1509 = btb_wr_addr == 8'he0; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1510 = _T_1509 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1513 = btb_wr_addr == 8'he1; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1514 = _T_1513 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1517 = btb_wr_addr == 8'he2; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1518 = _T_1517 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1521 = btb_wr_addr == 8'he3; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1522 = _T_1521 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1525 = btb_wr_addr == 8'he4; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1526 = _T_1525 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1529 = btb_wr_addr == 8'he5; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1530 = _T_1529 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1533 = btb_wr_addr == 8'he6; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1534 = _T_1533 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1537 = btb_wr_addr == 8'he7; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1538 = _T_1537 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1541 = btb_wr_addr == 8'he8; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1542 = _T_1541 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1545 = btb_wr_addr == 8'he9; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1546 = _T_1545 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1549 = btb_wr_addr == 8'hea; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1550 = _T_1549 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1553 = btb_wr_addr == 8'heb; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1554 = _T_1553 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1557 = btb_wr_addr == 8'hec; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1558 = _T_1557 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1561 = btb_wr_addr == 8'hed; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1562 = _T_1561 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1565 = btb_wr_addr == 8'hee; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1566 = _T_1565 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1569 = btb_wr_addr == 8'hef; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1570 = _T_1569 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1573 = btb_wr_addr == 8'hf0; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1574 = _T_1573 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1577 = btb_wr_addr == 8'hf1; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1578 = _T_1577 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1581 = btb_wr_addr == 8'hf2; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1582 = _T_1581 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1585 = btb_wr_addr == 8'hf3; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1586 = _T_1585 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1589 = btb_wr_addr == 8'hf4; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1590 = _T_1589 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1593 = btb_wr_addr == 8'hf5; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1594 = _T_1593 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1597 = btb_wr_addr == 8'hf6; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1598 = _T_1597 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1601 = btb_wr_addr == 8'hf7; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1602 = _T_1601 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1605 = btb_wr_addr == 8'hf8; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1606 = _T_1605 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1609 = btb_wr_addr == 8'hf9; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1610 = _T_1609 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1613 = btb_wr_addr == 8'hfa; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1614 = _T_1613 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1617 = btb_wr_addr == 8'hfb; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1618 = _T_1617 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1621 = btb_wr_addr == 8'hfc; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1622 = _T_1621 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1625 = btb_wr_addr == 8'hfd; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1626 = _T_1625 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1629 = btb_wr_addr == 8'hfe; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1630 = _T_1629 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1633 = btb_wr_addr == 8'hff; // @[ifu_bp_ctl.scala 434:95]
  wire  _T_1634 = _T_1633 & btb_wr_en_way0; // @[ifu_bp_ctl.scala 434:104]
  wire  _T_1638 = _T_613 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1642 = _T_617 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1646 = _T_621 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1650 = _T_625 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1654 = _T_629 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1658 = _T_633 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1662 = _T_637 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1666 = _T_641 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1670 = _T_645 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1674 = _T_649 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1678 = _T_653 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1682 = _T_657 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1686 = _T_661 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1690 = _T_665 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1694 = _T_669 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1698 = _T_673 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1702 = _T_677 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1706 = _T_681 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1710 = _T_685 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1714 = _T_689 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1718 = _T_693 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1722 = _T_697 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1726 = _T_701 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1730 = _T_705 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1734 = _T_709 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1738 = _T_713 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1742 = _T_717 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1746 = _T_721 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1750 = _T_725 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1754 = _T_729 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1758 = _T_733 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1762 = _T_737 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1766 = _T_741 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1770 = _T_745 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1774 = _T_749 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1778 = _T_753 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1782 = _T_757 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1786 = _T_761 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1790 = _T_765 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1794 = _T_769 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1798 = _T_773 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1802 = _T_777 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1806 = _T_781 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1810 = _T_785 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1814 = _T_789 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1818 = _T_793 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1822 = _T_797 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1826 = _T_801 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1830 = _T_805 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1834 = _T_809 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1838 = _T_813 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1842 = _T_817 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1846 = _T_821 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1850 = _T_825 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1854 = _T_829 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1858 = _T_833 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1862 = _T_837 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1866 = _T_841 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1870 = _T_845 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1874 = _T_849 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1878 = _T_853 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1882 = _T_857 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1886 = _T_861 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1890 = _T_865 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1894 = _T_869 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1898 = _T_873 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1902 = _T_877 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1906 = _T_881 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1910 = _T_885 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1914 = _T_889 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1918 = _T_893 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1922 = _T_897 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1926 = _T_901 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1930 = _T_905 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1934 = _T_909 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1938 = _T_913 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1942 = _T_917 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1946 = _T_921 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1950 = _T_925 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1954 = _T_929 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1958 = _T_933 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1962 = _T_937 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1966 = _T_941 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1970 = _T_945 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1974 = _T_949 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1978 = _T_953 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1982 = _T_957 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1986 = _T_961 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1990 = _T_965 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1994 = _T_969 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_1998 = _T_973 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2002 = _T_977 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2006 = _T_981 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2010 = _T_985 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2014 = _T_989 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2018 = _T_993 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2022 = _T_997 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2026 = _T_1001 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2030 = _T_1005 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2034 = _T_1009 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2038 = _T_1013 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2042 = _T_1017 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2046 = _T_1021 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2050 = _T_1025 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2054 = _T_1029 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2058 = _T_1033 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2062 = _T_1037 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2066 = _T_1041 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2070 = _T_1045 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2074 = _T_1049 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2078 = _T_1053 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2082 = _T_1057 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2086 = _T_1061 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2090 = _T_1065 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2094 = _T_1069 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2098 = _T_1073 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2102 = _T_1077 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2106 = _T_1081 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2110 = _T_1085 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2114 = _T_1089 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2118 = _T_1093 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2122 = _T_1097 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2126 = _T_1101 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2130 = _T_1105 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2134 = _T_1109 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2138 = _T_1113 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2142 = _T_1117 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2146 = _T_1121 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2150 = _T_1125 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2154 = _T_1129 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2158 = _T_1133 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2162 = _T_1137 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2166 = _T_1141 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2170 = _T_1145 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2174 = _T_1149 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2178 = _T_1153 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2182 = _T_1157 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2186 = _T_1161 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2190 = _T_1165 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2194 = _T_1169 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2198 = _T_1173 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2202 = _T_1177 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2206 = _T_1181 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2210 = _T_1185 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2214 = _T_1189 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2218 = _T_1193 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2222 = _T_1197 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2226 = _T_1201 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2230 = _T_1205 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2234 = _T_1209 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2238 = _T_1213 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2242 = _T_1217 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2246 = _T_1221 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2250 = _T_1225 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2254 = _T_1229 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2258 = _T_1233 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2262 = _T_1237 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2266 = _T_1241 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2270 = _T_1245 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2274 = _T_1249 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2278 = _T_1253 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2282 = _T_1257 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2286 = _T_1261 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2290 = _T_1265 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2294 = _T_1269 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2298 = _T_1273 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2302 = _T_1277 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2306 = _T_1281 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2310 = _T_1285 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2314 = _T_1289 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2318 = _T_1293 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2322 = _T_1297 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2326 = _T_1301 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2330 = _T_1305 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2334 = _T_1309 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2338 = _T_1313 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2342 = _T_1317 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2346 = _T_1321 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2350 = _T_1325 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2354 = _T_1329 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2358 = _T_1333 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2362 = _T_1337 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2366 = _T_1341 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2370 = _T_1345 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2374 = _T_1349 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2378 = _T_1353 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2382 = _T_1357 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2386 = _T_1361 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2390 = _T_1365 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2394 = _T_1369 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2398 = _T_1373 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2402 = _T_1377 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2406 = _T_1381 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2410 = _T_1385 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2414 = _T_1389 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2418 = _T_1393 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2422 = _T_1397 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2426 = _T_1401 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2430 = _T_1405 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2434 = _T_1409 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2438 = _T_1413 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2442 = _T_1417 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2446 = _T_1421 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2450 = _T_1425 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2454 = _T_1429 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2458 = _T_1433 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2462 = _T_1437 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2466 = _T_1441 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2470 = _T_1445 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2474 = _T_1449 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2478 = _T_1453 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2482 = _T_1457 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2486 = _T_1461 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2490 = _T_1465 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2494 = _T_1469 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2498 = _T_1473 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2502 = _T_1477 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2506 = _T_1481 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2510 = _T_1485 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2514 = _T_1489 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2518 = _T_1493 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2522 = _T_1497 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2526 = _T_1501 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2530 = _T_1505 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2534 = _T_1509 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2538 = _T_1513 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2542 = _T_1517 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2546 = _T_1521 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2550 = _T_1525 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2554 = _T_1529 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2558 = _T_1533 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2562 = _T_1537 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2566 = _T_1541 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2570 = _T_1545 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2574 = _T_1549 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2578 = _T_1553 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2582 = _T_1557 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2586 = _T_1561 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2590 = _T_1565 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2594 = _T_1569 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2598 = _T_1573 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2602 = _T_1577 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2606 = _T_1581 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2610 = _T_1585 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2614 = _T_1589 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2618 = _T_1593 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2622 = _T_1597 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2626 = _T_1601 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2630 = _T_1605 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2634 = _T_1609 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2638 = _T_1613 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2642 = _T_1617 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2646 = _T_1621 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2650 = _T_1625 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2654 = _T_1629 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_2658 = _T_1633 & btb_wr_en_way1; // @[ifu_bp_ctl.scala 435:104]
  wire  _T_6759 = mp_hashed[7:4] == 4'h0; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6761 = bht_wr_en0[0] & _T_6759; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6764 = br0_hashed_wb[7:4] == 4'h0; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6766 = bht_wr_en2[0] & _T_6764; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6770 = mp_hashed[7:4] == 4'h1; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6772 = bht_wr_en0[0] & _T_6770; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6775 = br0_hashed_wb[7:4] == 4'h1; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6777 = bht_wr_en2[0] & _T_6775; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6781 = mp_hashed[7:4] == 4'h2; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6783 = bht_wr_en0[0] & _T_6781; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6786 = br0_hashed_wb[7:4] == 4'h2; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6788 = bht_wr_en2[0] & _T_6786; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6792 = mp_hashed[7:4] == 4'h3; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6794 = bht_wr_en0[0] & _T_6792; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6797 = br0_hashed_wb[7:4] == 4'h3; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6799 = bht_wr_en2[0] & _T_6797; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6803 = mp_hashed[7:4] == 4'h4; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6805 = bht_wr_en0[0] & _T_6803; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6808 = br0_hashed_wb[7:4] == 4'h4; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6810 = bht_wr_en2[0] & _T_6808; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6814 = mp_hashed[7:4] == 4'h5; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6816 = bht_wr_en0[0] & _T_6814; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6819 = br0_hashed_wb[7:4] == 4'h5; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6821 = bht_wr_en2[0] & _T_6819; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6825 = mp_hashed[7:4] == 4'h6; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6827 = bht_wr_en0[0] & _T_6825; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6830 = br0_hashed_wb[7:4] == 4'h6; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6832 = bht_wr_en2[0] & _T_6830; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6836 = mp_hashed[7:4] == 4'h7; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6838 = bht_wr_en0[0] & _T_6836; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6841 = br0_hashed_wb[7:4] == 4'h7; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6843 = bht_wr_en2[0] & _T_6841; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6847 = mp_hashed[7:4] == 4'h8; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6849 = bht_wr_en0[0] & _T_6847; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6852 = br0_hashed_wb[7:4] == 4'h8; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6854 = bht_wr_en2[0] & _T_6852; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6858 = mp_hashed[7:4] == 4'h9; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6860 = bht_wr_en0[0] & _T_6858; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6863 = br0_hashed_wb[7:4] == 4'h9; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6865 = bht_wr_en2[0] & _T_6863; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6869 = mp_hashed[7:4] == 4'ha; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6871 = bht_wr_en0[0] & _T_6869; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6874 = br0_hashed_wb[7:4] == 4'ha; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6876 = bht_wr_en2[0] & _T_6874; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6880 = mp_hashed[7:4] == 4'hb; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6882 = bht_wr_en0[0] & _T_6880; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6885 = br0_hashed_wb[7:4] == 4'hb; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6887 = bht_wr_en2[0] & _T_6885; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6891 = mp_hashed[7:4] == 4'hc; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6893 = bht_wr_en0[0] & _T_6891; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6896 = br0_hashed_wb[7:4] == 4'hc; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6898 = bht_wr_en2[0] & _T_6896; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6902 = mp_hashed[7:4] == 4'hd; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6904 = bht_wr_en0[0] & _T_6902; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6907 = br0_hashed_wb[7:4] == 4'hd; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6909 = bht_wr_en2[0] & _T_6907; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6913 = mp_hashed[7:4] == 4'he; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6915 = bht_wr_en0[0] & _T_6913; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6918 = br0_hashed_wb[7:4] == 4'he; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6920 = bht_wr_en2[0] & _T_6918; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6924 = mp_hashed[7:4] == 4'hf; // @[ifu_bp_ctl.scala 507:109]
  wire  _T_6926 = bht_wr_en0[0] & _T_6924; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6929 = br0_hashed_wb[7:4] == 4'hf; // @[ifu_bp_ctl.scala 508:109]
  wire  _T_6931 = bht_wr_en2[0] & _T_6929; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6937 = bht_wr_en0[1] & _T_6759; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6942 = bht_wr_en2[1] & _T_6764; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6948 = bht_wr_en0[1] & _T_6770; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6953 = bht_wr_en2[1] & _T_6775; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6959 = bht_wr_en0[1] & _T_6781; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6964 = bht_wr_en2[1] & _T_6786; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6970 = bht_wr_en0[1] & _T_6792; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6975 = bht_wr_en2[1] & _T_6797; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6981 = bht_wr_en0[1] & _T_6803; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6986 = bht_wr_en2[1] & _T_6808; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_6992 = bht_wr_en0[1] & _T_6814; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_6997 = bht_wr_en2[1] & _T_6819; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7003 = bht_wr_en0[1] & _T_6825; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7008 = bht_wr_en2[1] & _T_6830; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7014 = bht_wr_en0[1] & _T_6836; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7019 = bht_wr_en2[1] & _T_6841; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7025 = bht_wr_en0[1] & _T_6847; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7030 = bht_wr_en2[1] & _T_6852; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7036 = bht_wr_en0[1] & _T_6858; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7041 = bht_wr_en2[1] & _T_6863; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7047 = bht_wr_en0[1] & _T_6869; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7052 = bht_wr_en2[1] & _T_6874; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7058 = bht_wr_en0[1] & _T_6880; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7063 = bht_wr_en2[1] & _T_6885; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7069 = bht_wr_en0[1] & _T_6891; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7074 = bht_wr_en2[1] & _T_6896; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7080 = bht_wr_en0[1] & _T_6902; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7085 = bht_wr_en2[1] & _T_6907; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7091 = bht_wr_en0[1] & _T_6913; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7096 = bht_wr_en2[1] & _T_6918; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7102 = bht_wr_en0[1] & _T_6924; // @[ifu_bp_ctl.scala 507:44]
  wire  _T_7107 = bht_wr_en2[1] & _T_6929; // @[ifu_bp_ctl.scala 508:44]
  wire  _T_7111 = br0_hashed_wb[3:0] == 4'h0; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7112 = bht_wr_en2[0] & _T_7111; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7116 = _T_7112 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7120 = br0_hashed_wb[3:0] == 4'h1; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7121 = bht_wr_en2[0] & _T_7120; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7125 = _T_7121 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7129 = br0_hashed_wb[3:0] == 4'h2; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7130 = bht_wr_en2[0] & _T_7129; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7134 = _T_7130 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7138 = br0_hashed_wb[3:0] == 4'h3; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7139 = bht_wr_en2[0] & _T_7138; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7143 = _T_7139 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7147 = br0_hashed_wb[3:0] == 4'h4; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7148 = bht_wr_en2[0] & _T_7147; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7152 = _T_7148 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7156 = br0_hashed_wb[3:0] == 4'h5; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7157 = bht_wr_en2[0] & _T_7156; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7161 = _T_7157 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7165 = br0_hashed_wb[3:0] == 4'h6; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7166 = bht_wr_en2[0] & _T_7165; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7170 = _T_7166 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7174 = br0_hashed_wb[3:0] == 4'h7; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7175 = bht_wr_en2[0] & _T_7174; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7179 = _T_7175 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7183 = br0_hashed_wb[3:0] == 4'h8; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7184 = bht_wr_en2[0] & _T_7183; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7188 = _T_7184 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7192 = br0_hashed_wb[3:0] == 4'h9; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7193 = bht_wr_en2[0] & _T_7192; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7197 = _T_7193 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7201 = br0_hashed_wb[3:0] == 4'ha; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7202 = bht_wr_en2[0] & _T_7201; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7206 = _T_7202 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7210 = br0_hashed_wb[3:0] == 4'hb; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7211 = bht_wr_en2[0] & _T_7210; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7215 = _T_7211 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7219 = br0_hashed_wb[3:0] == 4'hc; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7220 = bht_wr_en2[0] & _T_7219; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7224 = _T_7220 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7228 = br0_hashed_wb[3:0] == 4'hd; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7229 = bht_wr_en2[0] & _T_7228; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7233 = _T_7229 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7237 = br0_hashed_wb[3:0] == 4'he; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7238 = bht_wr_en2[0] & _T_7237; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7242 = _T_7238 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7246 = br0_hashed_wb[3:0] == 4'hf; // @[ifu_bp_ctl.scala 512:74]
  wire  _T_7247 = bht_wr_en2[0] & _T_7246; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_7251 = _T_7247 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7260 = _T_7112 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7269 = _T_7121 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7278 = _T_7130 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7287 = _T_7139 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7296 = _T_7148 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7305 = _T_7157 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7314 = _T_7166 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7323 = _T_7175 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7332 = _T_7184 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7341 = _T_7193 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7350 = _T_7202 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7359 = _T_7211 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7368 = _T_7220 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7377 = _T_7229 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7386 = _T_7238 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7395 = _T_7247 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7404 = _T_7112 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7413 = _T_7121 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7422 = _T_7130 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7431 = _T_7139 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7440 = _T_7148 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7449 = _T_7157 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7458 = _T_7166 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7467 = _T_7175 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7476 = _T_7184 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7485 = _T_7193 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7494 = _T_7202 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7503 = _T_7211 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7512 = _T_7220 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7521 = _T_7229 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7530 = _T_7238 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7539 = _T_7247 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7548 = _T_7112 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7557 = _T_7121 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7566 = _T_7130 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7575 = _T_7139 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7584 = _T_7148 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7593 = _T_7157 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7602 = _T_7166 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7611 = _T_7175 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7620 = _T_7184 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7629 = _T_7193 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7638 = _T_7202 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7647 = _T_7211 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7656 = _T_7220 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7665 = _T_7229 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7674 = _T_7238 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7683 = _T_7247 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7692 = _T_7112 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7701 = _T_7121 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7710 = _T_7130 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7719 = _T_7139 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7728 = _T_7148 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7737 = _T_7157 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7746 = _T_7166 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7755 = _T_7175 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7764 = _T_7184 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7773 = _T_7193 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7782 = _T_7202 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7791 = _T_7211 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7800 = _T_7220 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7809 = _T_7229 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7818 = _T_7238 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7827 = _T_7247 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7836 = _T_7112 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7845 = _T_7121 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7854 = _T_7130 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7863 = _T_7139 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7872 = _T_7148 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7881 = _T_7157 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7890 = _T_7166 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7899 = _T_7175 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7908 = _T_7184 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7917 = _T_7193 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7926 = _T_7202 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7935 = _T_7211 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7944 = _T_7220 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7953 = _T_7229 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7962 = _T_7238 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7971 = _T_7247 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7980 = _T_7112 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7989 = _T_7121 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_7998 = _T_7130 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8007 = _T_7139 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8016 = _T_7148 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8025 = _T_7157 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8034 = _T_7166 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8043 = _T_7175 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8052 = _T_7184 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8061 = _T_7193 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8070 = _T_7202 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8079 = _T_7211 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8088 = _T_7220 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8097 = _T_7229 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8106 = _T_7238 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8115 = _T_7247 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8124 = _T_7112 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8133 = _T_7121 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8142 = _T_7130 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8151 = _T_7139 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8160 = _T_7148 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8169 = _T_7157 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8178 = _T_7166 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8187 = _T_7175 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8196 = _T_7184 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8205 = _T_7193 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8214 = _T_7202 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8223 = _T_7211 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8232 = _T_7220 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8241 = _T_7229 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8250 = _T_7238 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8259 = _T_7247 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8268 = _T_7112 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8277 = _T_7121 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8286 = _T_7130 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8295 = _T_7139 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8304 = _T_7148 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8313 = _T_7157 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8322 = _T_7166 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8331 = _T_7175 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8340 = _T_7184 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8349 = _T_7193 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8358 = _T_7202 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8367 = _T_7211 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8376 = _T_7220 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8385 = _T_7229 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8394 = _T_7238 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8403 = _T_7247 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8412 = _T_7112 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8421 = _T_7121 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8430 = _T_7130 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8439 = _T_7139 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8448 = _T_7148 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8457 = _T_7157 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8466 = _T_7166 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8475 = _T_7175 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8484 = _T_7184 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8493 = _T_7193 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8502 = _T_7202 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8511 = _T_7211 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8520 = _T_7220 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8529 = _T_7229 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8538 = _T_7238 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8547 = _T_7247 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8556 = _T_7112 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8565 = _T_7121 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8574 = _T_7130 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8583 = _T_7139 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8592 = _T_7148 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8601 = _T_7157 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8610 = _T_7166 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8619 = _T_7175 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8628 = _T_7184 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8637 = _T_7193 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8646 = _T_7202 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8655 = _T_7211 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8664 = _T_7220 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8673 = _T_7229 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8682 = _T_7238 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8691 = _T_7247 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8700 = _T_7112 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8709 = _T_7121 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8718 = _T_7130 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8727 = _T_7139 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8736 = _T_7148 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8745 = _T_7157 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8754 = _T_7166 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8763 = _T_7175 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8772 = _T_7184 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8781 = _T_7193 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8790 = _T_7202 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8799 = _T_7211 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8808 = _T_7220 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8817 = _T_7229 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8826 = _T_7238 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8835 = _T_7247 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8844 = _T_7112 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8853 = _T_7121 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8862 = _T_7130 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8871 = _T_7139 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8880 = _T_7148 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8889 = _T_7157 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8898 = _T_7166 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8907 = _T_7175 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8916 = _T_7184 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8925 = _T_7193 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8934 = _T_7202 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8943 = _T_7211 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8952 = _T_7220 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8961 = _T_7229 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8970 = _T_7238 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8979 = _T_7247 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8988 = _T_7112 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_8997 = _T_7121 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9006 = _T_7130 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9015 = _T_7139 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9024 = _T_7148 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9033 = _T_7157 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9042 = _T_7166 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9051 = _T_7175 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9060 = _T_7184 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9069 = _T_7193 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9078 = _T_7202 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9087 = _T_7211 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9096 = _T_7220 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9105 = _T_7229 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9114 = _T_7238 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9123 = _T_7247 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9132 = _T_7112 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9141 = _T_7121 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9150 = _T_7130 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9159 = _T_7139 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9168 = _T_7148 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9177 = _T_7157 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9186 = _T_7166 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9195 = _T_7175 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9204 = _T_7184 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9213 = _T_7193 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9222 = _T_7202 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9231 = _T_7211 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9240 = _T_7220 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9249 = _T_7229 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9258 = _T_7238 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9267 = _T_7247 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9276 = _T_7112 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9285 = _T_7121 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9294 = _T_7130 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9303 = _T_7139 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9312 = _T_7148 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9321 = _T_7157 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9330 = _T_7166 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9339 = _T_7175 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9348 = _T_7184 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9357 = _T_7193 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9366 = _T_7202 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9375 = _T_7211 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9384 = _T_7220 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9393 = _T_7229 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9402 = _T_7238 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9411 = _T_7247 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9416 = bht_wr_en2[1] & _T_7111; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9420 = _T_9416 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9425 = bht_wr_en2[1] & _T_7120; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9429 = _T_9425 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9434 = bht_wr_en2[1] & _T_7129; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9438 = _T_9434 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9443 = bht_wr_en2[1] & _T_7138; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9447 = _T_9443 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9452 = bht_wr_en2[1] & _T_7147; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9456 = _T_9452 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9461 = bht_wr_en2[1] & _T_7156; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9465 = _T_9461 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9470 = bht_wr_en2[1] & _T_7165; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9474 = _T_9470 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9479 = bht_wr_en2[1] & _T_7174; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9483 = _T_9479 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9488 = bht_wr_en2[1] & _T_7183; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9492 = _T_9488 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9497 = bht_wr_en2[1] & _T_7192; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9501 = _T_9497 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9506 = bht_wr_en2[1] & _T_7201; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9510 = _T_9506 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9515 = bht_wr_en2[1] & _T_7210; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9519 = _T_9515 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9524 = bht_wr_en2[1] & _T_7219; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9528 = _T_9524 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9533 = bht_wr_en2[1] & _T_7228; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9537 = _T_9533 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9542 = bht_wr_en2[1] & _T_7237; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9546 = _T_9542 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9551 = bht_wr_en2[1] & _T_7246; // @[ifu_bp_ctl.scala 512:23]
  wire  _T_9555 = _T_9551 & _T_6764; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9564 = _T_9416 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9573 = _T_9425 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9582 = _T_9434 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9591 = _T_9443 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9600 = _T_9452 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9609 = _T_9461 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9618 = _T_9470 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9627 = _T_9479 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9636 = _T_9488 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9645 = _T_9497 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9654 = _T_9506 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9663 = _T_9515 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9672 = _T_9524 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9681 = _T_9533 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9690 = _T_9542 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9699 = _T_9551 & _T_6775; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9708 = _T_9416 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9717 = _T_9425 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9726 = _T_9434 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9735 = _T_9443 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9744 = _T_9452 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9753 = _T_9461 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9762 = _T_9470 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9771 = _T_9479 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9780 = _T_9488 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9789 = _T_9497 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9798 = _T_9506 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9807 = _T_9515 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9816 = _T_9524 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9825 = _T_9533 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9834 = _T_9542 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9843 = _T_9551 & _T_6786; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9852 = _T_9416 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9861 = _T_9425 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9870 = _T_9434 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9879 = _T_9443 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9888 = _T_9452 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9897 = _T_9461 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9906 = _T_9470 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9915 = _T_9479 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9924 = _T_9488 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9933 = _T_9497 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9942 = _T_9506 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9951 = _T_9515 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9960 = _T_9524 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9969 = _T_9533 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9978 = _T_9542 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9987 = _T_9551 & _T_6797; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_9996 = _T_9416 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10005 = _T_9425 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10014 = _T_9434 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10023 = _T_9443 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10032 = _T_9452 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10041 = _T_9461 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10050 = _T_9470 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10059 = _T_9479 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10068 = _T_9488 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10077 = _T_9497 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10086 = _T_9506 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10095 = _T_9515 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10104 = _T_9524 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10113 = _T_9533 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10122 = _T_9542 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10131 = _T_9551 & _T_6808; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10140 = _T_9416 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10149 = _T_9425 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10158 = _T_9434 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10167 = _T_9443 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10176 = _T_9452 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10185 = _T_9461 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10194 = _T_9470 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10203 = _T_9479 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10212 = _T_9488 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10221 = _T_9497 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10230 = _T_9506 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10239 = _T_9515 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10248 = _T_9524 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10257 = _T_9533 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10266 = _T_9542 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10275 = _T_9551 & _T_6819; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10284 = _T_9416 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10293 = _T_9425 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10302 = _T_9434 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10311 = _T_9443 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10320 = _T_9452 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10329 = _T_9461 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10338 = _T_9470 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10347 = _T_9479 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10356 = _T_9488 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10365 = _T_9497 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10374 = _T_9506 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10383 = _T_9515 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10392 = _T_9524 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10401 = _T_9533 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10410 = _T_9542 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10419 = _T_9551 & _T_6830; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10428 = _T_9416 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10437 = _T_9425 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10446 = _T_9434 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10455 = _T_9443 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10464 = _T_9452 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10473 = _T_9461 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10482 = _T_9470 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10491 = _T_9479 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10500 = _T_9488 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10509 = _T_9497 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10518 = _T_9506 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10527 = _T_9515 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10536 = _T_9524 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10545 = _T_9533 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10554 = _T_9542 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10563 = _T_9551 & _T_6841; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10572 = _T_9416 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10581 = _T_9425 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10590 = _T_9434 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10599 = _T_9443 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10608 = _T_9452 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10617 = _T_9461 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10626 = _T_9470 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10635 = _T_9479 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10644 = _T_9488 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10653 = _T_9497 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10662 = _T_9506 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10671 = _T_9515 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10680 = _T_9524 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10689 = _T_9533 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10698 = _T_9542 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10707 = _T_9551 & _T_6852; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10716 = _T_9416 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10725 = _T_9425 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10734 = _T_9434 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10743 = _T_9443 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10752 = _T_9452 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10761 = _T_9461 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10770 = _T_9470 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10779 = _T_9479 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10788 = _T_9488 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10797 = _T_9497 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10806 = _T_9506 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10815 = _T_9515 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10824 = _T_9524 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10833 = _T_9533 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10842 = _T_9542 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10851 = _T_9551 & _T_6863; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10860 = _T_9416 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10869 = _T_9425 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10878 = _T_9434 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10887 = _T_9443 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10896 = _T_9452 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10905 = _T_9461 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10914 = _T_9470 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10923 = _T_9479 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10932 = _T_9488 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10941 = _T_9497 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10950 = _T_9506 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10959 = _T_9515 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10968 = _T_9524 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10977 = _T_9533 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10986 = _T_9542 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_10995 = _T_9551 & _T_6874; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11004 = _T_9416 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11013 = _T_9425 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11022 = _T_9434 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11031 = _T_9443 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11040 = _T_9452 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11049 = _T_9461 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11058 = _T_9470 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11067 = _T_9479 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11076 = _T_9488 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11085 = _T_9497 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11094 = _T_9506 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11103 = _T_9515 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11112 = _T_9524 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11121 = _T_9533 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11130 = _T_9542 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11139 = _T_9551 & _T_6885; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11148 = _T_9416 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11157 = _T_9425 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11166 = _T_9434 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11175 = _T_9443 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11184 = _T_9452 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11193 = _T_9461 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11202 = _T_9470 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11211 = _T_9479 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11220 = _T_9488 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11229 = _T_9497 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11238 = _T_9506 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11247 = _T_9515 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11256 = _T_9524 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11265 = _T_9533 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11274 = _T_9542 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11283 = _T_9551 & _T_6896; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11292 = _T_9416 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11301 = _T_9425 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11310 = _T_9434 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11319 = _T_9443 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11328 = _T_9452 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11337 = _T_9461 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11346 = _T_9470 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11355 = _T_9479 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11364 = _T_9488 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11373 = _T_9497 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11382 = _T_9506 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11391 = _T_9515 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11400 = _T_9524 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11409 = _T_9533 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11418 = _T_9542 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11427 = _T_9551 & _T_6907; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11436 = _T_9416 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11445 = _T_9425 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11454 = _T_9434 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11463 = _T_9443 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11472 = _T_9452 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11481 = _T_9461 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11490 = _T_9470 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11499 = _T_9479 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11508 = _T_9488 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11517 = _T_9497 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11526 = _T_9506 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11535 = _T_9515 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11544 = _T_9524 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11553 = _T_9533 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11562 = _T_9542 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11571 = _T_9551 & _T_6918; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11580 = _T_9416 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11589 = _T_9425 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11598 = _T_9434 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11607 = _T_9443 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11616 = _T_9452 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11625 = _T_9461 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11634 = _T_9470 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11643 = _T_9479 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11652 = _T_9488 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11661 = _T_9497 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11670 = _T_9506 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11679 = _T_9515 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11688 = _T_9524 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11697 = _T_9533 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11706 = _T_9542 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11715 = _T_9551 & _T_6929; // @[ifu_bp_ctl.scala 512:81]
  wire  _T_11719 = mp_hashed[3:0] == 4'h0; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11720 = bht_wr_en0[0] & _T_11719; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11724 = _T_11720 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_0 = _T_11724 | _T_7116; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11736 = mp_hashed[3:0] == 4'h1; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11737 = bht_wr_en0[0] & _T_11736; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11741 = _T_11737 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_1 = _T_11741 | _T_7125; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11753 = mp_hashed[3:0] == 4'h2; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11754 = bht_wr_en0[0] & _T_11753; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11758 = _T_11754 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_2 = _T_11758 | _T_7134; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11770 = mp_hashed[3:0] == 4'h3; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11771 = bht_wr_en0[0] & _T_11770; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11775 = _T_11771 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_3 = _T_11775 | _T_7143; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11787 = mp_hashed[3:0] == 4'h4; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11788 = bht_wr_en0[0] & _T_11787; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11792 = _T_11788 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_4 = _T_11792 | _T_7152; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11804 = mp_hashed[3:0] == 4'h5; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11805 = bht_wr_en0[0] & _T_11804; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11809 = _T_11805 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_5 = _T_11809 | _T_7161; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11821 = mp_hashed[3:0] == 4'h6; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11822 = bht_wr_en0[0] & _T_11821; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11826 = _T_11822 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_6 = _T_11826 | _T_7170; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11838 = mp_hashed[3:0] == 4'h7; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11839 = bht_wr_en0[0] & _T_11838; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11843 = _T_11839 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_7 = _T_11843 | _T_7179; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11855 = mp_hashed[3:0] == 4'h8; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11856 = bht_wr_en0[0] & _T_11855; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11860 = _T_11856 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_8 = _T_11860 | _T_7188; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11872 = mp_hashed[3:0] == 4'h9; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11873 = bht_wr_en0[0] & _T_11872; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11877 = _T_11873 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_9 = _T_11877 | _T_7197; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11889 = mp_hashed[3:0] == 4'ha; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11890 = bht_wr_en0[0] & _T_11889; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11894 = _T_11890 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_10 = _T_11894 | _T_7206; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11906 = mp_hashed[3:0] == 4'hb; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11907 = bht_wr_en0[0] & _T_11906; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11911 = _T_11907 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_11 = _T_11911 | _T_7215; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11923 = mp_hashed[3:0] == 4'hc; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11924 = bht_wr_en0[0] & _T_11923; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11928 = _T_11924 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_12 = _T_11928 | _T_7224; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11940 = mp_hashed[3:0] == 4'hd; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11941 = bht_wr_en0[0] & _T_11940; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11945 = _T_11941 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_13 = _T_11945 | _T_7233; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11957 = mp_hashed[3:0] == 4'he; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11958 = bht_wr_en0[0] & _T_11957; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11962 = _T_11958 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_14 = _T_11962 | _T_7242; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11974 = mp_hashed[3:0] == 4'hf; // @[ifu_bp_ctl.scala 521:97]
  wire  _T_11975 = bht_wr_en0[0] & _T_11974; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_11979 = _T_11975 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_0_15 = _T_11979 | _T_7251; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_11996 = _T_11720 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_0 = _T_11996 | _T_7260; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12013 = _T_11737 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_1 = _T_12013 | _T_7269; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12030 = _T_11754 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_2 = _T_12030 | _T_7278; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12047 = _T_11771 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_3 = _T_12047 | _T_7287; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12064 = _T_11788 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_4 = _T_12064 | _T_7296; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12081 = _T_11805 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_5 = _T_12081 | _T_7305; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12098 = _T_11822 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_6 = _T_12098 | _T_7314; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12115 = _T_11839 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_7 = _T_12115 | _T_7323; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12132 = _T_11856 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_8 = _T_12132 | _T_7332; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12149 = _T_11873 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_9 = _T_12149 | _T_7341; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12166 = _T_11890 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_10 = _T_12166 | _T_7350; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12183 = _T_11907 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_11 = _T_12183 | _T_7359; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12200 = _T_11924 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_12 = _T_12200 | _T_7368; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12217 = _T_11941 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_13 = _T_12217 | _T_7377; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12234 = _T_11958 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_14 = _T_12234 | _T_7386; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12251 = _T_11975 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_1_15 = _T_12251 | _T_7395; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12268 = _T_11720 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_0 = _T_12268 | _T_7404; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12285 = _T_11737 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_1 = _T_12285 | _T_7413; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12302 = _T_11754 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_2 = _T_12302 | _T_7422; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12319 = _T_11771 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_3 = _T_12319 | _T_7431; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12336 = _T_11788 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_4 = _T_12336 | _T_7440; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12353 = _T_11805 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_5 = _T_12353 | _T_7449; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12370 = _T_11822 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_6 = _T_12370 | _T_7458; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12387 = _T_11839 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_7 = _T_12387 | _T_7467; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12404 = _T_11856 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_8 = _T_12404 | _T_7476; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12421 = _T_11873 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_9 = _T_12421 | _T_7485; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12438 = _T_11890 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_10 = _T_12438 | _T_7494; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12455 = _T_11907 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_11 = _T_12455 | _T_7503; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12472 = _T_11924 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_12 = _T_12472 | _T_7512; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12489 = _T_11941 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_13 = _T_12489 | _T_7521; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12506 = _T_11958 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_14 = _T_12506 | _T_7530; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12523 = _T_11975 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_2_15 = _T_12523 | _T_7539; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12540 = _T_11720 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_0 = _T_12540 | _T_7548; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12557 = _T_11737 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_1 = _T_12557 | _T_7557; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12574 = _T_11754 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_2 = _T_12574 | _T_7566; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12591 = _T_11771 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_3 = _T_12591 | _T_7575; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12608 = _T_11788 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_4 = _T_12608 | _T_7584; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12625 = _T_11805 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_5 = _T_12625 | _T_7593; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12642 = _T_11822 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_6 = _T_12642 | _T_7602; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12659 = _T_11839 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_7 = _T_12659 | _T_7611; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12676 = _T_11856 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_8 = _T_12676 | _T_7620; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12693 = _T_11873 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_9 = _T_12693 | _T_7629; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12710 = _T_11890 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_10 = _T_12710 | _T_7638; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12727 = _T_11907 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_11 = _T_12727 | _T_7647; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12744 = _T_11924 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_12 = _T_12744 | _T_7656; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12761 = _T_11941 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_13 = _T_12761 | _T_7665; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12778 = _T_11958 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_14 = _T_12778 | _T_7674; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12795 = _T_11975 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_3_15 = _T_12795 | _T_7683; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12812 = _T_11720 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_0 = _T_12812 | _T_7692; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12829 = _T_11737 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_1 = _T_12829 | _T_7701; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12846 = _T_11754 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_2 = _T_12846 | _T_7710; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12863 = _T_11771 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_3 = _T_12863 | _T_7719; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12880 = _T_11788 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_4 = _T_12880 | _T_7728; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12897 = _T_11805 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_5 = _T_12897 | _T_7737; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12914 = _T_11822 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_6 = _T_12914 | _T_7746; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12931 = _T_11839 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_7 = _T_12931 | _T_7755; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12948 = _T_11856 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_8 = _T_12948 | _T_7764; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12965 = _T_11873 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_9 = _T_12965 | _T_7773; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12982 = _T_11890 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_10 = _T_12982 | _T_7782; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_12999 = _T_11907 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_11 = _T_12999 | _T_7791; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13016 = _T_11924 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_12 = _T_13016 | _T_7800; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13033 = _T_11941 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_13 = _T_13033 | _T_7809; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13050 = _T_11958 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_14 = _T_13050 | _T_7818; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13067 = _T_11975 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_4_15 = _T_13067 | _T_7827; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13084 = _T_11720 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_0 = _T_13084 | _T_7836; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13101 = _T_11737 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_1 = _T_13101 | _T_7845; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13118 = _T_11754 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_2 = _T_13118 | _T_7854; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13135 = _T_11771 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_3 = _T_13135 | _T_7863; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13152 = _T_11788 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_4 = _T_13152 | _T_7872; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13169 = _T_11805 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_5 = _T_13169 | _T_7881; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13186 = _T_11822 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_6 = _T_13186 | _T_7890; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13203 = _T_11839 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_7 = _T_13203 | _T_7899; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13220 = _T_11856 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_8 = _T_13220 | _T_7908; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13237 = _T_11873 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_9 = _T_13237 | _T_7917; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13254 = _T_11890 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_10 = _T_13254 | _T_7926; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13271 = _T_11907 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_11 = _T_13271 | _T_7935; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13288 = _T_11924 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_12 = _T_13288 | _T_7944; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13305 = _T_11941 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_13 = _T_13305 | _T_7953; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13322 = _T_11958 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_14 = _T_13322 | _T_7962; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13339 = _T_11975 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_5_15 = _T_13339 | _T_7971; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13356 = _T_11720 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_0 = _T_13356 | _T_7980; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13373 = _T_11737 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_1 = _T_13373 | _T_7989; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13390 = _T_11754 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_2 = _T_13390 | _T_7998; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13407 = _T_11771 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_3 = _T_13407 | _T_8007; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13424 = _T_11788 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_4 = _T_13424 | _T_8016; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13441 = _T_11805 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_5 = _T_13441 | _T_8025; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13458 = _T_11822 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_6 = _T_13458 | _T_8034; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13475 = _T_11839 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_7 = _T_13475 | _T_8043; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13492 = _T_11856 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_8 = _T_13492 | _T_8052; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13509 = _T_11873 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_9 = _T_13509 | _T_8061; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13526 = _T_11890 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_10 = _T_13526 | _T_8070; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13543 = _T_11907 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_11 = _T_13543 | _T_8079; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13560 = _T_11924 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_12 = _T_13560 | _T_8088; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13577 = _T_11941 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_13 = _T_13577 | _T_8097; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13594 = _T_11958 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_14 = _T_13594 | _T_8106; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13611 = _T_11975 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_6_15 = _T_13611 | _T_8115; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13628 = _T_11720 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_0 = _T_13628 | _T_8124; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13645 = _T_11737 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_1 = _T_13645 | _T_8133; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13662 = _T_11754 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_2 = _T_13662 | _T_8142; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13679 = _T_11771 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_3 = _T_13679 | _T_8151; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13696 = _T_11788 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_4 = _T_13696 | _T_8160; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13713 = _T_11805 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_5 = _T_13713 | _T_8169; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13730 = _T_11822 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_6 = _T_13730 | _T_8178; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13747 = _T_11839 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_7 = _T_13747 | _T_8187; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13764 = _T_11856 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_8 = _T_13764 | _T_8196; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13781 = _T_11873 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_9 = _T_13781 | _T_8205; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13798 = _T_11890 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_10 = _T_13798 | _T_8214; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13815 = _T_11907 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_11 = _T_13815 | _T_8223; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13832 = _T_11924 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_12 = _T_13832 | _T_8232; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13849 = _T_11941 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_13 = _T_13849 | _T_8241; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13866 = _T_11958 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_14 = _T_13866 | _T_8250; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13883 = _T_11975 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_7_15 = _T_13883 | _T_8259; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13900 = _T_11720 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_0 = _T_13900 | _T_8268; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13917 = _T_11737 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_1 = _T_13917 | _T_8277; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13934 = _T_11754 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_2 = _T_13934 | _T_8286; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13951 = _T_11771 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_3 = _T_13951 | _T_8295; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13968 = _T_11788 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_4 = _T_13968 | _T_8304; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_13985 = _T_11805 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_5 = _T_13985 | _T_8313; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14002 = _T_11822 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_6 = _T_14002 | _T_8322; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14019 = _T_11839 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_7 = _T_14019 | _T_8331; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14036 = _T_11856 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_8 = _T_14036 | _T_8340; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14053 = _T_11873 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_9 = _T_14053 | _T_8349; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14070 = _T_11890 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_10 = _T_14070 | _T_8358; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14087 = _T_11907 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_11 = _T_14087 | _T_8367; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14104 = _T_11924 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_12 = _T_14104 | _T_8376; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14121 = _T_11941 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_13 = _T_14121 | _T_8385; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14138 = _T_11958 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_14 = _T_14138 | _T_8394; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14155 = _T_11975 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_8_15 = _T_14155 | _T_8403; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14172 = _T_11720 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_0 = _T_14172 | _T_8412; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14189 = _T_11737 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_1 = _T_14189 | _T_8421; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14206 = _T_11754 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_2 = _T_14206 | _T_8430; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14223 = _T_11771 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_3 = _T_14223 | _T_8439; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14240 = _T_11788 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_4 = _T_14240 | _T_8448; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14257 = _T_11805 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_5 = _T_14257 | _T_8457; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14274 = _T_11822 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_6 = _T_14274 | _T_8466; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14291 = _T_11839 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_7 = _T_14291 | _T_8475; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14308 = _T_11856 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_8 = _T_14308 | _T_8484; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14325 = _T_11873 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_9 = _T_14325 | _T_8493; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14342 = _T_11890 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_10 = _T_14342 | _T_8502; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14359 = _T_11907 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_11 = _T_14359 | _T_8511; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14376 = _T_11924 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_12 = _T_14376 | _T_8520; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14393 = _T_11941 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_13 = _T_14393 | _T_8529; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14410 = _T_11958 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_14 = _T_14410 | _T_8538; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14427 = _T_11975 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_9_15 = _T_14427 | _T_8547; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14444 = _T_11720 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_0 = _T_14444 | _T_8556; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14461 = _T_11737 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_1 = _T_14461 | _T_8565; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14478 = _T_11754 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_2 = _T_14478 | _T_8574; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14495 = _T_11771 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_3 = _T_14495 | _T_8583; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14512 = _T_11788 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_4 = _T_14512 | _T_8592; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14529 = _T_11805 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_5 = _T_14529 | _T_8601; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14546 = _T_11822 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_6 = _T_14546 | _T_8610; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14563 = _T_11839 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_7 = _T_14563 | _T_8619; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14580 = _T_11856 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_8 = _T_14580 | _T_8628; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14597 = _T_11873 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_9 = _T_14597 | _T_8637; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14614 = _T_11890 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_10 = _T_14614 | _T_8646; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14631 = _T_11907 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_11 = _T_14631 | _T_8655; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14648 = _T_11924 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_12 = _T_14648 | _T_8664; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14665 = _T_11941 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_13 = _T_14665 | _T_8673; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14682 = _T_11958 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_14 = _T_14682 | _T_8682; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14699 = _T_11975 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_10_15 = _T_14699 | _T_8691; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14716 = _T_11720 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_0 = _T_14716 | _T_8700; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14733 = _T_11737 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_1 = _T_14733 | _T_8709; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14750 = _T_11754 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_2 = _T_14750 | _T_8718; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14767 = _T_11771 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_3 = _T_14767 | _T_8727; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14784 = _T_11788 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_4 = _T_14784 | _T_8736; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14801 = _T_11805 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_5 = _T_14801 | _T_8745; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14818 = _T_11822 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_6 = _T_14818 | _T_8754; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14835 = _T_11839 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_7 = _T_14835 | _T_8763; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14852 = _T_11856 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_8 = _T_14852 | _T_8772; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14869 = _T_11873 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_9 = _T_14869 | _T_8781; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14886 = _T_11890 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_10 = _T_14886 | _T_8790; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14903 = _T_11907 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_11 = _T_14903 | _T_8799; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14920 = _T_11924 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_12 = _T_14920 | _T_8808; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14937 = _T_11941 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_13 = _T_14937 | _T_8817; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14954 = _T_11958 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_14 = _T_14954 | _T_8826; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14971 = _T_11975 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_11_15 = _T_14971 | _T_8835; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_14988 = _T_11720 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_0 = _T_14988 | _T_8844; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15005 = _T_11737 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_1 = _T_15005 | _T_8853; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15022 = _T_11754 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_2 = _T_15022 | _T_8862; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15039 = _T_11771 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_3 = _T_15039 | _T_8871; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15056 = _T_11788 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_4 = _T_15056 | _T_8880; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15073 = _T_11805 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_5 = _T_15073 | _T_8889; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15090 = _T_11822 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_6 = _T_15090 | _T_8898; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15107 = _T_11839 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_7 = _T_15107 | _T_8907; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15124 = _T_11856 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_8 = _T_15124 | _T_8916; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15141 = _T_11873 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_9 = _T_15141 | _T_8925; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15158 = _T_11890 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_10 = _T_15158 | _T_8934; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15175 = _T_11907 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_11 = _T_15175 | _T_8943; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15192 = _T_11924 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_12 = _T_15192 | _T_8952; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15209 = _T_11941 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_13 = _T_15209 | _T_8961; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15226 = _T_11958 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_14 = _T_15226 | _T_8970; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15243 = _T_11975 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_12_15 = _T_15243 | _T_8979; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15260 = _T_11720 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_0 = _T_15260 | _T_8988; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15277 = _T_11737 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_1 = _T_15277 | _T_8997; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15294 = _T_11754 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_2 = _T_15294 | _T_9006; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15311 = _T_11771 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_3 = _T_15311 | _T_9015; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15328 = _T_11788 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_4 = _T_15328 | _T_9024; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15345 = _T_11805 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_5 = _T_15345 | _T_9033; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15362 = _T_11822 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_6 = _T_15362 | _T_9042; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15379 = _T_11839 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_7 = _T_15379 | _T_9051; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15396 = _T_11856 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_8 = _T_15396 | _T_9060; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15413 = _T_11873 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_9 = _T_15413 | _T_9069; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15430 = _T_11890 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_10 = _T_15430 | _T_9078; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15447 = _T_11907 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_11 = _T_15447 | _T_9087; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15464 = _T_11924 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_12 = _T_15464 | _T_9096; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15481 = _T_11941 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_13 = _T_15481 | _T_9105; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15498 = _T_11958 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_14 = _T_15498 | _T_9114; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15515 = _T_11975 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_13_15 = _T_15515 | _T_9123; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15532 = _T_11720 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_0 = _T_15532 | _T_9132; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15549 = _T_11737 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_1 = _T_15549 | _T_9141; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15566 = _T_11754 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_2 = _T_15566 | _T_9150; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15583 = _T_11771 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_3 = _T_15583 | _T_9159; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15600 = _T_11788 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_4 = _T_15600 | _T_9168; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15617 = _T_11805 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_5 = _T_15617 | _T_9177; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15634 = _T_11822 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_6 = _T_15634 | _T_9186; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15651 = _T_11839 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_7 = _T_15651 | _T_9195; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15668 = _T_11856 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_8 = _T_15668 | _T_9204; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15685 = _T_11873 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_9 = _T_15685 | _T_9213; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15702 = _T_11890 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_10 = _T_15702 | _T_9222; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15719 = _T_11907 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_11 = _T_15719 | _T_9231; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15736 = _T_11924 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_12 = _T_15736 | _T_9240; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15753 = _T_11941 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_13 = _T_15753 | _T_9249; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15770 = _T_11958 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_14 = _T_15770 | _T_9258; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15787 = _T_11975 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_14_15 = _T_15787 | _T_9267; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15804 = _T_11720 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_0 = _T_15804 | _T_9276; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15821 = _T_11737 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_1 = _T_15821 | _T_9285; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15838 = _T_11754 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_2 = _T_15838 | _T_9294; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15855 = _T_11771 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_3 = _T_15855 | _T_9303; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15872 = _T_11788 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_4 = _T_15872 | _T_9312; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15889 = _T_11805 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_5 = _T_15889 | _T_9321; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15906 = _T_11822 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_6 = _T_15906 | _T_9330; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15923 = _T_11839 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_7 = _T_15923 | _T_9339; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15940 = _T_11856 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_8 = _T_15940 | _T_9348; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15957 = _T_11873 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_9 = _T_15957 | _T_9357; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15974 = _T_11890 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_10 = _T_15974 | _T_9366; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_15991 = _T_11907 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_11 = _T_15991 | _T_9375; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16008 = _T_11924 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_12 = _T_16008 | _T_9384; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16025 = _T_11941 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_13 = _T_16025 | _T_9393; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16042 = _T_11958 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_14 = _T_16042 | _T_9402; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16059 = _T_11975 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_0_15_15 = _T_16059 | _T_9411; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16072 = bht_wr_en0[1] & _T_11719; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16076 = _T_16072 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_0 = _T_16076 | _T_9420; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16089 = bht_wr_en0[1] & _T_11736; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16093 = _T_16089 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_1 = _T_16093 | _T_9429; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16106 = bht_wr_en0[1] & _T_11753; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16110 = _T_16106 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_2 = _T_16110 | _T_9438; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16123 = bht_wr_en0[1] & _T_11770; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16127 = _T_16123 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_3 = _T_16127 | _T_9447; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16140 = bht_wr_en0[1] & _T_11787; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16144 = _T_16140 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_4 = _T_16144 | _T_9456; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16157 = bht_wr_en0[1] & _T_11804; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16161 = _T_16157 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_5 = _T_16161 | _T_9465; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16174 = bht_wr_en0[1] & _T_11821; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16178 = _T_16174 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_6 = _T_16178 | _T_9474; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16191 = bht_wr_en0[1] & _T_11838; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16195 = _T_16191 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_7 = _T_16195 | _T_9483; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16208 = bht_wr_en0[1] & _T_11855; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16212 = _T_16208 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_8 = _T_16212 | _T_9492; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16225 = bht_wr_en0[1] & _T_11872; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16229 = _T_16225 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_9 = _T_16229 | _T_9501; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16242 = bht_wr_en0[1] & _T_11889; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16246 = _T_16242 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_10 = _T_16246 | _T_9510; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16259 = bht_wr_en0[1] & _T_11906; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16263 = _T_16259 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_11 = _T_16263 | _T_9519; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16276 = bht_wr_en0[1] & _T_11923; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16280 = _T_16276 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_12 = _T_16280 | _T_9528; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16293 = bht_wr_en0[1] & _T_11940; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16297 = _T_16293 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_13 = _T_16297 | _T_9537; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16310 = bht_wr_en0[1] & _T_11957; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16314 = _T_16310 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_14 = _T_16314 | _T_9546; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16327 = bht_wr_en0[1] & _T_11974; // @[ifu_bp_ctl.scala 521:45]
  wire  _T_16331 = _T_16327 & _T_6759; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_0_15 = _T_16331 | _T_9555; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16348 = _T_16072 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_0 = _T_16348 | _T_9564; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16365 = _T_16089 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_1 = _T_16365 | _T_9573; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16382 = _T_16106 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_2 = _T_16382 | _T_9582; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16399 = _T_16123 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_3 = _T_16399 | _T_9591; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16416 = _T_16140 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_4 = _T_16416 | _T_9600; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16433 = _T_16157 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_5 = _T_16433 | _T_9609; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16450 = _T_16174 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_6 = _T_16450 | _T_9618; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16467 = _T_16191 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_7 = _T_16467 | _T_9627; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16484 = _T_16208 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_8 = _T_16484 | _T_9636; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16501 = _T_16225 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_9 = _T_16501 | _T_9645; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16518 = _T_16242 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_10 = _T_16518 | _T_9654; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16535 = _T_16259 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_11 = _T_16535 | _T_9663; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16552 = _T_16276 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_12 = _T_16552 | _T_9672; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16569 = _T_16293 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_13 = _T_16569 | _T_9681; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16586 = _T_16310 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_14 = _T_16586 | _T_9690; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16603 = _T_16327 & _T_6770; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_1_15 = _T_16603 | _T_9699; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16620 = _T_16072 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_0 = _T_16620 | _T_9708; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16637 = _T_16089 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_1 = _T_16637 | _T_9717; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16654 = _T_16106 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_2 = _T_16654 | _T_9726; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16671 = _T_16123 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_3 = _T_16671 | _T_9735; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16688 = _T_16140 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_4 = _T_16688 | _T_9744; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16705 = _T_16157 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_5 = _T_16705 | _T_9753; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16722 = _T_16174 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_6 = _T_16722 | _T_9762; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16739 = _T_16191 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_7 = _T_16739 | _T_9771; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16756 = _T_16208 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_8 = _T_16756 | _T_9780; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16773 = _T_16225 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_9 = _T_16773 | _T_9789; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16790 = _T_16242 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_10 = _T_16790 | _T_9798; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16807 = _T_16259 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_11 = _T_16807 | _T_9807; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16824 = _T_16276 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_12 = _T_16824 | _T_9816; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16841 = _T_16293 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_13 = _T_16841 | _T_9825; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16858 = _T_16310 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_14 = _T_16858 | _T_9834; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16875 = _T_16327 & _T_6781; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_2_15 = _T_16875 | _T_9843; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16892 = _T_16072 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_0 = _T_16892 | _T_9852; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16909 = _T_16089 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_1 = _T_16909 | _T_9861; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16926 = _T_16106 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_2 = _T_16926 | _T_9870; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16943 = _T_16123 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_3 = _T_16943 | _T_9879; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16960 = _T_16140 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_4 = _T_16960 | _T_9888; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16977 = _T_16157 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_5 = _T_16977 | _T_9897; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_16994 = _T_16174 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_6 = _T_16994 | _T_9906; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17011 = _T_16191 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_7 = _T_17011 | _T_9915; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17028 = _T_16208 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_8 = _T_17028 | _T_9924; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17045 = _T_16225 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_9 = _T_17045 | _T_9933; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17062 = _T_16242 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_10 = _T_17062 | _T_9942; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17079 = _T_16259 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_11 = _T_17079 | _T_9951; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17096 = _T_16276 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_12 = _T_17096 | _T_9960; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17113 = _T_16293 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_13 = _T_17113 | _T_9969; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17130 = _T_16310 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_14 = _T_17130 | _T_9978; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17147 = _T_16327 & _T_6792; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_3_15 = _T_17147 | _T_9987; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17164 = _T_16072 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_0 = _T_17164 | _T_9996; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17181 = _T_16089 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_1 = _T_17181 | _T_10005; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17198 = _T_16106 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_2 = _T_17198 | _T_10014; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17215 = _T_16123 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_3 = _T_17215 | _T_10023; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17232 = _T_16140 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_4 = _T_17232 | _T_10032; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17249 = _T_16157 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_5 = _T_17249 | _T_10041; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17266 = _T_16174 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_6 = _T_17266 | _T_10050; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17283 = _T_16191 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_7 = _T_17283 | _T_10059; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17300 = _T_16208 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_8 = _T_17300 | _T_10068; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17317 = _T_16225 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_9 = _T_17317 | _T_10077; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17334 = _T_16242 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_10 = _T_17334 | _T_10086; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17351 = _T_16259 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_11 = _T_17351 | _T_10095; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17368 = _T_16276 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_12 = _T_17368 | _T_10104; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17385 = _T_16293 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_13 = _T_17385 | _T_10113; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17402 = _T_16310 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_14 = _T_17402 | _T_10122; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17419 = _T_16327 & _T_6803; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_4_15 = _T_17419 | _T_10131; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17436 = _T_16072 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_0 = _T_17436 | _T_10140; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17453 = _T_16089 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_1 = _T_17453 | _T_10149; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17470 = _T_16106 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_2 = _T_17470 | _T_10158; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17487 = _T_16123 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_3 = _T_17487 | _T_10167; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17504 = _T_16140 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_4 = _T_17504 | _T_10176; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17521 = _T_16157 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_5 = _T_17521 | _T_10185; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17538 = _T_16174 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_6 = _T_17538 | _T_10194; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17555 = _T_16191 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_7 = _T_17555 | _T_10203; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17572 = _T_16208 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_8 = _T_17572 | _T_10212; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17589 = _T_16225 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_9 = _T_17589 | _T_10221; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17606 = _T_16242 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_10 = _T_17606 | _T_10230; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17623 = _T_16259 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_11 = _T_17623 | _T_10239; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17640 = _T_16276 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_12 = _T_17640 | _T_10248; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17657 = _T_16293 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_13 = _T_17657 | _T_10257; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17674 = _T_16310 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_14 = _T_17674 | _T_10266; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17691 = _T_16327 & _T_6814; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_5_15 = _T_17691 | _T_10275; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17708 = _T_16072 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_0 = _T_17708 | _T_10284; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17725 = _T_16089 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_1 = _T_17725 | _T_10293; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17742 = _T_16106 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_2 = _T_17742 | _T_10302; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17759 = _T_16123 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_3 = _T_17759 | _T_10311; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17776 = _T_16140 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_4 = _T_17776 | _T_10320; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17793 = _T_16157 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_5 = _T_17793 | _T_10329; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17810 = _T_16174 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_6 = _T_17810 | _T_10338; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17827 = _T_16191 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_7 = _T_17827 | _T_10347; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17844 = _T_16208 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_8 = _T_17844 | _T_10356; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17861 = _T_16225 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_9 = _T_17861 | _T_10365; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17878 = _T_16242 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_10 = _T_17878 | _T_10374; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17895 = _T_16259 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_11 = _T_17895 | _T_10383; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17912 = _T_16276 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_12 = _T_17912 | _T_10392; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17929 = _T_16293 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_13 = _T_17929 | _T_10401; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17946 = _T_16310 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_14 = _T_17946 | _T_10410; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17963 = _T_16327 & _T_6825; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_6_15 = _T_17963 | _T_10419; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17980 = _T_16072 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_0 = _T_17980 | _T_10428; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_17997 = _T_16089 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_1 = _T_17997 | _T_10437; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18014 = _T_16106 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_2 = _T_18014 | _T_10446; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18031 = _T_16123 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_3 = _T_18031 | _T_10455; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18048 = _T_16140 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_4 = _T_18048 | _T_10464; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18065 = _T_16157 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_5 = _T_18065 | _T_10473; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18082 = _T_16174 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_6 = _T_18082 | _T_10482; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18099 = _T_16191 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_7 = _T_18099 | _T_10491; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18116 = _T_16208 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_8 = _T_18116 | _T_10500; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18133 = _T_16225 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_9 = _T_18133 | _T_10509; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18150 = _T_16242 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_10 = _T_18150 | _T_10518; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18167 = _T_16259 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_11 = _T_18167 | _T_10527; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18184 = _T_16276 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_12 = _T_18184 | _T_10536; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18201 = _T_16293 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_13 = _T_18201 | _T_10545; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18218 = _T_16310 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_14 = _T_18218 | _T_10554; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18235 = _T_16327 & _T_6836; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_7_15 = _T_18235 | _T_10563; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18252 = _T_16072 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_0 = _T_18252 | _T_10572; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18269 = _T_16089 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_1 = _T_18269 | _T_10581; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18286 = _T_16106 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_2 = _T_18286 | _T_10590; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18303 = _T_16123 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_3 = _T_18303 | _T_10599; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18320 = _T_16140 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_4 = _T_18320 | _T_10608; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18337 = _T_16157 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_5 = _T_18337 | _T_10617; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18354 = _T_16174 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_6 = _T_18354 | _T_10626; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18371 = _T_16191 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_7 = _T_18371 | _T_10635; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18388 = _T_16208 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_8 = _T_18388 | _T_10644; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18405 = _T_16225 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_9 = _T_18405 | _T_10653; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18422 = _T_16242 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_10 = _T_18422 | _T_10662; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18439 = _T_16259 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_11 = _T_18439 | _T_10671; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18456 = _T_16276 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_12 = _T_18456 | _T_10680; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18473 = _T_16293 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_13 = _T_18473 | _T_10689; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18490 = _T_16310 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_14 = _T_18490 | _T_10698; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18507 = _T_16327 & _T_6847; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_8_15 = _T_18507 | _T_10707; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18524 = _T_16072 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_0 = _T_18524 | _T_10716; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18541 = _T_16089 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_1 = _T_18541 | _T_10725; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18558 = _T_16106 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_2 = _T_18558 | _T_10734; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18575 = _T_16123 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_3 = _T_18575 | _T_10743; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18592 = _T_16140 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_4 = _T_18592 | _T_10752; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18609 = _T_16157 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_5 = _T_18609 | _T_10761; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18626 = _T_16174 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_6 = _T_18626 | _T_10770; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18643 = _T_16191 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_7 = _T_18643 | _T_10779; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18660 = _T_16208 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_8 = _T_18660 | _T_10788; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18677 = _T_16225 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_9 = _T_18677 | _T_10797; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18694 = _T_16242 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_10 = _T_18694 | _T_10806; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18711 = _T_16259 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_11 = _T_18711 | _T_10815; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18728 = _T_16276 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_12 = _T_18728 | _T_10824; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18745 = _T_16293 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_13 = _T_18745 | _T_10833; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18762 = _T_16310 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_14 = _T_18762 | _T_10842; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18779 = _T_16327 & _T_6858; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_9_15 = _T_18779 | _T_10851; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18796 = _T_16072 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_0 = _T_18796 | _T_10860; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18813 = _T_16089 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_1 = _T_18813 | _T_10869; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18830 = _T_16106 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_2 = _T_18830 | _T_10878; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18847 = _T_16123 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_3 = _T_18847 | _T_10887; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18864 = _T_16140 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_4 = _T_18864 | _T_10896; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18881 = _T_16157 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_5 = _T_18881 | _T_10905; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18898 = _T_16174 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_6 = _T_18898 | _T_10914; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18915 = _T_16191 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_7 = _T_18915 | _T_10923; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18932 = _T_16208 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_8 = _T_18932 | _T_10932; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18949 = _T_16225 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_9 = _T_18949 | _T_10941; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18966 = _T_16242 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_10 = _T_18966 | _T_10950; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_18983 = _T_16259 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_11 = _T_18983 | _T_10959; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19000 = _T_16276 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_12 = _T_19000 | _T_10968; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19017 = _T_16293 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_13 = _T_19017 | _T_10977; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19034 = _T_16310 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_14 = _T_19034 | _T_10986; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19051 = _T_16327 & _T_6869; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_10_15 = _T_19051 | _T_10995; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19068 = _T_16072 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_0 = _T_19068 | _T_11004; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19085 = _T_16089 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_1 = _T_19085 | _T_11013; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19102 = _T_16106 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_2 = _T_19102 | _T_11022; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19119 = _T_16123 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_3 = _T_19119 | _T_11031; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19136 = _T_16140 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_4 = _T_19136 | _T_11040; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19153 = _T_16157 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_5 = _T_19153 | _T_11049; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19170 = _T_16174 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_6 = _T_19170 | _T_11058; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19187 = _T_16191 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_7 = _T_19187 | _T_11067; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19204 = _T_16208 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_8 = _T_19204 | _T_11076; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19221 = _T_16225 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_9 = _T_19221 | _T_11085; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19238 = _T_16242 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_10 = _T_19238 | _T_11094; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19255 = _T_16259 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_11 = _T_19255 | _T_11103; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19272 = _T_16276 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_12 = _T_19272 | _T_11112; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19289 = _T_16293 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_13 = _T_19289 | _T_11121; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19306 = _T_16310 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_14 = _T_19306 | _T_11130; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19323 = _T_16327 & _T_6880; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_11_15 = _T_19323 | _T_11139; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19340 = _T_16072 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_0 = _T_19340 | _T_11148; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19357 = _T_16089 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_1 = _T_19357 | _T_11157; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19374 = _T_16106 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_2 = _T_19374 | _T_11166; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19391 = _T_16123 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_3 = _T_19391 | _T_11175; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19408 = _T_16140 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_4 = _T_19408 | _T_11184; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19425 = _T_16157 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_5 = _T_19425 | _T_11193; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19442 = _T_16174 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_6 = _T_19442 | _T_11202; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19459 = _T_16191 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_7 = _T_19459 | _T_11211; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19476 = _T_16208 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_8 = _T_19476 | _T_11220; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19493 = _T_16225 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_9 = _T_19493 | _T_11229; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19510 = _T_16242 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_10 = _T_19510 | _T_11238; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19527 = _T_16259 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_11 = _T_19527 | _T_11247; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19544 = _T_16276 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_12 = _T_19544 | _T_11256; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19561 = _T_16293 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_13 = _T_19561 | _T_11265; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19578 = _T_16310 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_14 = _T_19578 | _T_11274; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19595 = _T_16327 & _T_6891; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_12_15 = _T_19595 | _T_11283; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19612 = _T_16072 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_0 = _T_19612 | _T_11292; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19629 = _T_16089 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_1 = _T_19629 | _T_11301; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19646 = _T_16106 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_2 = _T_19646 | _T_11310; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19663 = _T_16123 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_3 = _T_19663 | _T_11319; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19680 = _T_16140 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_4 = _T_19680 | _T_11328; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19697 = _T_16157 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_5 = _T_19697 | _T_11337; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19714 = _T_16174 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_6 = _T_19714 | _T_11346; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19731 = _T_16191 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_7 = _T_19731 | _T_11355; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19748 = _T_16208 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_8 = _T_19748 | _T_11364; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19765 = _T_16225 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_9 = _T_19765 | _T_11373; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19782 = _T_16242 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_10 = _T_19782 | _T_11382; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19799 = _T_16259 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_11 = _T_19799 | _T_11391; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19816 = _T_16276 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_12 = _T_19816 | _T_11400; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19833 = _T_16293 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_13 = _T_19833 | _T_11409; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19850 = _T_16310 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_14 = _T_19850 | _T_11418; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19867 = _T_16327 & _T_6902; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_13_15 = _T_19867 | _T_11427; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19884 = _T_16072 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_0 = _T_19884 | _T_11436; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19901 = _T_16089 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_1 = _T_19901 | _T_11445; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19918 = _T_16106 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_2 = _T_19918 | _T_11454; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19935 = _T_16123 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_3 = _T_19935 | _T_11463; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19952 = _T_16140 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_4 = _T_19952 | _T_11472; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19969 = _T_16157 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_5 = _T_19969 | _T_11481; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_19986 = _T_16174 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_6 = _T_19986 | _T_11490; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20003 = _T_16191 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_7 = _T_20003 | _T_11499; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20020 = _T_16208 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_8 = _T_20020 | _T_11508; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20037 = _T_16225 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_9 = _T_20037 | _T_11517; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20054 = _T_16242 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_10 = _T_20054 | _T_11526; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20071 = _T_16259 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_11 = _T_20071 | _T_11535; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20088 = _T_16276 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_12 = _T_20088 | _T_11544; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20105 = _T_16293 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_13 = _T_20105 | _T_11553; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20122 = _T_16310 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_14 = _T_20122 | _T_11562; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20139 = _T_16327 & _T_6913; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_14_15 = _T_20139 | _T_11571; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20156 = _T_16072 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_0 = _T_20156 | _T_11580; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20173 = _T_16089 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_1 = _T_20173 | _T_11589; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20190 = _T_16106 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_2 = _T_20190 | _T_11598; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20207 = _T_16123 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_3 = _T_20207 | _T_11607; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20224 = _T_16140 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_4 = _T_20224 | _T_11616; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20241 = _T_16157 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_5 = _T_20241 | _T_11625; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20258 = _T_16174 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_6 = _T_20258 | _T_11634; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20275 = _T_16191 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_7 = _T_20275 | _T_11643; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20292 = _T_16208 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_8 = _T_20292 | _T_11652; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20309 = _T_16225 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_9 = _T_20309 | _T_11661; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20326 = _T_16242 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_10 = _T_20326 | _T_11670; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20343 = _T_16259 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_11 = _T_20343 | _T_11679; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20360 = _T_16276 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_12 = _T_20360 | _T_11688; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20377 = _T_16293 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_13 = _T_20377 | _T_11697; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20394 = _T_16310 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_14 = _T_20394 | _T_11706; // @[ifu_bp_ctl.scala 521:223]
  wire  _T_20411 = _T_16327 & _T_6924; // @[ifu_bp_ctl.scala 521:110]
  wire  bht_bank_sel_1_15_15 = _T_20411 | _T_11715; // @[ifu_bp_ctl.scala 521:223]
  rvclkhdr rvclkhdr ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en)
  );
  rvclkhdr rvclkhdr_1 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en)
  );
  rvclkhdr rvclkhdr_2 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en)
  );
  rvclkhdr rvclkhdr_3 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en)
  );
  rvclkhdr rvclkhdr_4 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_4_io_clk),
    .io_en(rvclkhdr_4_io_en)
  );
  rvclkhdr rvclkhdr_5 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_5_io_clk),
    .io_en(rvclkhdr_5_io_en)
  );
  rvclkhdr rvclkhdr_6 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_6_io_clk),
    .io_en(rvclkhdr_6_io_en)
  );
  rvclkhdr rvclkhdr_7 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_7_io_clk),
    .io_en(rvclkhdr_7_io_en)
  );
  rvclkhdr rvclkhdr_8 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_8_io_clk),
    .io_en(rvclkhdr_8_io_en)
  );
  rvclkhdr rvclkhdr_9 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_9_io_clk),
    .io_en(rvclkhdr_9_io_en)
  );
  rvclkhdr rvclkhdr_10 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_10_io_clk),
    .io_en(rvclkhdr_10_io_en)
  );
  rvclkhdr rvclkhdr_11 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_11_io_clk),
    .io_en(rvclkhdr_11_io_en)
  );
  rvclkhdr rvclkhdr_12 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_12_io_clk),
    .io_en(rvclkhdr_12_io_en)
  );
  rvclkhdr rvclkhdr_13 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_13_io_clk),
    .io_en(rvclkhdr_13_io_en)
  );
  rvclkhdr rvclkhdr_14 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_14_io_clk),
    .io_en(rvclkhdr_14_io_en)
  );
  rvclkhdr rvclkhdr_15 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_15_io_clk),
    .io_en(rvclkhdr_15_io_en)
  );
  rvclkhdr rvclkhdr_16 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_16_io_clk),
    .io_en(rvclkhdr_16_io_en)
  );
  rvclkhdr rvclkhdr_17 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_17_io_clk),
    .io_en(rvclkhdr_17_io_en)
  );
  rvclkhdr rvclkhdr_18 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_18_io_clk),
    .io_en(rvclkhdr_18_io_en)
  );
  rvclkhdr rvclkhdr_19 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_19_io_clk),
    .io_en(rvclkhdr_19_io_en)
  );
  rvclkhdr rvclkhdr_20 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_20_io_clk),
    .io_en(rvclkhdr_20_io_en)
  );
  rvclkhdr rvclkhdr_21 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_21_io_clk),
    .io_en(rvclkhdr_21_io_en)
  );
  rvclkhdr rvclkhdr_22 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_22_io_clk),
    .io_en(rvclkhdr_22_io_en)
  );
  rvclkhdr rvclkhdr_23 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_23_io_clk),
    .io_en(rvclkhdr_23_io_en)
  );
  rvclkhdr rvclkhdr_24 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_24_io_clk),
    .io_en(rvclkhdr_24_io_en)
  );
  rvclkhdr rvclkhdr_25 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_25_io_clk),
    .io_en(rvclkhdr_25_io_en)
  );
  rvclkhdr rvclkhdr_26 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_26_io_clk),
    .io_en(rvclkhdr_26_io_en)
  );
  rvclkhdr rvclkhdr_27 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_27_io_clk),
    .io_en(rvclkhdr_27_io_en)
  );
  rvclkhdr rvclkhdr_28 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_28_io_clk),
    .io_en(rvclkhdr_28_io_en)
  );
  rvclkhdr rvclkhdr_29 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_29_io_clk),
    .io_en(rvclkhdr_29_io_en)
  );
  rvclkhdr rvclkhdr_30 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_30_io_clk),
    .io_en(rvclkhdr_30_io_en)
  );
  rvclkhdr rvclkhdr_31 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_31_io_clk),
    .io_en(rvclkhdr_31_io_en)
  );
  rvclkhdr rvclkhdr_32 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_32_io_clk),
    .io_en(rvclkhdr_32_io_en)
  );
  rvclkhdr rvclkhdr_33 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_33_io_clk),
    .io_en(rvclkhdr_33_io_en)
  );
  rvclkhdr rvclkhdr_34 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_34_io_clk),
    .io_en(rvclkhdr_34_io_en)
  );
  rvclkhdr rvclkhdr_35 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_35_io_clk),
    .io_en(rvclkhdr_35_io_en)
  );
  rvclkhdr rvclkhdr_36 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_36_io_clk),
    .io_en(rvclkhdr_36_io_en)
  );
  rvclkhdr rvclkhdr_37 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_37_io_clk),
    .io_en(rvclkhdr_37_io_en)
  );
  rvclkhdr rvclkhdr_38 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_38_io_clk),
    .io_en(rvclkhdr_38_io_en)
  );
  rvclkhdr rvclkhdr_39 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_39_io_clk),
    .io_en(rvclkhdr_39_io_en)
  );
  rvclkhdr rvclkhdr_40 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_40_io_clk),
    .io_en(rvclkhdr_40_io_en)
  );
  rvclkhdr rvclkhdr_41 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_41_io_clk),
    .io_en(rvclkhdr_41_io_en)
  );
  rvclkhdr rvclkhdr_42 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_42_io_clk),
    .io_en(rvclkhdr_42_io_en)
  );
  rvclkhdr rvclkhdr_43 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_43_io_clk),
    .io_en(rvclkhdr_43_io_en)
  );
  rvclkhdr rvclkhdr_44 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_44_io_clk),
    .io_en(rvclkhdr_44_io_en)
  );
  rvclkhdr rvclkhdr_45 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_45_io_clk),
    .io_en(rvclkhdr_45_io_en)
  );
  rvclkhdr rvclkhdr_46 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_46_io_clk),
    .io_en(rvclkhdr_46_io_en)
  );
  rvclkhdr rvclkhdr_47 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_47_io_clk),
    .io_en(rvclkhdr_47_io_en)
  );
  rvclkhdr rvclkhdr_48 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_48_io_clk),
    .io_en(rvclkhdr_48_io_en)
  );
  rvclkhdr rvclkhdr_49 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_49_io_clk),
    .io_en(rvclkhdr_49_io_en)
  );
  rvclkhdr rvclkhdr_50 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_50_io_clk),
    .io_en(rvclkhdr_50_io_en)
  );
  rvclkhdr rvclkhdr_51 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_51_io_clk),
    .io_en(rvclkhdr_51_io_en)
  );
  rvclkhdr rvclkhdr_52 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_52_io_clk),
    .io_en(rvclkhdr_52_io_en)
  );
  rvclkhdr rvclkhdr_53 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_53_io_clk),
    .io_en(rvclkhdr_53_io_en)
  );
  rvclkhdr rvclkhdr_54 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_54_io_clk),
    .io_en(rvclkhdr_54_io_en)
  );
  rvclkhdr rvclkhdr_55 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_55_io_clk),
    .io_en(rvclkhdr_55_io_en)
  );
  rvclkhdr rvclkhdr_56 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_56_io_clk),
    .io_en(rvclkhdr_56_io_en)
  );
  rvclkhdr rvclkhdr_57 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_57_io_clk),
    .io_en(rvclkhdr_57_io_en)
  );
  rvclkhdr rvclkhdr_58 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_58_io_clk),
    .io_en(rvclkhdr_58_io_en)
  );
  rvclkhdr rvclkhdr_59 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_59_io_clk),
    .io_en(rvclkhdr_59_io_en)
  );
  rvclkhdr rvclkhdr_60 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_60_io_clk),
    .io_en(rvclkhdr_60_io_en)
  );
  rvclkhdr rvclkhdr_61 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_61_io_clk),
    .io_en(rvclkhdr_61_io_en)
  );
  rvclkhdr rvclkhdr_62 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_62_io_clk),
    .io_en(rvclkhdr_62_io_en)
  );
  rvclkhdr rvclkhdr_63 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_63_io_clk),
    .io_en(rvclkhdr_63_io_en)
  );
  rvclkhdr rvclkhdr_64 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_64_io_clk),
    .io_en(rvclkhdr_64_io_en)
  );
  rvclkhdr rvclkhdr_65 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_65_io_clk),
    .io_en(rvclkhdr_65_io_en)
  );
  rvclkhdr rvclkhdr_66 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_66_io_clk),
    .io_en(rvclkhdr_66_io_en)
  );
  rvclkhdr rvclkhdr_67 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_67_io_clk),
    .io_en(rvclkhdr_67_io_en)
  );
  rvclkhdr rvclkhdr_68 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_68_io_clk),
    .io_en(rvclkhdr_68_io_en)
  );
  rvclkhdr rvclkhdr_69 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_69_io_clk),
    .io_en(rvclkhdr_69_io_en)
  );
  rvclkhdr rvclkhdr_70 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_70_io_clk),
    .io_en(rvclkhdr_70_io_en)
  );
  rvclkhdr rvclkhdr_71 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_71_io_clk),
    .io_en(rvclkhdr_71_io_en)
  );
  rvclkhdr rvclkhdr_72 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_72_io_clk),
    .io_en(rvclkhdr_72_io_en)
  );
  rvclkhdr rvclkhdr_73 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_73_io_clk),
    .io_en(rvclkhdr_73_io_en)
  );
  rvclkhdr rvclkhdr_74 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_74_io_clk),
    .io_en(rvclkhdr_74_io_en)
  );
  rvclkhdr rvclkhdr_75 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_75_io_clk),
    .io_en(rvclkhdr_75_io_en)
  );
  rvclkhdr rvclkhdr_76 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_76_io_clk),
    .io_en(rvclkhdr_76_io_en)
  );
  rvclkhdr rvclkhdr_77 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_77_io_clk),
    .io_en(rvclkhdr_77_io_en)
  );
  rvclkhdr rvclkhdr_78 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_78_io_clk),
    .io_en(rvclkhdr_78_io_en)
  );
  rvclkhdr rvclkhdr_79 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_79_io_clk),
    .io_en(rvclkhdr_79_io_en)
  );
  rvclkhdr rvclkhdr_80 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_80_io_clk),
    .io_en(rvclkhdr_80_io_en)
  );
  rvclkhdr rvclkhdr_81 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_81_io_clk),
    .io_en(rvclkhdr_81_io_en)
  );
  rvclkhdr rvclkhdr_82 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_82_io_clk),
    .io_en(rvclkhdr_82_io_en)
  );
  rvclkhdr rvclkhdr_83 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_83_io_clk),
    .io_en(rvclkhdr_83_io_en)
  );
  rvclkhdr rvclkhdr_84 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_84_io_clk),
    .io_en(rvclkhdr_84_io_en)
  );
  rvclkhdr rvclkhdr_85 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_85_io_clk),
    .io_en(rvclkhdr_85_io_en)
  );
  rvclkhdr rvclkhdr_86 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_86_io_clk),
    .io_en(rvclkhdr_86_io_en)
  );
  rvclkhdr rvclkhdr_87 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_87_io_clk),
    .io_en(rvclkhdr_87_io_en)
  );
  rvclkhdr rvclkhdr_88 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_88_io_clk),
    .io_en(rvclkhdr_88_io_en)
  );
  rvclkhdr rvclkhdr_89 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_89_io_clk),
    .io_en(rvclkhdr_89_io_en)
  );
  rvclkhdr rvclkhdr_90 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_90_io_clk),
    .io_en(rvclkhdr_90_io_en)
  );
  rvclkhdr rvclkhdr_91 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_91_io_clk),
    .io_en(rvclkhdr_91_io_en)
  );
  rvclkhdr rvclkhdr_92 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_92_io_clk),
    .io_en(rvclkhdr_92_io_en)
  );
  rvclkhdr rvclkhdr_93 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_93_io_clk),
    .io_en(rvclkhdr_93_io_en)
  );
  rvclkhdr rvclkhdr_94 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_94_io_clk),
    .io_en(rvclkhdr_94_io_en)
  );
  rvclkhdr rvclkhdr_95 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_95_io_clk),
    .io_en(rvclkhdr_95_io_en)
  );
  rvclkhdr rvclkhdr_96 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_96_io_clk),
    .io_en(rvclkhdr_96_io_en)
  );
  rvclkhdr rvclkhdr_97 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_97_io_clk),
    .io_en(rvclkhdr_97_io_en)
  );
  rvclkhdr rvclkhdr_98 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_98_io_clk),
    .io_en(rvclkhdr_98_io_en)
  );
  rvclkhdr rvclkhdr_99 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_99_io_clk),
    .io_en(rvclkhdr_99_io_en)
  );
  rvclkhdr rvclkhdr_100 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_100_io_clk),
    .io_en(rvclkhdr_100_io_en)
  );
  rvclkhdr rvclkhdr_101 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_101_io_clk),
    .io_en(rvclkhdr_101_io_en)
  );
  rvclkhdr rvclkhdr_102 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_102_io_clk),
    .io_en(rvclkhdr_102_io_en)
  );
  rvclkhdr rvclkhdr_103 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_103_io_clk),
    .io_en(rvclkhdr_103_io_en)
  );
  rvclkhdr rvclkhdr_104 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_104_io_clk),
    .io_en(rvclkhdr_104_io_en)
  );
  rvclkhdr rvclkhdr_105 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_105_io_clk),
    .io_en(rvclkhdr_105_io_en)
  );
  rvclkhdr rvclkhdr_106 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_106_io_clk),
    .io_en(rvclkhdr_106_io_en)
  );
  rvclkhdr rvclkhdr_107 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_107_io_clk),
    .io_en(rvclkhdr_107_io_en)
  );
  rvclkhdr rvclkhdr_108 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_108_io_clk),
    .io_en(rvclkhdr_108_io_en)
  );
  rvclkhdr rvclkhdr_109 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_109_io_clk),
    .io_en(rvclkhdr_109_io_en)
  );
  rvclkhdr rvclkhdr_110 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_110_io_clk),
    .io_en(rvclkhdr_110_io_en)
  );
  rvclkhdr rvclkhdr_111 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_111_io_clk),
    .io_en(rvclkhdr_111_io_en)
  );
  rvclkhdr rvclkhdr_112 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_112_io_clk),
    .io_en(rvclkhdr_112_io_en)
  );
  rvclkhdr rvclkhdr_113 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_113_io_clk),
    .io_en(rvclkhdr_113_io_en)
  );
  rvclkhdr rvclkhdr_114 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_114_io_clk),
    .io_en(rvclkhdr_114_io_en)
  );
  rvclkhdr rvclkhdr_115 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_115_io_clk),
    .io_en(rvclkhdr_115_io_en)
  );
  rvclkhdr rvclkhdr_116 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_116_io_clk),
    .io_en(rvclkhdr_116_io_en)
  );
  rvclkhdr rvclkhdr_117 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_117_io_clk),
    .io_en(rvclkhdr_117_io_en)
  );
  rvclkhdr rvclkhdr_118 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_118_io_clk),
    .io_en(rvclkhdr_118_io_en)
  );
  rvclkhdr rvclkhdr_119 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_119_io_clk),
    .io_en(rvclkhdr_119_io_en)
  );
  rvclkhdr rvclkhdr_120 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_120_io_clk),
    .io_en(rvclkhdr_120_io_en)
  );
  rvclkhdr rvclkhdr_121 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_121_io_clk),
    .io_en(rvclkhdr_121_io_en)
  );
  rvclkhdr rvclkhdr_122 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_122_io_clk),
    .io_en(rvclkhdr_122_io_en)
  );
  rvclkhdr rvclkhdr_123 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_123_io_clk),
    .io_en(rvclkhdr_123_io_en)
  );
  rvclkhdr rvclkhdr_124 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_124_io_clk),
    .io_en(rvclkhdr_124_io_en)
  );
  rvclkhdr rvclkhdr_125 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_125_io_clk),
    .io_en(rvclkhdr_125_io_en)
  );
  rvclkhdr rvclkhdr_126 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_126_io_clk),
    .io_en(rvclkhdr_126_io_en)
  );
  rvclkhdr rvclkhdr_127 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_127_io_clk),
    .io_en(rvclkhdr_127_io_en)
  );
  rvclkhdr rvclkhdr_128 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_128_io_clk),
    .io_en(rvclkhdr_128_io_en)
  );
  rvclkhdr rvclkhdr_129 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_129_io_clk),
    .io_en(rvclkhdr_129_io_en)
  );
  rvclkhdr rvclkhdr_130 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_130_io_clk),
    .io_en(rvclkhdr_130_io_en)
  );
  rvclkhdr rvclkhdr_131 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_131_io_clk),
    .io_en(rvclkhdr_131_io_en)
  );
  rvclkhdr rvclkhdr_132 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_132_io_clk),
    .io_en(rvclkhdr_132_io_en)
  );
  rvclkhdr rvclkhdr_133 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_133_io_clk),
    .io_en(rvclkhdr_133_io_en)
  );
  rvclkhdr rvclkhdr_134 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_134_io_clk),
    .io_en(rvclkhdr_134_io_en)
  );
  rvclkhdr rvclkhdr_135 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_135_io_clk),
    .io_en(rvclkhdr_135_io_en)
  );
  rvclkhdr rvclkhdr_136 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_136_io_clk),
    .io_en(rvclkhdr_136_io_en)
  );
  rvclkhdr rvclkhdr_137 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_137_io_clk),
    .io_en(rvclkhdr_137_io_en)
  );
  rvclkhdr rvclkhdr_138 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_138_io_clk),
    .io_en(rvclkhdr_138_io_en)
  );
  rvclkhdr rvclkhdr_139 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_139_io_clk),
    .io_en(rvclkhdr_139_io_en)
  );
  rvclkhdr rvclkhdr_140 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_140_io_clk),
    .io_en(rvclkhdr_140_io_en)
  );
  rvclkhdr rvclkhdr_141 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_141_io_clk),
    .io_en(rvclkhdr_141_io_en)
  );
  rvclkhdr rvclkhdr_142 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_142_io_clk),
    .io_en(rvclkhdr_142_io_en)
  );
  rvclkhdr rvclkhdr_143 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_143_io_clk),
    .io_en(rvclkhdr_143_io_en)
  );
  rvclkhdr rvclkhdr_144 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_144_io_clk),
    .io_en(rvclkhdr_144_io_en)
  );
  rvclkhdr rvclkhdr_145 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_145_io_clk),
    .io_en(rvclkhdr_145_io_en)
  );
  rvclkhdr rvclkhdr_146 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_146_io_clk),
    .io_en(rvclkhdr_146_io_en)
  );
  rvclkhdr rvclkhdr_147 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_147_io_clk),
    .io_en(rvclkhdr_147_io_en)
  );
  rvclkhdr rvclkhdr_148 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_148_io_clk),
    .io_en(rvclkhdr_148_io_en)
  );
  rvclkhdr rvclkhdr_149 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_149_io_clk),
    .io_en(rvclkhdr_149_io_en)
  );
  rvclkhdr rvclkhdr_150 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_150_io_clk),
    .io_en(rvclkhdr_150_io_en)
  );
  rvclkhdr rvclkhdr_151 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_151_io_clk),
    .io_en(rvclkhdr_151_io_en)
  );
  rvclkhdr rvclkhdr_152 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_152_io_clk),
    .io_en(rvclkhdr_152_io_en)
  );
  rvclkhdr rvclkhdr_153 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_153_io_clk),
    .io_en(rvclkhdr_153_io_en)
  );
  rvclkhdr rvclkhdr_154 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_154_io_clk),
    .io_en(rvclkhdr_154_io_en)
  );
  rvclkhdr rvclkhdr_155 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_155_io_clk),
    .io_en(rvclkhdr_155_io_en)
  );
  rvclkhdr rvclkhdr_156 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_156_io_clk),
    .io_en(rvclkhdr_156_io_en)
  );
  rvclkhdr rvclkhdr_157 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_157_io_clk),
    .io_en(rvclkhdr_157_io_en)
  );
  rvclkhdr rvclkhdr_158 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_158_io_clk),
    .io_en(rvclkhdr_158_io_en)
  );
  rvclkhdr rvclkhdr_159 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_159_io_clk),
    .io_en(rvclkhdr_159_io_en)
  );
  rvclkhdr rvclkhdr_160 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_160_io_clk),
    .io_en(rvclkhdr_160_io_en)
  );
  rvclkhdr rvclkhdr_161 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_161_io_clk),
    .io_en(rvclkhdr_161_io_en)
  );
  rvclkhdr rvclkhdr_162 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_162_io_clk),
    .io_en(rvclkhdr_162_io_en)
  );
  rvclkhdr rvclkhdr_163 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_163_io_clk),
    .io_en(rvclkhdr_163_io_en)
  );
  rvclkhdr rvclkhdr_164 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_164_io_clk),
    .io_en(rvclkhdr_164_io_en)
  );
  rvclkhdr rvclkhdr_165 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_165_io_clk),
    .io_en(rvclkhdr_165_io_en)
  );
  rvclkhdr rvclkhdr_166 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_166_io_clk),
    .io_en(rvclkhdr_166_io_en)
  );
  rvclkhdr rvclkhdr_167 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_167_io_clk),
    .io_en(rvclkhdr_167_io_en)
  );
  rvclkhdr rvclkhdr_168 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_168_io_clk),
    .io_en(rvclkhdr_168_io_en)
  );
  rvclkhdr rvclkhdr_169 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_169_io_clk),
    .io_en(rvclkhdr_169_io_en)
  );
  rvclkhdr rvclkhdr_170 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_170_io_clk),
    .io_en(rvclkhdr_170_io_en)
  );
  rvclkhdr rvclkhdr_171 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_171_io_clk),
    .io_en(rvclkhdr_171_io_en)
  );
  rvclkhdr rvclkhdr_172 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_172_io_clk),
    .io_en(rvclkhdr_172_io_en)
  );
  rvclkhdr rvclkhdr_173 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_173_io_clk),
    .io_en(rvclkhdr_173_io_en)
  );
  rvclkhdr rvclkhdr_174 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_174_io_clk),
    .io_en(rvclkhdr_174_io_en)
  );
  rvclkhdr rvclkhdr_175 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_175_io_clk),
    .io_en(rvclkhdr_175_io_en)
  );
  rvclkhdr rvclkhdr_176 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_176_io_clk),
    .io_en(rvclkhdr_176_io_en)
  );
  rvclkhdr rvclkhdr_177 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_177_io_clk),
    .io_en(rvclkhdr_177_io_en)
  );
  rvclkhdr rvclkhdr_178 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_178_io_clk),
    .io_en(rvclkhdr_178_io_en)
  );
  rvclkhdr rvclkhdr_179 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_179_io_clk),
    .io_en(rvclkhdr_179_io_en)
  );
  rvclkhdr rvclkhdr_180 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_180_io_clk),
    .io_en(rvclkhdr_180_io_en)
  );
  rvclkhdr rvclkhdr_181 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_181_io_clk),
    .io_en(rvclkhdr_181_io_en)
  );
  rvclkhdr rvclkhdr_182 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_182_io_clk),
    .io_en(rvclkhdr_182_io_en)
  );
  rvclkhdr rvclkhdr_183 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_183_io_clk),
    .io_en(rvclkhdr_183_io_en)
  );
  rvclkhdr rvclkhdr_184 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_184_io_clk),
    .io_en(rvclkhdr_184_io_en)
  );
  rvclkhdr rvclkhdr_185 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_185_io_clk),
    .io_en(rvclkhdr_185_io_en)
  );
  rvclkhdr rvclkhdr_186 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_186_io_clk),
    .io_en(rvclkhdr_186_io_en)
  );
  rvclkhdr rvclkhdr_187 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_187_io_clk),
    .io_en(rvclkhdr_187_io_en)
  );
  rvclkhdr rvclkhdr_188 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_188_io_clk),
    .io_en(rvclkhdr_188_io_en)
  );
  rvclkhdr rvclkhdr_189 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_189_io_clk),
    .io_en(rvclkhdr_189_io_en)
  );
  rvclkhdr rvclkhdr_190 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_190_io_clk),
    .io_en(rvclkhdr_190_io_en)
  );
  rvclkhdr rvclkhdr_191 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_191_io_clk),
    .io_en(rvclkhdr_191_io_en)
  );
  rvclkhdr rvclkhdr_192 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_192_io_clk),
    .io_en(rvclkhdr_192_io_en)
  );
  rvclkhdr rvclkhdr_193 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_193_io_clk),
    .io_en(rvclkhdr_193_io_en)
  );
  rvclkhdr rvclkhdr_194 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_194_io_clk),
    .io_en(rvclkhdr_194_io_en)
  );
  rvclkhdr rvclkhdr_195 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_195_io_clk),
    .io_en(rvclkhdr_195_io_en)
  );
  rvclkhdr rvclkhdr_196 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_196_io_clk),
    .io_en(rvclkhdr_196_io_en)
  );
  rvclkhdr rvclkhdr_197 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_197_io_clk),
    .io_en(rvclkhdr_197_io_en)
  );
  rvclkhdr rvclkhdr_198 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_198_io_clk),
    .io_en(rvclkhdr_198_io_en)
  );
  rvclkhdr rvclkhdr_199 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_199_io_clk),
    .io_en(rvclkhdr_199_io_en)
  );
  rvclkhdr rvclkhdr_200 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_200_io_clk),
    .io_en(rvclkhdr_200_io_en)
  );
  rvclkhdr rvclkhdr_201 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_201_io_clk),
    .io_en(rvclkhdr_201_io_en)
  );
  rvclkhdr rvclkhdr_202 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_202_io_clk),
    .io_en(rvclkhdr_202_io_en)
  );
  rvclkhdr rvclkhdr_203 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_203_io_clk),
    .io_en(rvclkhdr_203_io_en)
  );
  rvclkhdr rvclkhdr_204 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_204_io_clk),
    .io_en(rvclkhdr_204_io_en)
  );
  rvclkhdr rvclkhdr_205 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_205_io_clk),
    .io_en(rvclkhdr_205_io_en)
  );
  rvclkhdr rvclkhdr_206 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_206_io_clk),
    .io_en(rvclkhdr_206_io_en)
  );
  rvclkhdr rvclkhdr_207 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_207_io_clk),
    .io_en(rvclkhdr_207_io_en)
  );
  rvclkhdr rvclkhdr_208 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_208_io_clk),
    .io_en(rvclkhdr_208_io_en)
  );
  rvclkhdr rvclkhdr_209 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_209_io_clk),
    .io_en(rvclkhdr_209_io_en)
  );
  rvclkhdr rvclkhdr_210 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_210_io_clk),
    .io_en(rvclkhdr_210_io_en)
  );
  rvclkhdr rvclkhdr_211 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_211_io_clk),
    .io_en(rvclkhdr_211_io_en)
  );
  rvclkhdr rvclkhdr_212 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_212_io_clk),
    .io_en(rvclkhdr_212_io_en)
  );
  rvclkhdr rvclkhdr_213 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_213_io_clk),
    .io_en(rvclkhdr_213_io_en)
  );
  rvclkhdr rvclkhdr_214 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_214_io_clk),
    .io_en(rvclkhdr_214_io_en)
  );
  rvclkhdr rvclkhdr_215 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_215_io_clk),
    .io_en(rvclkhdr_215_io_en)
  );
  rvclkhdr rvclkhdr_216 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_216_io_clk),
    .io_en(rvclkhdr_216_io_en)
  );
  rvclkhdr rvclkhdr_217 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_217_io_clk),
    .io_en(rvclkhdr_217_io_en)
  );
  rvclkhdr rvclkhdr_218 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_218_io_clk),
    .io_en(rvclkhdr_218_io_en)
  );
  rvclkhdr rvclkhdr_219 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_219_io_clk),
    .io_en(rvclkhdr_219_io_en)
  );
  rvclkhdr rvclkhdr_220 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_220_io_clk),
    .io_en(rvclkhdr_220_io_en)
  );
  rvclkhdr rvclkhdr_221 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_221_io_clk),
    .io_en(rvclkhdr_221_io_en)
  );
  rvclkhdr rvclkhdr_222 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_222_io_clk),
    .io_en(rvclkhdr_222_io_en)
  );
  rvclkhdr rvclkhdr_223 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_223_io_clk),
    .io_en(rvclkhdr_223_io_en)
  );
  rvclkhdr rvclkhdr_224 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_224_io_clk),
    .io_en(rvclkhdr_224_io_en)
  );
  rvclkhdr rvclkhdr_225 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_225_io_clk),
    .io_en(rvclkhdr_225_io_en)
  );
  rvclkhdr rvclkhdr_226 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_226_io_clk),
    .io_en(rvclkhdr_226_io_en)
  );
  rvclkhdr rvclkhdr_227 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_227_io_clk),
    .io_en(rvclkhdr_227_io_en)
  );
  rvclkhdr rvclkhdr_228 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_228_io_clk),
    .io_en(rvclkhdr_228_io_en)
  );
  rvclkhdr rvclkhdr_229 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_229_io_clk),
    .io_en(rvclkhdr_229_io_en)
  );
  rvclkhdr rvclkhdr_230 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_230_io_clk),
    .io_en(rvclkhdr_230_io_en)
  );
  rvclkhdr rvclkhdr_231 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_231_io_clk),
    .io_en(rvclkhdr_231_io_en)
  );
  rvclkhdr rvclkhdr_232 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_232_io_clk),
    .io_en(rvclkhdr_232_io_en)
  );
  rvclkhdr rvclkhdr_233 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_233_io_clk),
    .io_en(rvclkhdr_233_io_en)
  );
  rvclkhdr rvclkhdr_234 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_234_io_clk),
    .io_en(rvclkhdr_234_io_en)
  );
  rvclkhdr rvclkhdr_235 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_235_io_clk),
    .io_en(rvclkhdr_235_io_en)
  );
  rvclkhdr rvclkhdr_236 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_236_io_clk),
    .io_en(rvclkhdr_236_io_en)
  );
  rvclkhdr rvclkhdr_237 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_237_io_clk),
    .io_en(rvclkhdr_237_io_en)
  );
  rvclkhdr rvclkhdr_238 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_238_io_clk),
    .io_en(rvclkhdr_238_io_en)
  );
  rvclkhdr rvclkhdr_239 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_239_io_clk),
    .io_en(rvclkhdr_239_io_en)
  );
  rvclkhdr rvclkhdr_240 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_240_io_clk),
    .io_en(rvclkhdr_240_io_en)
  );
  rvclkhdr rvclkhdr_241 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_241_io_clk),
    .io_en(rvclkhdr_241_io_en)
  );
  rvclkhdr rvclkhdr_242 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_242_io_clk),
    .io_en(rvclkhdr_242_io_en)
  );
  rvclkhdr rvclkhdr_243 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_243_io_clk),
    .io_en(rvclkhdr_243_io_en)
  );
  rvclkhdr rvclkhdr_244 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_244_io_clk),
    .io_en(rvclkhdr_244_io_en)
  );
  rvclkhdr rvclkhdr_245 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_245_io_clk),
    .io_en(rvclkhdr_245_io_en)
  );
  rvclkhdr rvclkhdr_246 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_246_io_clk),
    .io_en(rvclkhdr_246_io_en)
  );
  rvclkhdr rvclkhdr_247 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_247_io_clk),
    .io_en(rvclkhdr_247_io_en)
  );
  rvclkhdr rvclkhdr_248 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_248_io_clk),
    .io_en(rvclkhdr_248_io_en)
  );
  rvclkhdr rvclkhdr_249 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_249_io_clk),
    .io_en(rvclkhdr_249_io_en)
  );
  rvclkhdr rvclkhdr_250 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_250_io_clk),
    .io_en(rvclkhdr_250_io_en)
  );
  rvclkhdr rvclkhdr_251 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_251_io_clk),
    .io_en(rvclkhdr_251_io_en)
  );
  rvclkhdr rvclkhdr_252 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_252_io_clk),
    .io_en(rvclkhdr_252_io_en)
  );
  rvclkhdr rvclkhdr_253 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_253_io_clk),
    .io_en(rvclkhdr_253_io_en)
  );
  rvclkhdr rvclkhdr_254 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_254_io_clk),
    .io_en(rvclkhdr_254_io_en)
  );
  rvclkhdr rvclkhdr_255 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_255_io_clk),
    .io_en(rvclkhdr_255_io_en)
  );
  rvclkhdr rvclkhdr_256 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_256_io_clk),
    .io_en(rvclkhdr_256_io_en)
  );
  rvclkhdr rvclkhdr_257 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_257_io_clk),
    .io_en(rvclkhdr_257_io_en)
  );
  rvclkhdr rvclkhdr_258 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_258_io_clk),
    .io_en(rvclkhdr_258_io_en)
  );
  rvclkhdr rvclkhdr_259 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_259_io_clk),
    .io_en(rvclkhdr_259_io_en)
  );
  rvclkhdr rvclkhdr_260 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_260_io_clk),
    .io_en(rvclkhdr_260_io_en)
  );
  rvclkhdr rvclkhdr_261 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_261_io_clk),
    .io_en(rvclkhdr_261_io_en)
  );
  rvclkhdr rvclkhdr_262 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_262_io_clk),
    .io_en(rvclkhdr_262_io_en)
  );
  rvclkhdr rvclkhdr_263 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_263_io_clk),
    .io_en(rvclkhdr_263_io_en)
  );
  rvclkhdr rvclkhdr_264 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_264_io_clk),
    .io_en(rvclkhdr_264_io_en)
  );
  rvclkhdr rvclkhdr_265 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_265_io_clk),
    .io_en(rvclkhdr_265_io_en)
  );
  rvclkhdr rvclkhdr_266 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_266_io_clk),
    .io_en(rvclkhdr_266_io_en)
  );
  rvclkhdr rvclkhdr_267 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_267_io_clk),
    .io_en(rvclkhdr_267_io_en)
  );
  rvclkhdr rvclkhdr_268 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_268_io_clk),
    .io_en(rvclkhdr_268_io_en)
  );
  rvclkhdr rvclkhdr_269 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_269_io_clk),
    .io_en(rvclkhdr_269_io_en)
  );
  rvclkhdr rvclkhdr_270 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_270_io_clk),
    .io_en(rvclkhdr_270_io_en)
  );
  rvclkhdr rvclkhdr_271 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_271_io_clk),
    .io_en(rvclkhdr_271_io_en)
  );
  rvclkhdr rvclkhdr_272 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_272_io_clk),
    .io_en(rvclkhdr_272_io_en)
  );
  rvclkhdr rvclkhdr_273 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_273_io_clk),
    .io_en(rvclkhdr_273_io_en)
  );
  rvclkhdr rvclkhdr_274 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_274_io_clk),
    .io_en(rvclkhdr_274_io_en)
  );
  rvclkhdr rvclkhdr_275 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_275_io_clk),
    .io_en(rvclkhdr_275_io_en)
  );
  rvclkhdr rvclkhdr_276 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_276_io_clk),
    .io_en(rvclkhdr_276_io_en)
  );
  rvclkhdr rvclkhdr_277 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_277_io_clk),
    .io_en(rvclkhdr_277_io_en)
  );
  rvclkhdr rvclkhdr_278 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_278_io_clk),
    .io_en(rvclkhdr_278_io_en)
  );
  rvclkhdr rvclkhdr_279 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_279_io_clk),
    .io_en(rvclkhdr_279_io_en)
  );
  rvclkhdr rvclkhdr_280 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_280_io_clk),
    .io_en(rvclkhdr_280_io_en)
  );
  rvclkhdr rvclkhdr_281 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_281_io_clk),
    .io_en(rvclkhdr_281_io_en)
  );
  rvclkhdr rvclkhdr_282 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_282_io_clk),
    .io_en(rvclkhdr_282_io_en)
  );
  rvclkhdr rvclkhdr_283 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_283_io_clk),
    .io_en(rvclkhdr_283_io_en)
  );
  rvclkhdr rvclkhdr_284 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_284_io_clk),
    .io_en(rvclkhdr_284_io_en)
  );
  rvclkhdr rvclkhdr_285 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_285_io_clk),
    .io_en(rvclkhdr_285_io_en)
  );
  rvclkhdr rvclkhdr_286 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_286_io_clk),
    .io_en(rvclkhdr_286_io_en)
  );
  rvclkhdr rvclkhdr_287 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_287_io_clk),
    .io_en(rvclkhdr_287_io_en)
  );
  rvclkhdr rvclkhdr_288 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_288_io_clk),
    .io_en(rvclkhdr_288_io_en)
  );
  rvclkhdr rvclkhdr_289 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_289_io_clk),
    .io_en(rvclkhdr_289_io_en)
  );
  rvclkhdr rvclkhdr_290 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_290_io_clk),
    .io_en(rvclkhdr_290_io_en)
  );
  rvclkhdr rvclkhdr_291 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_291_io_clk),
    .io_en(rvclkhdr_291_io_en)
  );
  rvclkhdr rvclkhdr_292 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_292_io_clk),
    .io_en(rvclkhdr_292_io_en)
  );
  rvclkhdr rvclkhdr_293 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_293_io_clk),
    .io_en(rvclkhdr_293_io_en)
  );
  rvclkhdr rvclkhdr_294 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_294_io_clk),
    .io_en(rvclkhdr_294_io_en)
  );
  rvclkhdr rvclkhdr_295 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_295_io_clk),
    .io_en(rvclkhdr_295_io_en)
  );
  rvclkhdr rvclkhdr_296 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_296_io_clk),
    .io_en(rvclkhdr_296_io_en)
  );
  rvclkhdr rvclkhdr_297 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_297_io_clk),
    .io_en(rvclkhdr_297_io_en)
  );
  rvclkhdr rvclkhdr_298 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_298_io_clk),
    .io_en(rvclkhdr_298_io_en)
  );
  rvclkhdr rvclkhdr_299 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_299_io_clk),
    .io_en(rvclkhdr_299_io_en)
  );
  rvclkhdr rvclkhdr_300 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_300_io_clk),
    .io_en(rvclkhdr_300_io_en)
  );
  rvclkhdr rvclkhdr_301 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_301_io_clk),
    .io_en(rvclkhdr_301_io_en)
  );
  rvclkhdr rvclkhdr_302 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_302_io_clk),
    .io_en(rvclkhdr_302_io_en)
  );
  rvclkhdr rvclkhdr_303 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_303_io_clk),
    .io_en(rvclkhdr_303_io_en)
  );
  rvclkhdr rvclkhdr_304 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_304_io_clk),
    .io_en(rvclkhdr_304_io_en)
  );
  rvclkhdr rvclkhdr_305 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_305_io_clk),
    .io_en(rvclkhdr_305_io_en)
  );
  rvclkhdr rvclkhdr_306 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_306_io_clk),
    .io_en(rvclkhdr_306_io_en)
  );
  rvclkhdr rvclkhdr_307 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_307_io_clk),
    .io_en(rvclkhdr_307_io_en)
  );
  rvclkhdr rvclkhdr_308 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_308_io_clk),
    .io_en(rvclkhdr_308_io_en)
  );
  rvclkhdr rvclkhdr_309 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_309_io_clk),
    .io_en(rvclkhdr_309_io_en)
  );
  rvclkhdr rvclkhdr_310 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_310_io_clk),
    .io_en(rvclkhdr_310_io_en)
  );
  rvclkhdr rvclkhdr_311 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_311_io_clk),
    .io_en(rvclkhdr_311_io_en)
  );
  rvclkhdr rvclkhdr_312 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_312_io_clk),
    .io_en(rvclkhdr_312_io_en)
  );
  rvclkhdr rvclkhdr_313 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_313_io_clk),
    .io_en(rvclkhdr_313_io_en)
  );
  rvclkhdr rvclkhdr_314 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_314_io_clk),
    .io_en(rvclkhdr_314_io_en)
  );
  rvclkhdr rvclkhdr_315 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_315_io_clk),
    .io_en(rvclkhdr_315_io_en)
  );
  rvclkhdr rvclkhdr_316 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_316_io_clk),
    .io_en(rvclkhdr_316_io_en)
  );
  rvclkhdr rvclkhdr_317 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_317_io_clk),
    .io_en(rvclkhdr_317_io_en)
  );
  rvclkhdr rvclkhdr_318 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_318_io_clk),
    .io_en(rvclkhdr_318_io_en)
  );
  rvclkhdr rvclkhdr_319 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_319_io_clk),
    .io_en(rvclkhdr_319_io_en)
  );
  rvclkhdr rvclkhdr_320 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_320_io_clk),
    .io_en(rvclkhdr_320_io_en)
  );
  rvclkhdr rvclkhdr_321 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_321_io_clk),
    .io_en(rvclkhdr_321_io_en)
  );
  rvclkhdr rvclkhdr_322 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_322_io_clk),
    .io_en(rvclkhdr_322_io_en)
  );
  rvclkhdr rvclkhdr_323 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_323_io_clk),
    .io_en(rvclkhdr_323_io_en)
  );
  rvclkhdr rvclkhdr_324 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_324_io_clk),
    .io_en(rvclkhdr_324_io_en)
  );
  rvclkhdr rvclkhdr_325 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_325_io_clk),
    .io_en(rvclkhdr_325_io_en)
  );
  rvclkhdr rvclkhdr_326 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_326_io_clk),
    .io_en(rvclkhdr_326_io_en)
  );
  rvclkhdr rvclkhdr_327 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_327_io_clk),
    .io_en(rvclkhdr_327_io_en)
  );
  rvclkhdr rvclkhdr_328 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_328_io_clk),
    .io_en(rvclkhdr_328_io_en)
  );
  rvclkhdr rvclkhdr_329 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_329_io_clk),
    .io_en(rvclkhdr_329_io_en)
  );
  rvclkhdr rvclkhdr_330 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_330_io_clk),
    .io_en(rvclkhdr_330_io_en)
  );
  rvclkhdr rvclkhdr_331 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_331_io_clk),
    .io_en(rvclkhdr_331_io_en)
  );
  rvclkhdr rvclkhdr_332 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_332_io_clk),
    .io_en(rvclkhdr_332_io_en)
  );
  rvclkhdr rvclkhdr_333 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_333_io_clk),
    .io_en(rvclkhdr_333_io_en)
  );
  rvclkhdr rvclkhdr_334 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_334_io_clk),
    .io_en(rvclkhdr_334_io_en)
  );
  rvclkhdr rvclkhdr_335 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_335_io_clk),
    .io_en(rvclkhdr_335_io_en)
  );
  rvclkhdr rvclkhdr_336 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_336_io_clk),
    .io_en(rvclkhdr_336_io_en)
  );
  rvclkhdr rvclkhdr_337 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_337_io_clk),
    .io_en(rvclkhdr_337_io_en)
  );
  rvclkhdr rvclkhdr_338 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_338_io_clk),
    .io_en(rvclkhdr_338_io_en)
  );
  rvclkhdr rvclkhdr_339 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_339_io_clk),
    .io_en(rvclkhdr_339_io_en)
  );
  rvclkhdr rvclkhdr_340 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_340_io_clk),
    .io_en(rvclkhdr_340_io_en)
  );
  rvclkhdr rvclkhdr_341 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_341_io_clk),
    .io_en(rvclkhdr_341_io_en)
  );
  rvclkhdr rvclkhdr_342 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_342_io_clk),
    .io_en(rvclkhdr_342_io_en)
  );
  rvclkhdr rvclkhdr_343 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_343_io_clk),
    .io_en(rvclkhdr_343_io_en)
  );
  rvclkhdr rvclkhdr_344 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_344_io_clk),
    .io_en(rvclkhdr_344_io_en)
  );
  rvclkhdr rvclkhdr_345 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_345_io_clk),
    .io_en(rvclkhdr_345_io_en)
  );
  rvclkhdr rvclkhdr_346 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_346_io_clk),
    .io_en(rvclkhdr_346_io_en)
  );
  rvclkhdr rvclkhdr_347 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_347_io_clk),
    .io_en(rvclkhdr_347_io_en)
  );
  rvclkhdr rvclkhdr_348 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_348_io_clk),
    .io_en(rvclkhdr_348_io_en)
  );
  rvclkhdr rvclkhdr_349 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_349_io_clk),
    .io_en(rvclkhdr_349_io_en)
  );
  rvclkhdr rvclkhdr_350 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_350_io_clk),
    .io_en(rvclkhdr_350_io_en)
  );
  rvclkhdr rvclkhdr_351 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_351_io_clk),
    .io_en(rvclkhdr_351_io_en)
  );
  rvclkhdr rvclkhdr_352 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_352_io_clk),
    .io_en(rvclkhdr_352_io_en)
  );
  rvclkhdr rvclkhdr_353 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_353_io_clk),
    .io_en(rvclkhdr_353_io_en)
  );
  rvclkhdr rvclkhdr_354 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_354_io_clk),
    .io_en(rvclkhdr_354_io_en)
  );
  rvclkhdr rvclkhdr_355 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_355_io_clk),
    .io_en(rvclkhdr_355_io_en)
  );
  rvclkhdr rvclkhdr_356 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_356_io_clk),
    .io_en(rvclkhdr_356_io_en)
  );
  rvclkhdr rvclkhdr_357 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_357_io_clk),
    .io_en(rvclkhdr_357_io_en)
  );
  rvclkhdr rvclkhdr_358 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_358_io_clk),
    .io_en(rvclkhdr_358_io_en)
  );
  rvclkhdr rvclkhdr_359 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_359_io_clk),
    .io_en(rvclkhdr_359_io_en)
  );
  rvclkhdr rvclkhdr_360 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_360_io_clk),
    .io_en(rvclkhdr_360_io_en)
  );
  rvclkhdr rvclkhdr_361 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_361_io_clk),
    .io_en(rvclkhdr_361_io_en)
  );
  rvclkhdr rvclkhdr_362 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_362_io_clk),
    .io_en(rvclkhdr_362_io_en)
  );
  rvclkhdr rvclkhdr_363 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_363_io_clk),
    .io_en(rvclkhdr_363_io_en)
  );
  rvclkhdr rvclkhdr_364 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_364_io_clk),
    .io_en(rvclkhdr_364_io_en)
  );
  rvclkhdr rvclkhdr_365 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_365_io_clk),
    .io_en(rvclkhdr_365_io_en)
  );
  rvclkhdr rvclkhdr_366 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_366_io_clk),
    .io_en(rvclkhdr_366_io_en)
  );
  rvclkhdr rvclkhdr_367 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_367_io_clk),
    .io_en(rvclkhdr_367_io_en)
  );
  rvclkhdr rvclkhdr_368 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_368_io_clk),
    .io_en(rvclkhdr_368_io_en)
  );
  rvclkhdr rvclkhdr_369 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_369_io_clk),
    .io_en(rvclkhdr_369_io_en)
  );
  rvclkhdr rvclkhdr_370 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_370_io_clk),
    .io_en(rvclkhdr_370_io_en)
  );
  rvclkhdr rvclkhdr_371 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_371_io_clk),
    .io_en(rvclkhdr_371_io_en)
  );
  rvclkhdr rvclkhdr_372 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_372_io_clk),
    .io_en(rvclkhdr_372_io_en)
  );
  rvclkhdr rvclkhdr_373 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_373_io_clk),
    .io_en(rvclkhdr_373_io_en)
  );
  rvclkhdr rvclkhdr_374 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_374_io_clk),
    .io_en(rvclkhdr_374_io_en)
  );
  rvclkhdr rvclkhdr_375 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_375_io_clk),
    .io_en(rvclkhdr_375_io_en)
  );
  rvclkhdr rvclkhdr_376 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_376_io_clk),
    .io_en(rvclkhdr_376_io_en)
  );
  rvclkhdr rvclkhdr_377 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_377_io_clk),
    .io_en(rvclkhdr_377_io_en)
  );
  rvclkhdr rvclkhdr_378 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_378_io_clk),
    .io_en(rvclkhdr_378_io_en)
  );
  rvclkhdr rvclkhdr_379 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_379_io_clk),
    .io_en(rvclkhdr_379_io_en)
  );
  rvclkhdr rvclkhdr_380 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_380_io_clk),
    .io_en(rvclkhdr_380_io_en)
  );
  rvclkhdr rvclkhdr_381 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_381_io_clk),
    .io_en(rvclkhdr_381_io_en)
  );
  rvclkhdr rvclkhdr_382 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_382_io_clk),
    .io_en(rvclkhdr_382_io_en)
  );
  rvclkhdr rvclkhdr_383 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_383_io_clk),
    .io_en(rvclkhdr_383_io_en)
  );
  rvclkhdr rvclkhdr_384 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_384_io_clk),
    .io_en(rvclkhdr_384_io_en)
  );
  rvclkhdr rvclkhdr_385 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_385_io_clk),
    .io_en(rvclkhdr_385_io_en)
  );
  rvclkhdr rvclkhdr_386 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_386_io_clk),
    .io_en(rvclkhdr_386_io_en)
  );
  rvclkhdr rvclkhdr_387 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_387_io_clk),
    .io_en(rvclkhdr_387_io_en)
  );
  rvclkhdr rvclkhdr_388 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_388_io_clk),
    .io_en(rvclkhdr_388_io_en)
  );
  rvclkhdr rvclkhdr_389 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_389_io_clk),
    .io_en(rvclkhdr_389_io_en)
  );
  rvclkhdr rvclkhdr_390 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_390_io_clk),
    .io_en(rvclkhdr_390_io_en)
  );
  rvclkhdr rvclkhdr_391 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_391_io_clk),
    .io_en(rvclkhdr_391_io_en)
  );
  rvclkhdr rvclkhdr_392 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_392_io_clk),
    .io_en(rvclkhdr_392_io_en)
  );
  rvclkhdr rvclkhdr_393 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_393_io_clk),
    .io_en(rvclkhdr_393_io_en)
  );
  rvclkhdr rvclkhdr_394 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_394_io_clk),
    .io_en(rvclkhdr_394_io_en)
  );
  rvclkhdr rvclkhdr_395 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_395_io_clk),
    .io_en(rvclkhdr_395_io_en)
  );
  rvclkhdr rvclkhdr_396 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_396_io_clk),
    .io_en(rvclkhdr_396_io_en)
  );
  rvclkhdr rvclkhdr_397 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_397_io_clk),
    .io_en(rvclkhdr_397_io_en)
  );
  rvclkhdr rvclkhdr_398 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_398_io_clk),
    .io_en(rvclkhdr_398_io_en)
  );
  rvclkhdr rvclkhdr_399 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_399_io_clk),
    .io_en(rvclkhdr_399_io_en)
  );
  rvclkhdr rvclkhdr_400 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_400_io_clk),
    .io_en(rvclkhdr_400_io_en)
  );
  rvclkhdr rvclkhdr_401 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_401_io_clk),
    .io_en(rvclkhdr_401_io_en)
  );
  rvclkhdr rvclkhdr_402 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_402_io_clk),
    .io_en(rvclkhdr_402_io_en)
  );
  rvclkhdr rvclkhdr_403 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_403_io_clk),
    .io_en(rvclkhdr_403_io_en)
  );
  rvclkhdr rvclkhdr_404 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_404_io_clk),
    .io_en(rvclkhdr_404_io_en)
  );
  rvclkhdr rvclkhdr_405 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_405_io_clk),
    .io_en(rvclkhdr_405_io_en)
  );
  rvclkhdr rvclkhdr_406 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_406_io_clk),
    .io_en(rvclkhdr_406_io_en)
  );
  rvclkhdr rvclkhdr_407 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_407_io_clk),
    .io_en(rvclkhdr_407_io_en)
  );
  rvclkhdr rvclkhdr_408 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_408_io_clk),
    .io_en(rvclkhdr_408_io_en)
  );
  rvclkhdr rvclkhdr_409 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_409_io_clk),
    .io_en(rvclkhdr_409_io_en)
  );
  rvclkhdr rvclkhdr_410 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_410_io_clk),
    .io_en(rvclkhdr_410_io_en)
  );
  rvclkhdr rvclkhdr_411 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_411_io_clk),
    .io_en(rvclkhdr_411_io_en)
  );
  rvclkhdr rvclkhdr_412 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_412_io_clk),
    .io_en(rvclkhdr_412_io_en)
  );
  rvclkhdr rvclkhdr_413 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_413_io_clk),
    .io_en(rvclkhdr_413_io_en)
  );
  rvclkhdr rvclkhdr_414 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_414_io_clk),
    .io_en(rvclkhdr_414_io_en)
  );
  rvclkhdr rvclkhdr_415 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_415_io_clk),
    .io_en(rvclkhdr_415_io_en)
  );
  rvclkhdr rvclkhdr_416 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_416_io_clk),
    .io_en(rvclkhdr_416_io_en)
  );
  rvclkhdr rvclkhdr_417 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_417_io_clk),
    .io_en(rvclkhdr_417_io_en)
  );
  rvclkhdr rvclkhdr_418 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_418_io_clk),
    .io_en(rvclkhdr_418_io_en)
  );
  rvclkhdr rvclkhdr_419 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_419_io_clk),
    .io_en(rvclkhdr_419_io_en)
  );
  rvclkhdr rvclkhdr_420 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_420_io_clk),
    .io_en(rvclkhdr_420_io_en)
  );
  rvclkhdr rvclkhdr_421 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_421_io_clk),
    .io_en(rvclkhdr_421_io_en)
  );
  rvclkhdr rvclkhdr_422 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_422_io_clk),
    .io_en(rvclkhdr_422_io_en)
  );
  rvclkhdr rvclkhdr_423 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_423_io_clk),
    .io_en(rvclkhdr_423_io_en)
  );
  rvclkhdr rvclkhdr_424 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_424_io_clk),
    .io_en(rvclkhdr_424_io_en)
  );
  rvclkhdr rvclkhdr_425 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_425_io_clk),
    .io_en(rvclkhdr_425_io_en)
  );
  rvclkhdr rvclkhdr_426 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_426_io_clk),
    .io_en(rvclkhdr_426_io_en)
  );
  rvclkhdr rvclkhdr_427 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_427_io_clk),
    .io_en(rvclkhdr_427_io_en)
  );
  rvclkhdr rvclkhdr_428 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_428_io_clk),
    .io_en(rvclkhdr_428_io_en)
  );
  rvclkhdr rvclkhdr_429 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_429_io_clk),
    .io_en(rvclkhdr_429_io_en)
  );
  rvclkhdr rvclkhdr_430 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_430_io_clk),
    .io_en(rvclkhdr_430_io_en)
  );
  rvclkhdr rvclkhdr_431 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_431_io_clk),
    .io_en(rvclkhdr_431_io_en)
  );
  rvclkhdr rvclkhdr_432 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_432_io_clk),
    .io_en(rvclkhdr_432_io_en)
  );
  rvclkhdr rvclkhdr_433 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_433_io_clk),
    .io_en(rvclkhdr_433_io_en)
  );
  rvclkhdr rvclkhdr_434 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_434_io_clk),
    .io_en(rvclkhdr_434_io_en)
  );
  rvclkhdr rvclkhdr_435 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_435_io_clk),
    .io_en(rvclkhdr_435_io_en)
  );
  rvclkhdr rvclkhdr_436 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_436_io_clk),
    .io_en(rvclkhdr_436_io_en)
  );
  rvclkhdr rvclkhdr_437 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_437_io_clk),
    .io_en(rvclkhdr_437_io_en)
  );
  rvclkhdr rvclkhdr_438 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_438_io_clk),
    .io_en(rvclkhdr_438_io_en)
  );
  rvclkhdr rvclkhdr_439 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_439_io_clk),
    .io_en(rvclkhdr_439_io_en)
  );
  rvclkhdr rvclkhdr_440 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_440_io_clk),
    .io_en(rvclkhdr_440_io_en)
  );
  rvclkhdr rvclkhdr_441 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_441_io_clk),
    .io_en(rvclkhdr_441_io_en)
  );
  rvclkhdr rvclkhdr_442 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_442_io_clk),
    .io_en(rvclkhdr_442_io_en)
  );
  rvclkhdr rvclkhdr_443 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_443_io_clk),
    .io_en(rvclkhdr_443_io_en)
  );
  rvclkhdr rvclkhdr_444 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_444_io_clk),
    .io_en(rvclkhdr_444_io_en)
  );
  rvclkhdr rvclkhdr_445 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_445_io_clk),
    .io_en(rvclkhdr_445_io_en)
  );
  rvclkhdr rvclkhdr_446 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_446_io_clk),
    .io_en(rvclkhdr_446_io_en)
  );
  rvclkhdr rvclkhdr_447 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_447_io_clk),
    .io_en(rvclkhdr_447_io_en)
  );
  rvclkhdr rvclkhdr_448 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_448_io_clk),
    .io_en(rvclkhdr_448_io_en)
  );
  rvclkhdr rvclkhdr_449 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_449_io_clk),
    .io_en(rvclkhdr_449_io_en)
  );
  rvclkhdr rvclkhdr_450 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_450_io_clk),
    .io_en(rvclkhdr_450_io_en)
  );
  rvclkhdr rvclkhdr_451 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_451_io_clk),
    .io_en(rvclkhdr_451_io_en)
  );
  rvclkhdr rvclkhdr_452 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_452_io_clk),
    .io_en(rvclkhdr_452_io_en)
  );
  rvclkhdr rvclkhdr_453 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_453_io_clk),
    .io_en(rvclkhdr_453_io_en)
  );
  rvclkhdr rvclkhdr_454 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_454_io_clk),
    .io_en(rvclkhdr_454_io_en)
  );
  rvclkhdr rvclkhdr_455 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_455_io_clk),
    .io_en(rvclkhdr_455_io_en)
  );
  rvclkhdr rvclkhdr_456 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_456_io_clk),
    .io_en(rvclkhdr_456_io_en)
  );
  rvclkhdr rvclkhdr_457 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_457_io_clk),
    .io_en(rvclkhdr_457_io_en)
  );
  rvclkhdr rvclkhdr_458 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_458_io_clk),
    .io_en(rvclkhdr_458_io_en)
  );
  rvclkhdr rvclkhdr_459 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_459_io_clk),
    .io_en(rvclkhdr_459_io_en)
  );
  rvclkhdr rvclkhdr_460 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_460_io_clk),
    .io_en(rvclkhdr_460_io_en)
  );
  rvclkhdr rvclkhdr_461 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_461_io_clk),
    .io_en(rvclkhdr_461_io_en)
  );
  rvclkhdr rvclkhdr_462 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_462_io_clk),
    .io_en(rvclkhdr_462_io_en)
  );
  rvclkhdr rvclkhdr_463 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_463_io_clk),
    .io_en(rvclkhdr_463_io_en)
  );
  rvclkhdr rvclkhdr_464 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_464_io_clk),
    .io_en(rvclkhdr_464_io_en)
  );
  rvclkhdr rvclkhdr_465 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_465_io_clk),
    .io_en(rvclkhdr_465_io_en)
  );
  rvclkhdr rvclkhdr_466 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_466_io_clk),
    .io_en(rvclkhdr_466_io_en)
  );
  rvclkhdr rvclkhdr_467 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_467_io_clk),
    .io_en(rvclkhdr_467_io_en)
  );
  rvclkhdr rvclkhdr_468 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_468_io_clk),
    .io_en(rvclkhdr_468_io_en)
  );
  rvclkhdr rvclkhdr_469 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_469_io_clk),
    .io_en(rvclkhdr_469_io_en)
  );
  rvclkhdr rvclkhdr_470 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_470_io_clk),
    .io_en(rvclkhdr_470_io_en)
  );
  rvclkhdr rvclkhdr_471 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_471_io_clk),
    .io_en(rvclkhdr_471_io_en)
  );
  rvclkhdr rvclkhdr_472 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_472_io_clk),
    .io_en(rvclkhdr_472_io_en)
  );
  rvclkhdr rvclkhdr_473 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_473_io_clk),
    .io_en(rvclkhdr_473_io_en)
  );
  rvclkhdr rvclkhdr_474 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_474_io_clk),
    .io_en(rvclkhdr_474_io_en)
  );
  rvclkhdr rvclkhdr_475 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_475_io_clk),
    .io_en(rvclkhdr_475_io_en)
  );
  rvclkhdr rvclkhdr_476 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_476_io_clk),
    .io_en(rvclkhdr_476_io_en)
  );
  rvclkhdr rvclkhdr_477 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_477_io_clk),
    .io_en(rvclkhdr_477_io_en)
  );
  rvclkhdr rvclkhdr_478 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_478_io_clk),
    .io_en(rvclkhdr_478_io_en)
  );
  rvclkhdr rvclkhdr_479 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_479_io_clk),
    .io_en(rvclkhdr_479_io_en)
  );
  rvclkhdr rvclkhdr_480 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_480_io_clk),
    .io_en(rvclkhdr_480_io_en)
  );
  rvclkhdr rvclkhdr_481 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_481_io_clk),
    .io_en(rvclkhdr_481_io_en)
  );
  rvclkhdr rvclkhdr_482 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_482_io_clk),
    .io_en(rvclkhdr_482_io_en)
  );
  rvclkhdr rvclkhdr_483 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_483_io_clk),
    .io_en(rvclkhdr_483_io_en)
  );
  rvclkhdr rvclkhdr_484 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_484_io_clk),
    .io_en(rvclkhdr_484_io_en)
  );
  rvclkhdr rvclkhdr_485 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_485_io_clk),
    .io_en(rvclkhdr_485_io_en)
  );
  rvclkhdr rvclkhdr_486 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_486_io_clk),
    .io_en(rvclkhdr_486_io_en)
  );
  rvclkhdr rvclkhdr_487 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_487_io_clk),
    .io_en(rvclkhdr_487_io_en)
  );
  rvclkhdr rvclkhdr_488 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_488_io_clk),
    .io_en(rvclkhdr_488_io_en)
  );
  rvclkhdr rvclkhdr_489 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_489_io_clk),
    .io_en(rvclkhdr_489_io_en)
  );
  rvclkhdr rvclkhdr_490 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_490_io_clk),
    .io_en(rvclkhdr_490_io_en)
  );
  rvclkhdr rvclkhdr_491 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_491_io_clk),
    .io_en(rvclkhdr_491_io_en)
  );
  rvclkhdr rvclkhdr_492 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_492_io_clk),
    .io_en(rvclkhdr_492_io_en)
  );
  rvclkhdr rvclkhdr_493 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_493_io_clk),
    .io_en(rvclkhdr_493_io_en)
  );
  rvclkhdr rvclkhdr_494 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_494_io_clk),
    .io_en(rvclkhdr_494_io_en)
  );
  rvclkhdr rvclkhdr_495 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_495_io_clk),
    .io_en(rvclkhdr_495_io_en)
  );
  rvclkhdr rvclkhdr_496 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_496_io_clk),
    .io_en(rvclkhdr_496_io_en)
  );
  rvclkhdr rvclkhdr_497 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_497_io_clk),
    .io_en(rvclkhdr_497_io_en)
  );
  rvclkhdr rvclkhdr_498 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_498_io_clk),
    .io_en(rvclkhdr_498_io_en)
  );
  rvclkhdr rvclkhdr_499 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_499_io_clk),
    .io_en(rvclkhdr_499_io_en)
  );
  rvclkhdr rvclkhdr_500 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_500_io_clk),
    .io_en(rvclkhdr_500_io_en)
  );
  rvclkhdr rvclkhdr_501 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_501_io_clk),
    .io_en(rvclkhdr_501_io_en)
  );
  rvclkhdr rvclkhdr_502 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_502_io_clk),
    .io_en(rvclkhdr_502_io_en)
  );
  rvclkhdr rvclkhdr_503 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_503_io_clk),
    .io_en(rvclkhdr_503_io_en)
  );
  rvclkhdr rvclkhdr_504 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_504_io_clk),
    .io_en(rvclkhdr_504_io_en)
  );
  rvclkhdr rvclkhdr_505 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_505_io_clk),
    .io_en(rvclkhdr_505_io_en)
  );
  rvclkhdr rvclkhdr_506 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_506_io_clk),
    .io_en(rvclkhdr_506_io_en)
  );
  rvclkhdr rvclkhdr_507 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_507_io_clk),
    .io_en(rvclkhdr_507_io_en)
  );
  rvclkhdr rvclkhdr_508 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_508_io_clk),
    .io_en(rvclkhdr_508_io_en)
  );
  rvclkhdr rvclkhdr_509 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_509_io_clk),
    .io_en(rvclkhdr_509_io_en)
  );
  rvclkhdr rvclkhdr_510 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_510_io_clk),
    .io_en(rvclkhdr_510_io_en)
  );
  rvclkhdr rvclkhdr_511 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_511_io_clk),
    .io_en(rvclkhdr_511_io_en)
  );
  rvclkhdr rvclkhdr_512 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_512_io_clk),
    .io_en(rvclkhdr_512_io_en)
  );
  rvclkhdr rvclkhdr_513 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_513_io_clk),
    .io_en(rvclkhdr_513_io_en)
  );
  rvclkhdr rvclkhdr_514 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_514_io_clk),
    .io_en(rvclkhdr_514_io_en)
  );
  rvclkhdr rvclkhdr_515 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_515_io_clk),
    .io_en(rvclkhdr_515_io_en)
  );
  rvclkhdr rvclkhdr_516 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_516_io_clk),
    .io_en(rvclkhdr_516_io_en)
  );
  rvclkhdr rvclkhdr_517 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_517_io_clk),
    .io_en(rvclkhdr_517_io_en)
  );
  rvclkhdr rvclkhdr_518 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_518_io_clk),
    .io_en(rvclkhdr_518_io_en)
  );
  rvclkhdr rvclkhdr_519 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_519_io_clk),
    .io_en(rvclkhdr_519_io_en)
  );
  rvclkhdr rvclkhdr_520 ( // @[lib.scala 409:23]
    .io_clk(rvclkhdr_520_io_clk),
    .io_en(rvclkhdr_520_io_en)
  );
  rvclkhdr rvclkhdr_521 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_521_io_clk),
    .io_en(rvclkhdr_521_io_en)
  );
  rvclkhdr rvclkhdr_522 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_522_io_clk),
    .io_en(rvclkhdr_522_io_en)
  );
  rvclkhdr rvclkhdr_523 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_523_io_clk),
    .io_en(rvclkhdr_523_io_en)
  );
  rvclkhdr rvclkhdr_524 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_524_io_clk),
    .io_en(rvclkhdr_524_io_en)
  );
  rvclkhdr rvclkhdr_525 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_525_io_clk),
    .io_en(rvclkhdr_525_io_en)
  );
  rvclkhdr rvclkhdr_526 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_526_io_clk),
    .io_en(rvclkhdr_526_io_en)
  );
  rvclkhdr rvclkhdr_527 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_527_io_clk),
    .io_en(rvclkhdr_527_io_en)
  );
  rvclkhdr rvclkhdr_528 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_528_io_clk),
    .io_en(rvclkhdr_528_io_en)
  );
  rvclkhdr rvclkhdr_529 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_529_io_clk),
    .io_en(rvclkhdr_529_io_en)
  );
  rvclkhdr rvclkhdr_530 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_530_io_clk),
    .io_en(rvclkhdr_530_io_en)
  );
  rvclkhdr rvclkhdr_531 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_531_io_clk),
    .io_en(rvclkhdr_531_io_en)
  );
  rvclkhdr rvclkhdr_532 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_532_io_clk),
    .io_en(rvclkhdr_532_io_en)
  );
  rvclkhdr rvclkhdr_533 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_533_io_clk),
    .io_en(rvclkhdr_533_io_en)
  );
  rvclkhdr rvclkhdr_534 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_534_io_clk),
    .io_en(rvclkhdr_534_io_en)
  );
  rvclkhdr rvclkhdr_535 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_535_io_clk),
    .io_en(rvclkhdr_535_io_en)
  );
  rvclkhdr rvclkhdr_536 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_536_io_clk),
    .io_en(rvclkhdr_536_io_en)
  );
  rvclkhdr rvclkhdr_537 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_537_io_clk),
    .io_en(rvclkhdr_537_io_en)
  );
  rvclkhdr rvclkhdr_538 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_538_io_clk),
    .io_en(rvclkhdr_538_io_en)
  );
  rvclkhdr rvclkhdr_539 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_539_io_clk),
    .io_en(rvclkhdr_539_io_en)
  );
  rvclkhdr rvclkhdr_540 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_540_io_clk),
    .io_en(rvclkhdr_540_io_en)
  );
  rvclkhdr rvclkhdr_541 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_541_io_clk),
    .io_en(rvclkhdr_541_io_en)
  );
  rvclkhdr rvclkhdr_542 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_542_io_clk),
    .io_en(rvclkhdr_542_io_en)
  );
  rvclkhdr rvclkhdr_543 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_543_io_clk),
    .io_en(rvclkhdr_543_io_en)
  );
  rvclkhdr rvclkhdr_544 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_544_io_clk),
    .io_en(rvclkhdr_544_io_en)
  );
  rvclkhdr rvclkhdr_545 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_545_io_clk),
    .io_en(rvclkhdr_545_io_en)
  );
  rvclkhdr rvclkhdr_546 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_546_io_clk),
    .io_en(rvclkhdr_546_io_en)
  );
  rvclkhdr rvclkhdr_547 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_547_io_clk),
    .io_en(rvclkhdr_547_io_en)
  );
  rvclkhdr rvclkhdr_548 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_548_io_clk),
    .io_en(rvclkhdr_548_io_en)
  );
  rvclkhdr rvclkhdr_549 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_549_io_clk),
    .io_en(rvclkhdr_549_io_en)
  );
  rvclkhdr rvclkhdr_550 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_550_io_clk),
    .io_en(rvclkhdr_550_io_en)
  );
  rvclkhdr rvclkhdr_551 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_551_io_clk),
    .io_en(rvclkhdr_551_io_en)
  );
  rvclkhdr rvclkhdr_552 ( // @[lib.scala 343:22]
    .io_clk(rvclkhdr_552_io_clk),
    .io_en(rvclkhdr_552_io_en)
  );
  assign io_ifu_bp_hit_taken_f = _T_231 & _T_232; // @[ifu_bp_ctl.scala 277:25]
  assign io_ifu_bp_btb_target_f = _T_443 | _T_453; // @[ifu_bp_ctl.scala 374:26]
  assign io_ifu_bp_inst_mask_f = _T_268 | _T_269; // @[ifu_bp_ctl.scala 302:25]
  assign io_ifu_bp_fghr_f = fghr; // @[ifu_bp_ctl.scala 345:20]
  assign io_ifu_bp_way_f = tag_match_vway1_expanded_f | _T_154; // @[ifu_bp_ctl.scala 254:19]
  assign io_ifu_bp_ret_f = {_T_288,_T_294}; // @[ifu_bp_ctl.scala 351:19]
  assign io_ifu_bp_hist1_f = bht_force_taken_f | _T_273; // @[ifu_bp_ctl.scala 346:21]
  assign io_ifu_bp_hist0_f = {bht_vbank1_rd_data_f[0],bht_vbank0_rd_data_f[0]}; // @[ifu_bp_ctl.scala 347:21]
  assign io_ifu_bp_pc4_f = {_T_279,_T_282}; // @[ifu_bp_ctl.scala 348:19]
  assign io_ifu_bp_valid_f = vwayhit_f & _T_353; // @[ifu_bp_ctl.scala 350:21]
  assign io_ifu_bp_poffset_f = btb_sel_data_f[15:4]; // @[ifu_bp_ctl.scala 362:23]
  assign io_ifu_bp_fa_index_f_0 = 9'h0; // @[ifu_bp_ctl.scala 35:24]
  assign io_ifu_bp_fa_index_f_1 = 9'h0; // @[ifu_bp_ctl.scala 35:24]
  assign rvclkhdr_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_io_en = io_ifc_fetch_req_f | exu_mp_valid; // @[lib.scala 412:17]
  assign rvclkhdr_1_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_1_io_en = ~rs_hold; // @[lib.scala 412:17]
  assign rvclkhdr_2_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_2_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_3_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_3_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_4_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_4_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_5_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_5_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_6_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_6_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_7_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_7_io_en = rs_push | rs_pop; // @[lib.scala 412:17]
  assign rvclkhdr_8_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_8_io_en = _T_494 & io_ifu_bp_hit_taken_f; // @[lib.scala 412:17]
  assign rvclkhdr_9_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_9_io_en = _T_613 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_10_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_10_io_en = _T_617 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_11_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_11_io_en = _T_621 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_12_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_12_io_en = _T_625 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_13_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_13_io_en = _T_629 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_14_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_14_io_en = _T_633 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_15_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_15_io_en = _T_637 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_16_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_16_io_en = _T_641 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_17_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_17_io_en = _T_645 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_18_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_18_io_en = _T_649 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_19_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_19_io_en = _T_653 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_20_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_20_io_en = _T_657 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_21_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_21_io_en = _T_661 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_22_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_22_io_en = _T_665 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_23_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_23_io_en = _T_669 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_24_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_24_io_en = _T_673 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_25_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_25_io_en = _T_677 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_26_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_26_io_en = _T_681 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_27_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_27_io_en = _T_685 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_28_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_28_io_en = _T_689 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_29_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_29_io_en = _T_693 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_30_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_30_io_en = _T_697 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_31_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_31_io_en = _T_701 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_32_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_32_io_en = _T_705 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_33_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_33_io_en = _T_709 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_34_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_34_io_en = _T_713 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_35_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_35_io_en = _T_717 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_36_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_36_io_en = _T_721 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_37_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_37_io_en = _T_725 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_38_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_38_io_en = _T_729 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_39_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_39_io_en = _T_733 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_40_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_40_io_en = _T_737 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_41_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_41_io_en = _T_741 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_42_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_42_io_en = _T_745 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_43_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_43_io_en = _T_749 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_44_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_44_io_en = _T_753 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_45_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_45_io_en = _T_757 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_46_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_46_io_en = _T_761 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_47_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_47_io_en = _T_765 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_48_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_48_io_en = _T_769 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_49_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_49_io_en = _T_773 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_50_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_50_io_en = _T_777 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_51_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_51_io_en = _T_781 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_52_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_52_io_en = _T_785 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_53_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_53_io_en = _T_789 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_54_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_54_io_en = _T_793 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_55_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_55_io_en = _T_797 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_56_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_56_io_en = _T_801 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_57_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_57_io_en = _T_805 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_58_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_58_io_en = _T_809 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_59_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_59_io_en = _T_813 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_60_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_60_io_en = _T_817 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_61_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_61_io_en = _T_821 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_62_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_62_io_en = _T_825 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_63_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_63_io_en = _T_829 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_64_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_64_io_en = _T_833 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_65_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_65_io_en = _T_837 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_66_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_66_io_en = _T_841 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_67_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_67_io_en = _T_845 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_68_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_68_io_en = _T_849 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_69_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_69_io_en = _T_853 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_70_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_70_io_en = _T_857 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_71_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_71_io_en = _T_861 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_72_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_72_io_en = _T_865 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_73_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_73_io_en = _T_869 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_74_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_74_io_en = _T_873 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_75_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_75_io_en = _T_877 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_76_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_76_io_en = _T_881 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_77_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_77_io_en = _T_885 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_78_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_78_io_en = _T_889 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_79_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_79_io_en = _T_893 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_80_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_80_io_en = _T_897 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_81_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_81_io_en = _T_901 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_82_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_82_io_en = _T_905 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_83_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_83_io_en = _T_909 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_84_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_84_io_en = _T_913 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_85_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_85_io_en = _T_917 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_86_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_86_io_en = _T_921 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_87_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_87_io_en = _T_925 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_88_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_88_io_en = _T_929 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_89_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_89_io_en = _T_933 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_90_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_90_io_en = _T_937 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_91_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_91_io_en = _T_941 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_92_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_92_io_en = _T_945 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_93_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_93_io_en = _T_949 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_94_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_94_io_en = _T_953 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_95_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_95_io_en = _T_957 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_96_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_96_io_en = _T_961 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_97_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_97_io_en = _T_965 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_98_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_98_io_en = _T_969 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_99_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_99_io_en = _T_973 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_100_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_100_io_en = _T_977 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_101_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_101_io_en = _T_981 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_102_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_102_io_en = _T_985 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_103_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_103_io_en = _T_989 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_104_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_104_io_en = _T_993 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_105_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_105_io_en = _T_997 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_106_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_106_io_en = _T_1001 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_107_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_107_io_en = _T_1005 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_108_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_108_io_en = _T_1009 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_109_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_109_io_en = _T_1013 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_110_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_110_io_en = _T_1017 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_111_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_111_io_en = _T_1021 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_112_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_112_io_en = _T_1025 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_113_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_113_io_en = _T_1029 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_114_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_114_io_en = _T_1033 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_115_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_115_io_en = _T_1037 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_116_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_116_io_en = _T_1041 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_117_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_117_io_en = _T_1045 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_118_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_118_io_en = _T_1049 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_119_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_119_io_en = _T_1053 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_120_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_120_io_en = _T_1057 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_121_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_121_io_en = _T_1061 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_122_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_122_io_en = _T_1065 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_123_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_123_io_en = _T_1069 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_124_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_124_io_en = _T_1073 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_125_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_125_io_en = _T_1077 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_126_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_126_io_en = _T_1081 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_127_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_127_io_en = _T_1085 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_128_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_128_io_en = _T_1089 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_129_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_129_io_en = _T_1093 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_130_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_130_io_en = _T_1097 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_131_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_131_io_en = _T_1101 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_132_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_132_io_en = _T_1105 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_133_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_133_io_en = _T_1109 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_134_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_134_io_en = _T_1113 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_135_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_135_io_en = _T_1117 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_136_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_136_io_en = _T_1121 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_137_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_137_io_en = _T_1125 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_138_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_138_io_en = _T_1129 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_139_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_139_io_en = _T_1133 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_140_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_140_io_en = _T_1137 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_141_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_141_io_en = _T_1141 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_142_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_142_io_en = _T_1145 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_143_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_143_io_en = _T_1149 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_144_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_144_io_en = _T_1153 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_145_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_145_io_en = _T_1157 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_146_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_146_io_en = _T_1161 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_147_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_147_io_en = _T_1165 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_148_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_148_io_en = _T_1169 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_149_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_149_io_en = _T_1173 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_150_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_150_io_en = _T_1177 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_151_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_151_io_en = _T_1181 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_152_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_152_io_en = _T_1185 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_153_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_153_io_en = _T_1189 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_154_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_154_io_en = _T_1193 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_155_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_155_io_en = _T_1197 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_156_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_156_io_en = _T_1201 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_157_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_157_io_en = _T_1205 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_158_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_158_io_en = _T_1209 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_159_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_159_io_en = _T_1213 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_160_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_160_io_en = _T_1217 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_161_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_161_io_en = _T_1221 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_162_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_162_io_en = _T_1225 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_163_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_163_io_en = _T_1229 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_164_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_164_io_en = _T_1233 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_165_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_165_io_en = _T_1237 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_166_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_166_io_en = _T_1241 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_167_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_167_io_en = _T_1245 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_168_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_168_io_en = _T_1249 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_169_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_169_io_en = _T_1253 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_170_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_170_io_en = _T_1257 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_171_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_171_io_en = _T_1261 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_172_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_172_io_en = _T_1265 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_173_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_173_io_en = _T_1269 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_174_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_174_io_en = _T_1273 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_175_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_175_io_en = _T_1277 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_176_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_176_io_en = _T_1281 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_177_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_177_io_en = _T_1285 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_178_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_178_io_en = _T_1289 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_179_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_179_io_en = _T_1293 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_180_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_180_io_en = _T_1297 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_181_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_181_io_en = _T_1301 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_182_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_182_io_en = _T_1305 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_183_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_183_io_en = _T_1309 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_184_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_184_io_en = _T_1313 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_185_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_185_io_en = _T_1317 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_186_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_186_io_en = _T_1321 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_187_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_187_io_en = _T_1325 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_188_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_188_io_en = _T_1329 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_189_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_189_io_en = _T_1333 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_190_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_190_io_en = _T_1337 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_191_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_191_io_en = _T_1341 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_192_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_192_io_en = _T_1345 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_193_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_193_io_en = _T_1349 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_194_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_194_io_en = _T_1353 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_195_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_195_io_en = _T_1357 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_196_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_196_io_en = _T_1361 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_197_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_197_io_en = _T_1365 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_198_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_198_io_en = _T_1369 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_199_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_199_io_en = _T_1373 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_200_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_200_io_en = _T_1377 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_201_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_201_io_en = _T_1381 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_202_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_202_io_en = _T_1385 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_203_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_203_io_en = _T_1389 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_204_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_204_io_en = _T_1393 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_205_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_205_io_en = _T_1397 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_206_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_206_io_en = _T_1401 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_207_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_207_io_en = _T_1405 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_208_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_208_io_en = _T_1409 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_209_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_209_io_en = _T_1413 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_210_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_210_io_en = _T_1417 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_211_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_211_io_en = _T_1421 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_212_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_212_io_en = _T_1425 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_213_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_213_io_en = _T_1429 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_214_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_214_io_en = _T_1433 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_215_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_215_io_en = _T_1437 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_216_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_216_io_en = _T_1441 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_217_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_217_io_en = _T_1445 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_218_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_218_io_en = _T_1449 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_219_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_219_io_en = _T_1453 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_220_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_220_io_en = _T_1457 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_221_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_221_io_en = _T_1461 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_222_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_222_io_en = _T_1465 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_223_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_223_io_en = _T_1469 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_224_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_224_io_en = _T_1473 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_225_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_225_io_en = _T_1477 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_226_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_226_io_en = _T_1481 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_227_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_227_io_en = _T_1485 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_228_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_228_io_en = _T_1489 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_229_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_229_io_en = _T_1493 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_230_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_230_io_en = _T_1497 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_231_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_231_io_en = _T_1501 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_232_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_232_io_en = _T_1505 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_233_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_233_io_en = _T_1509 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_234_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_234_io_en = _T_1513 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_235_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_235_io_en = _T_1517 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_236_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_236_io_en = _T_1521 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_237_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_237_io_en = _T_1525 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_238_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_238_io_en = _T_1529 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_239_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_239_io_en = _T_1533 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_240_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_240_io_en = _T_1537 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_241_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_241_io_en = _T_1541 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_242_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_242_io_en = _T_1545 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_243_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_243_io_en = _T_1549 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_244_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_244_io_en = _T_1553 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_245_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_245_io_en = _T_1557 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_246_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_246_io_en = _T_1561 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_247_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_247_io_en = _T_1565 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_248_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_248_io_en = _T_1569 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_249_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_249_io_en = _T_1573 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_250_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_250_io_en = _T_1577 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_251_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_251_io_en = _T_1581 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_252_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_252_io_en = _T_1585 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_253_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_253_io_en = _T_1589 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_254_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_254_io_en = _T_1593 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_255_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_255_io_en = _T_1597 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_256_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_256_io_en = _T_1601 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_257_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_257_io_en = _T_1605 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_258_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_258_io_en = _T_1609 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_259_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_259_io_en = _T_1613 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_260_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_260_io_en = _T_1617 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_261_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_261_io_en = _T_1621 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_262_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_262_io_en = _T_1625 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_263_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_263_io_en = _T_1629 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_264_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_264_io_en = _T_1633 & btb_wr_en_way0; // @[lib.scala 412:17]
  assign rvclkhdr_265_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_265_io_en = _T_613 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_266_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_266_io_en = _T_617 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_267_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_267_io_en = _T_621 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_268_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_268_io_en = _T_625 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_269_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_269_io_en = _T_629 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_270_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_270_io_en = _T_633 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_271_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_271_io_en = _T_637 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_272_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_272_io_en = _T_641 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_273_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_273_io_en = _T_645 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_274_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_274_io_en = _T_649 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_275_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_275_io_en = _T_653 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_276_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_276_io_en = _T_657 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_277_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_277_io_en = _T_661 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_278_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_278_io_en = _T_665 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_279_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_279_io_en = _T_669 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_280_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_280_io_en = _T_673 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_281_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_281_io_en = _T_677 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_282_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_282_io_en = _T_681 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_283_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_283_io_en = _T_685 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_284_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_284_io_en = _T_689 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_285_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_285_io_en = _T_693 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_286_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_286_io_en = _T_697 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_287_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_287_io_en = _T_701 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_288_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_288_io_en = _T_705 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_289_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_289_io_en = _T_709 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_290_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_290_io_en = _T_713 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_291_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_291_io_en = _T_717 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_292_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_292_io_en = _T_721 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_293_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_293_io_en = _T_725 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_294_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_294_io_en = _T_729 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_295_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_295_io_en = _T_733 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_296_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_296_io_en = _T_737 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_297_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_297_io_en = _T_741 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_298_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_298_io_en = _T_745 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_299_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_299_io_en = _T_749 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_300_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_300_io_en = _T_753 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_301_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_301_io_en = _T_757 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_302_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_302_io_en = _T_761 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_303_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_303_io_en = _T_765 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_304_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_304_io_en = _T_769 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_305_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_305_io_en = _T_773 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_306_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_306_io_en = _T_777 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_307_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_307_io_en = _T_781 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_308_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_308_io_en = _T_785 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_309_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_309_io_en = _T_789 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_310_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_310_io_en = _T_793 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_311_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_311_io_en = _T_797 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_312_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_312_io_en = _T_801 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_313_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_313_io_en = _T_805 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_314_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_314_io_en = _T_809 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_315_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_315_io_en = _T_813 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_316_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_316_io_en = _T_817 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_317_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_317_io_en = _T_821 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_318_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_318_io_en = _T_825 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_319_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_319_io_en = _T_829 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_320_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_320_io_en = _T_833 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_321_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_321_io_en = _T_837 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_322_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_322_io_en = _T_841 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_323_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_323_io_en = _T_845 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_324_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_324_io_en = _T_849 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_325_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_325_io_en = _T_853 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_326_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_326_io_en = _T_857 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_327_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_327_io_en = _T_861 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_328_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_328_io_en = _T_865 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_329_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_329_io_en = _T_869 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_330_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_330_io_en = _T_873 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_331_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_331_io_en = _T_877 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_332_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_332_io_en = _T_881 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_333_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_333_io_en = _T_885 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_334_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_334_io_en = _T_889 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_335_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_335_io_en = _T_893 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_336_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_336_io_en = _T_897 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_337_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_337_io_en = _T_901 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_338_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_338_io_en = _T_905 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_339_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_339_io_en = _T_909 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_340_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_340_io_en = _T_913 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_341_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_341_io_en = _T_917 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_342_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_342_io_en = _T_921 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_343_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_343_io_en = _T_925 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_344_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_344_io_en = _T_929 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_345_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_345_io_en = _T_933 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_346_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_346_io_en = _T_937 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_347_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_347_io_en = _T_941 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_348_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_348_io_en = _T_945 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_349_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_349_io_en = _T_949 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_350_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_350_io_en = _T_953 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_351_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_351_io_en = _T_957 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_352_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_352_io_en = _T_961 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_353_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_353_io_en = _T_965 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_354_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_354_io_en = _T_969 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_355_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_355_io_en = _T_973 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_356_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_356_io_en = _T_977 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_357_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_357_io_en = _T_981 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_358_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_358_io_en = _T_985 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_359_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_359_io_en = _T_989 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_360_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_360_io_en = _T_993 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_361_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_361_io_en = _T_997 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_362_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_362_io_en = _T_1001 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_363_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_363_io_en = _T_1005 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_364_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_364_io_en = _T_1009 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_365_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_365_io_en = _T_1013 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_366_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_366_io_en = _T_1017 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_367_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_367_io_en = _T_1021 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_368_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_368_io_en = _T_1025 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_369_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_369_io_en = _T_1029 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_370_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_370_io_en = _T_1033 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_371_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_371_io_en = _T_1037 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_372_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_372_io_en = _T_1041 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_373_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_373_io_en = _T_1045 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_374_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_374_io_en = _T_1049 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_375_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_375_io_en = _T_1053 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_376_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_376_io_en = _T_1057 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_377_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_377_io_en = _T_1061 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_378_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_378_io_en = _T_1065 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_379_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_379_io_en = _T_1069 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_380_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_380_io_en = _T_1073 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_381_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_381_io_en = _T_1077 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_382_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_382_io_en = _T_1081 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_383_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_383_io_en = _T_1085 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_384_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_384_io_en = _T_1089 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_385_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_385_io_en = _T_1093 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_386_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_386_io_en = _T_1097 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_387_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_387_io_en = _T_1101 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_388_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_388_io_en = _T_1105 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_389_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_389_io_en = _T_1109 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_390_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_390_io_en = _T_1113 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_391_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_391_io_en = _T_1117 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_392_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_392_io_en = _T_1121 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_393_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_393_io_en = _T_1125 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_394_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_394_io_en = _T_1129 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_395_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_395_io_en = _T_1133 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_396_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_396_io_en = _T_1137 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_397_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_397_io_en = _T_1141 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_398_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_398_io_en = _T_1145 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_399_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_399_io_en = _T_1149 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_400_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_400_io_en = _T_1153 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_401_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_401_io_en = _T_1157 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_402_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_402_io_en = _T_1161 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_403_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_403_io_en = _T_1165 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_404_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_404_io_en = _T_1169 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_405_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_405_io_en = _T_1173 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_406_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_406_io_en = _T_1177 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_407_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_407_io_en = _T_1181 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_408_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_408_io_en = _T_1185 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_409_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_409_io_en = _T_1189 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_410_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_410_io_en = _T_1193 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_411_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_411_io_en = _T_1197 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_412_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_412_io_en = _T_1201 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_413_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_413_io_en = _T_1205 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_414_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_414_io_en = _T_1209 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_415_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_415_io_en = _T_1213 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_416_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_416_io_en = _T_1217 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_417_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_417_io_en = _T_1221 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_418_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_418_io_en = _T_1225 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_419_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_419_io_en = _T_1229 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_420_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_420_io_en = _T_1233 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_421_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_421_io_en = _T_1237 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_422_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_422_io_en = _T_1241 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_423_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_423_io_en = _T_1245 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_424_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_424_io_en = _T_1249 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_425_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_425_io_en = _T_1253 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_426_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_426_io_en = _T_1257 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_427_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_427_io_en = _T_1261 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_428_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_428_io_en = _T_1265 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_429_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_429_io_en = _T_1269 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_430_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_430_io_en = _T_1273 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_431_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_431_io_en = _T_1277 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_432_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_432_io_en = _T_1281 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_433_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_433_io_en = _T_1285 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_434_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_434_io_en = _T_1289 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_435_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_435_io_en = _T_1293 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_436_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_436_io_en = _T_1297 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_437_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_437_io_en = _T_1301 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_438_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_438_io_en = _T_1305 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_439_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_439_io_en = _T_1309 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_440_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_440_io_en = _T_1313 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_441_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_441_io_en = _T_1317 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_442_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_442_io_en = _T_1321 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_443_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_443_io_en = _T_1325 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_444_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_444_io_en = _T_1329 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_445_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_445_io_en = _T_1333 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_446_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_446_io_en = _T_1337 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_447_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_447_io_en = _T_1341 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_448_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_448_io_en = _T_1345 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_449_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_449_io_en = _T_1349 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_450_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_450_io_en = _T_1353 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_451_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_451_io_en = _T_1357 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_452_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_452_io_en = _T_1361 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_453_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_453_io_en = _T_1365 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_454_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_454_io_en = _T_1369 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_455_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_455_io_en = _T_1373 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_456_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_456_io_en = _T_1377 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_457_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_457_io_en = _T_1381 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_458_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_458_io_en = _T_1385 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_459_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_459_io_en = _T_1389 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_460_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_460_io_en = _T_1393 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_461_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_461_io_en = _T_1397 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_462_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_462_io_en = _T_1401 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_463_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_463_io_en = _T_1405 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_464_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_464_io_en = _T_1409 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_465_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_465_io_en = _T_1413 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_466_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_466_io_en = _T_1417 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_467_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_467_io_en = _T_1421 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_468_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_468_io_en = _T_1425 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_469_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_469_io_en = _T_1429 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_470_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_470_io_en = _T_1433 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_471_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_471_io_en = _T_1437 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_472_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_472_io_en = _T_1441 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_473_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_473_io_en = _T_1445 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_474_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_474_io_en = _T_1449 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_475_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_475_io_en = _T_1453 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_476_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_476_io_en = _T_1457 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_477_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_477_io_en = _T_1461 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_478_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_478_io_en = _T_1465 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_479_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_479_io_en = _T_1469 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_480_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_480_io_en = _T_1473 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_481_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_481_io_en = _T_1477 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_482_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_482_io_en = _T_1481 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_483_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_483_io_en = _T_1485 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_484_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_484_io_en = _T_1489 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_485_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_485_io_en = _T_1493 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_486_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_486_io_en = _T_1497 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_487_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_487_io_en = _T_1501 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_488_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_488_io_en = _T_1505 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_489_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_489_io_en = _T_1509 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_490_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_490_io_en = _T_1513 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_491_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_491_io_en = _T_1517 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_492_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_492_io_en = _T_1521 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_493_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_493_io_en = _T_1525 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_494_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_494_io_en = _T_1529 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_495_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_495_io_en = _T_1533 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_496_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_496_io_en = _T_1537 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_497_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_497_io_en = _T_1541 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_498_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_498_io_en = _T_1545 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_499_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_499_io_en = _T_1549 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_500_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_500_io_en = _T_1553 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_501_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_501_io_en = _T_1557 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_502_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_502_io_en = _T_1561 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_503_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_503_io_en = _T_1565 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_504_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_504_io_en = _T_1569 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_505_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_505_io_en = _T_1573 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_506_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_506_io_en = _T_1577 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_507_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_507_io_en = _T_1581 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_508_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_508_io_en = _T_1585 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_509_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_509_io_en = _T_1589 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_510_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_510_io_en = _T_1593 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_511_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_511_io_en = _T_1597 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_512_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_512_io_en = _T_1601 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_513_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_513_io_en = _T_1605 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_514_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_514_io_en = _T_1609 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_515_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_515_io_en = _T_1613 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_516_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_516_io_en = _T_1617 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_517_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_517_io_en = _T_1621 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_518_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_518_io_en = _T_1625 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_519_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_519_io_en = _T_1629 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_520_io_clk = clock; // @[lib.scala 411:18]
  assign rvclkhdr_520_io_en = _T_1633 & btb_wr_en_way1; // @[lib.scala 412:17]
  assign rvclkhdr_521_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_521_io_en = _T_6761 | _T_6766; // @[lib.scala 345:16]
  assign rvclkhdr_522_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_522_io_en = _T_6772 | _T_6777; // @[lib.scala 345:16]
  assign rvclkhdr_523_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_523_io_en = _T_6783 | _T_6788; // @[lib.scala 345:16]
  assign rvclkhdr_524_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_524_io_en = _T_6794 | _T_6799; // @[lib.scala 345:16]
  assign rvclkhdr_525_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_525_io_en = _T_6805 | _T_6810; // @[lib.scala 345:16]
  assign rvclkhdr_526_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_526_io_en = _T_6816 | _T_6821; // @[lib.scala 345:16]
  assign rvclkhdr_527_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_527_io_en = _T_6827 | _T_6832; // @[lib.scala 345:16]
  assign rvclkhdr_528_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_528_io_en = _T_6838 | _T_6843; // @[lib.scala 345:16]
  assign rvclkhdr_529_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_529_io_en = _T_6849 | _T_6854; // @[lib.scala 345:16]
  assign rvclkhdr_530_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_530_io_en = _T_6860 | _T_6865; // @[lib.scala 345:16]
  assign rvclkhdr_531_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_531_io_en = _T_6871 | _T_6876; // @[lib.scala 345:16]
  assign rvclkhdr_532_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_532_io_en = _T_6882 | _T_6887; // @[lib.scala 345:16]
  assign rvclkhdr_533_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_533_io_en = _T_6893 | _T_6898; // @[lib.scala 345:16]
  assign rvclkhdr_534_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_534_io_en = _T_6904 | _T_6909; // @[lib.scala 345:16]
  assign rvclkhdr_535_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_535_io_en = _T_6915 | _T_6920; // @[lib.scala 345:16]
  assign rvclkhdr_536_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_536_io_en = _T_6926 | _T_6931; // @[lib.scala 345:16]
  assign rvclkhdr_537_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_537_io_en = _T_6937 | _T_6942; // @[lib.scala 345:16]
  assign rvclkhdr_538_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_538_io_en = _T_6948 | _T_6953; // @[lib.scala 345:16]
  assign rvclkhdr_539_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_539_io_en = _T_6959 | _T_6964; // @[lib.scala 345:16]
  assign rvclkhdr_540_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_540_io_en = _T_6970 | _T_6975; // @[lib.scala 345:16]
  assign rvclkhdr_541_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_541_io_en = _T_6981 | _T_6986; // @[lib.scala 345:16]
  assign rvclkhdr_542_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_542_io_en = _T_6992 | _T_6997; // @[lib.scala 345:16]
  assign rvclkhdr_543_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_543_io_en = _T_7003 | _T_7008; // @[lib.scala 345:16]
  assign rvclkhdr_544_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_544_io_en = _T_7014 | _T_7019; // @[lib.scala 345:16]
  assign rvclkhdr_545_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_545_io_en = _T_7025 | _T_7030; // @[lib.scala 345:16]
  assign rvclkhdr_546_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_546_io_en = _T_7036 | _T_7041; // @[lib.scala 345:16]
  assign rvclkhdr_547_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_547_io_en = _T_7047 | _T_7052; // @[lib.scala 345:16]
  assign rvclkhdr_548_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_548_io_en = _T_7058 | _T_7063; // @[lib.scala 345:16]
  assign rvclkhdr_549_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_549_io_en = _T_7069 | _T_7074; // @[lib.scala 345:16]
  assign rvclkhdr_550_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_550_io_en = _T_7080 | _T_7085; // @[lib.scala 345:16]
  assign rvclkhdr_551_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_551_io_en = _T_7091 | _T_7096; // @[lib.scala 345:16]
  assign rvclkhdr_552_io_clk = clock; // @[lib.scala 344:17]
  assign rvclkhdr_552_io_en = _T_7102 | _T_7107; // @[lib.scala 345:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  leak_one_f_d1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_0 = _RAND_1[21:0];
  _RAND_2 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_1 = _RAND_2[21:0];
  _RAND_3 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_2 = _RAND_3[21:0];
  _RAND_4 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_3 = _RAND_4[21:0];
  _RAND_5 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_4 = _RAND_5[21:0];
  _RAND_6 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_5 = _RAND_6[21:0];
  _RAND_7 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_6 = _RAND_7[21:0];
  _RAND_8 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_7 = _RAND_8[21:0];
  _RAND_9 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_8 = _RAND_9[21:0];
  _RAND_10 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_9 = _RAND_10[21:0];
  _RAND_11 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_10 = _RAND_11[21:0];
  _RAND_12 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_11 = _RAND_12[21:0];
  _RAND_13 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_12 = _RAND_13[21:0];
  _RAND_14 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_13 = _RAND_14[21:0];
  _RAND_15 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_14 = _RAND_15[21:0];
  _RAND_16 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_15 = _RAND_16[21:0];
  _RAND_17 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_16 = _RAND_17[21:0];
  _RAND_18 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_17 = _RAND_18[21:0];
  _RAND_19 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_18 = _RAND_19[21:0];
  _RAND_20 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_19 = _RAND_20[21:0];
  _RAND_21 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_20 = _RAND_21[21:0];
  _RAND_22 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_21 = _RAND_22[21:0];
  _RAND_23 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_22 = _RAND_23[21:0];
  _RAND_24 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_23 = _RAND_24[21:0];
  _RAND_25 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_24 = _RAND_25[21:0];
  _RAND_26 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_25 = _RAND_26[21:0];
  _RAND_27 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_26 = _RAND_27[21:0];
  _RAND_28 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_27 = _RAND_28[21:0];
  _RAND_29 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_28 = _RAND_29[21:0];
  _RAND_30 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_29 = _RAND_30[21:0];
  _RAND_31 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_30 = _RAND_31[21:0];
  _RAND_32 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_31 = _RAND_32[21:0];
  _RAND_33 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_32 = _RAND_33[21:0];
  _RAND_34 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_33 = _RAND_34[21:0];
  _RAND_35 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_34 = _RAND_35[21:0];
  _RAND_36 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_35 = _RAND_36[21:0];
  _RAND_37 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_36 = _RAND_37[21:0];
  _RAND_38 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_37 = _RAND_38[21:0];
  _RAND_39 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_38 = _RAND_39[21:0];
  _RAND_40 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_39 = _RAND_40[21:0];
  _RAND_41 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_40 = _RAND_41[21:0];
  _RAND_42 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_41 = _RAND_42[21:0];
  _RAND_43 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_42 = _RAND_43[21:0];
  _RAND_44 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_43 = _RAND_44[21:0];
  _RAND_45 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_44 = _RAND_45[21:0];
  _RAND_46 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_45 = _RAND_46[21:0];
  _RAND_47 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_46 = _RAND_47[21:0];
  _RAND_48 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_47 = _RAND_48[21:0];
  _RAND_49 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_48 = _RAND_49[21:0];
  _RAND_50 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_49 = _RAND_50[21:0];
  _RAND_51 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_50 = _RAND_51[21:0];
  _RAND_52 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_51 = _RAND_52[21:0];
  _RAND_53 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_52 = _RAND_53[21:0];
  _RAND_54 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_53 = _RAND_54[21:0];
  _RAND_55 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_54 = _RAND_55[21:0];
  _RAND_56 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_55 = _RAND_56[21:0];
  _RAND_57 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_56 = _RAND_57[21:0];
  _RAND_58 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_57 = _RAND_58[21:0];
  _RAND_59 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_58 = _RAND_59[21:0];
  _RAND_60 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_59 = _RAND_60[21:0];
  _RAND_61 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_60 = _RAND_61[21:0];
  _RAND_62 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_61 = _RAND_62[21:0];
  _RAND_63 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_62 = _RAND_63[21:0];
  _RAND_64 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_63 = _RAND_64[21:0];
  _RAND_65 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_64 = _RAND_65[21:0];
  _RAND_66 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_65 = _RAND_66[21:0];
  _RAND_67 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_66 = _RAND_67[21:0];
  _RAND_68 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_67 = _RAND_68[21:0];
  _RAND_69 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_68 = _RAND_69[21:0];
  _RAND_70 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_69 = _RAND_70[21:0];
  _RAND_71 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_70 = _RAND_71[21:0];
  _RAND_72 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_71 = _RAND_72[21:0];
  _RAND_73 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_72 = _RAND_73[21:0];
  _RAND_74 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_73 = _RAND_74[21:0];
  _RAND_75 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_74 = _RAND_75[21:0];
  _RAND_76 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_75 = _RAND_76[21:0];
  _RAND_77 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_76 = _RAND_77[21:0];
  _RAND_78 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_77 = _RAND_78[21:0];
  _RAND_79 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_78 = _RAND_79[21:0];
  _RAND_80 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_79 = _RAND_80[21:0];
  _RAND_81 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_80 = _RAND_81[21:0];
  _RAND_82 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_81 = _RAND_82[21:0];
  _RAND_83 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_82 = _RAND_83[21:0];
  _RAND_84 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_83 = _RAND_84[21:0];
  _RAND_85 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_84 = _RAND_85[21:0];
  _RAND_86 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_85 = _RAND_86[21:0];
  _RAND_87 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_86 = _RAND_87[21:0];
  _RAND_88 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_87 = _RAND_88[21:0];
  _RAND_89 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_88 = _RAND_89[21:0];
  _RAND_90 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_89 = _RAND_90[21:0];
  _RAND_91 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_90 = _RAND_91[21:0];
  _RAND_92 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_91 = _RAND_92[21:0];
  _RAND_93 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_92 = _RAND_93[21:0];
  _RAND_94 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_93 = _RAND_94[21:0];
  _RAND_95 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_94 = _RAND_95[21:0];
  _RAND_96 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_95 = _RAND_96[21:0];
  _RAND_97 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_96 = _RAND_97[21:0];
  _RAND_98 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_97 = _RAND_98[21:0];
  _RAND_99 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_98 = _RAND_99[21:0];
  _RAND_100 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_99 = _RAND_100[21:0];
  _RAND_101 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_100 = _RAND_101[21:0];
  _RAND_102 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_101 = _RAND_102[21:0];
  _RAND_103 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_102 = _RAND_103[21:0];
  _RAND_104 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_103 = _RAND_104[21:0];
  _RAND_105 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_104 = _RAND_105[21:0];
  _RAND_106 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_105 = _RAND_106[21:0];
  _RAND_107 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_106 = _RAND_107[21:0];
  _RAND_108 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_107 = _RAND_108[21:0];
  _RAND_109 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_108 = _RAND_109[21:0];
  _RAND_110 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_109 = _RAND_110[21:0];
  _RAND_111 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_110 = _RAND_111[21:0];
  _RAND_112 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_111 = _RAND_112[21:0];
  _RAND_113 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_112 = _RAND_113[21:0];
  _RAND_114 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_113 = _RAND_114[21:0];
  _RAND_115 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_114 = _RAND_115[21:0];
  _RAND_116 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_115 = _RAND_116[21:0];
  _RAND_117 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_116 = _RAND_117[21:0];
  _RAND_118 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_117 = _RAND_118[21:0];
  _RAND_119 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_118 = _RAND_119[21:0];
  _RAND_120 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_119 = _RAND_120[21:0];
  _RAND_121 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_120 = _RAND_121[21:0];
  _RAND_122 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_121 = _RAND_122[21:0];
  _RAND_123 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_122 = _RAND_123[21:0];
  _RAND_124 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_123 = _RAND_124[21:0];
  _RAND_125 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_124 = _RAND_125[21:0];
  _RAND_126 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_125 = _RAND_126[21:0];
  _RAND_127 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_126 = _RAND_127[21:0];
  _RAND_128 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_127 = _RAND_128[21:0];
  _RAND_129 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_128 = _RAND_129[21:0];
  _RAND_130 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_129 = _RAND_130[21:0];
  _RAND_131 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_130 = _RAND_131[21:0];
  _RAND_132 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_131 = _RAND_132[21:0];
  _RAND_133 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_132 = _RAND_133[21:0];
  _RAND_134 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_133 = _RAND_134[21:0];
  _RAND_135 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_134 = _RAND_135[21:0];
  _RAND_136 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_135 = _RAND_136[21:0];
  _RAND_137 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_136 = _RAND_137[21:0];
  _RAND_138 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_137 = _RAND_138[21:0];
  _RAND_139 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_138 = _RAND_139[21:0];
  _RAND_140 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_139 = _RAND_140[21:0];
  _RAND_141 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_140 = _RAND_141[21:0];
  _RAND_142 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_141 = _RAND_142[21:0];
  _RAND_143 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_142 = _RAND_143[21:0];
  _RAND_144 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_143 = _RAND_144[21:0];
  _RAND_145 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_144 = _RAND_145[21:0];
  _RAND_146 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_145 = _RAND_146[21:0];
  _RAND_147 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_146 = _RAND_147[21:0];
  _RAND_148 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_147 = _RAND_148[21:0];
  _RAND_149 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_148 = _RAND_149[21:0];
  _RAND_150 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_149 = _RAND_150[21:0];
  _RAND_151 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_150 = _RAND_151[21:0];
  _RAND_152 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_151 = _RAND_152[21:0];
  _RAND_153 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_152 = _RAND_153[21:0];
  _RAND_154 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_153 = _RAND_154[21:0];
  _RAND_155 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_154 = _RAND_155[21:0];
  _RAND_156 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_155 = _RAND_156[21:0];
  _RAND_157 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_156 = _RAND_157[21:0];
  _RAND_158 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_157 = _RAND_158[21:0];
  _RAND_159 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_158 = _RAND_159[21:0];
  _RAND_160 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_159 = _RAND_160[21:0];
  _RAND_161 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_160 = _RAND_161[21:0];
  _RAND_162 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_161 = _RAND_162[21:0];
  _RAND_163 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_162 = _RAND_163[21:0];
  _RAND_164 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_163 = _RAND_164[21:0];
  _RAND_165 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_164 = _RAND_165[21:0];
  _RAND_166 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_165 = _RAND_166[21:0];
  _RAND_167 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_166 = _RAND_167[21:0];
  _RAND_168 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_167 = _RAND_168[21:0];
  _RAND_169 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_168 = _RAND_169[21:0];
  _RAND_170 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_169 = _RAND_170[21:0];
  _RAND_171 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_170 = _RAND_171[21:0];
  _RAND_172 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_171 = _RAND_172[21:0];
  _RAND_173 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_172 = _RAND_173[21:0];
  _RAND_174 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_173 = _RAND_174[21:0];
  _RAND_175 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_174 = _RAND_175[21:0];
  _RAND_176 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_175 = _RAND_176[21:0];
  _RAND_177 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_176 = _RAND_177[21:0];
  _RAND_178 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_177 = _RAND_178[21:0];
  _RAND_179 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_178 = _RAND_179[21:0];
  _RAND_180 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_179 = _RAND_180[21:0];
  _RAND_181 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_180 = _RAND_181[21:0];
  _RAND_182 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_181 = _RAND_182[21:0];
  _RAND_183 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_182 = _RAND_183[21:0];
  _RAND_184 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_183 = _RAND_184[21:0];
  _RAND_185 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_184 = _RAND_185[21:0];
  _RAND_186 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_185 = _RAND_186[21:0];
  _RAND_187 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_186 = _RAND_187[21:0];
  _RAND_188 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_187 = _RAND_188[21:0];
  _RAND_189 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_188 = _RAND_189[21:0];
  _RAND_190 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_189 = _RAND_190[21:0];
  _RAND_191 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_190 = _RAND_191[21:0];
  _RAND_192 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_191 = _RAND_192[21:0];
  _RAND_193 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_192 = _RAND_193[21:0];
  _RAND_194 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_193 = _RAND_194[21:0];
  _RAND_195 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_194 = _RAND_195[21:0];
  _RAND_196 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_195 = _RAND_196[21:0];
  _RAND_197 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_196 = _RAND_197[21:0];
  _RAND_198 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_197 = _RAND_198[21:0];
  _RAND_199 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_198 = _RAND_199[21:0];
  _RAND_200 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_199 = _RAND_200[21:0];
  _RAND_201 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_200 = _RAND_201[21:0];
  _RAND_202 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_201 = _RAND_202[21:0];
  _RAND_203 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_202 = _RAND_203[21:0];
  _RAND_204 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_203 = _RAND_204[21:0];
  _RAND_205 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_204 = _RAND_205[21:0];
  _RAND_206 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_205 = _RAND_206[21:0];
  _RAND_207 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_206 = _RAND_207[21:0];
  _RAND_208 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_207 = _RAND_208[21:0];
  _RAND_209 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_208 = _RAND_209[21:0];
  _RAND_210 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_209 = _RAND_210[21:0];
  _RAND_211 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_210 = _RAND_211[21:0];
  _RAND_212 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_211 = _RAND_212[21:0];
  _RAND_213 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_212 = _RAND_213[21:0];
  _RAND_214 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_213 = _RAND_214[21:0];
  _RAND_215 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_214 = _RAND_215[21:0];
  _RAND_216 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_215 = _RAND_216[21:0];
  _RAND_217 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_216 = _RAND_217[21:0];
  _RAND_218 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_217 = _RAND_218[21:0];
  _RAND_219 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_218 = _RAND_219[21:0];
  _RAND_220 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_219 = _RAND_220[21:0];
  _RAND_221 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_220 = _RAND_221[21:0];
  _RAND_222 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_221 = _RAND_222[21:0];
  _RAND_223 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_222 = _RAND_223[21:0];
  _RAND_224 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_223 = _RAND_224[21:0];
  _RAND_225 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_224 = _RAND_225[21:0];
  _RAND_226 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_225 = _RAND_226[21:0];
  _RAND_227 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_226 = _RAND_227[21:0];
  _RAND_228 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_227 = _RAND_228[21:0];
  _RAND_229 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_228 = _RAND_229[21:0];
  _RAND_230 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_229 = _RAND_230[21:0];
  _RAND_231 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_230 = _RAND_231[21:0];
  _RAND_232 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_231 = _RAND_232[21:0];
  _RAND_233 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_232 = _RAND_233[21:0];
  _RAND_234 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_233 = _RAND_234[21:0];
  _RAND_235 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_234 = _RAND_235[21:0];
  _RAND_236 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_235 = _RAND_236[21:0];
  _RAND_237 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_236 = _RAND_237[21:0];
  _RAND_238 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_237 = _RAND_238[21:0];
  _RAND_239 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_238 = _RAND_239[21:0];
  _RAND_240 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_239 = _RAND_240[21:0];
  _RAND_241 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_240 = _RAND_241[21:0];
  _RAND_242 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_241 = _RAND_242[21:0];
  _RAND_243 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_242 = _RAND_243[21:0];
  _RAND_244 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_243 = _RAND_244[21:0];
  _RAND_245 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_244 = _RAND_245[21:0];
  _RAND_246 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_245 = _RAND_246[21:0];
  _RAND_247 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_246 = _RAND_247[21:0];
  _RAND_248 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_247 = _RAND_248[21:0];
  _RAND_249 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_248 = _RAND_249[21:0];
  _RAND_250 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_249 = _RAND_250[21:0];
  _RAND_251 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_250 = _RAND_251[21:0];
  _RAND_252 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_251 = _RAND_252[21:0];
  _RAND_253 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_252 = _RAND_253[21:0];
  _RAND_254 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_253 = _RAND_254[21:0];
  _RAND_255 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_254 = _RAND_255[21:0];
  _RAND_256 = {1{`RANDOM}};
  btb_bank0_rd_data_way0_out_255 = _RAND_256[21:0];
  _RAND_257 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_0 = _RAND_257[21:0];
  _RAND_258 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_1 = _RAND_258[21:0];
  _RAND_259 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_2 = _RAND_259[21:0];
  _RAND_260 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_3 = _RAND_260[21:0];
  _RAND_261 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_4 = _RAND_261[21:0];
  _RAND_262 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_5 = _RAND_262[21:0];
  _RAND_263 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_6 = _RAND_263[21:0];
  _RAND_264 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_7 = _RAND_264[21:0];
  _RAND_265 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_8 = _RAND_265[21:0];
  _RAND_266 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_9 = _RAND_266[21:0];
  _RAND_267 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_10 = _RAND_267[21:0];
  _RAND_268 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_11 = _RAND_268[21:0];
  _RAND_269 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_12 = _RAND_269[21:0];
  _RAND_270 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_13 = _RAND_270[21:0];
  _RAND_271 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_14 = _RAND_271[21:0];
  _RAND_272 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_15 = _RAND_272[21:0];
  _RAND_273 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_16 = _RAND_273[21:0];
  _RAND_274 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_17 = _RAND_274[21:0];
  _RAND_275 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_18 = _RAND_275[21:0];
  _RAND_276 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_19 = _RAND_276[21:0];
  _RAND_277 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_20 = _RAND_277[21:0];
  _RAND_278 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_21 = _RAND_278[21:0];
  _RAND_279 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_22 = _RAND_279[21:0];
  _RAND_280 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_23 = _RAND_280[21:0];
  _RAND_281 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_24 = _RAND_281[21:0];
  _RAND_282 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_25 = _RAND_282[21:0];
  _RAND_283 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_26 = _RAND_283[21:0];
  _RAND_284 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_27 = _RAND_284[21:0];
  _RAND_285 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_28 = _RAND_285[21:0];
  _RAND_286 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_29 = _RAND_286[21:0];
  _RAND_287 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_30 = _RAND_287[21:0];
  _RAND_288 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_31 = _RAND_288[21:0];
  _RAND_289 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_32 = _RAND_289[21:0];
  _RAND_290 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_33 = _RAND_290[21:0];
  _RAND_291 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_34 = _RAND_291[21:0];
  _RAND_292 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_35 = _RAND_292[21:0];
  _RAND_293 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_36 = _RAND_293[21:0];
  _RAND_294 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_37 = _RAND_294[21:0];
  _RAND_295 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_38 = _RAND_295[21:0];
  _RAND_296 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_39 = _RAND_296[21:0];
  _RAND_297 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_40 = _RAND_297[21:0];
  _RAND_298 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_41 = _RAND_298[21:0];
  _RAND_299 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_42 = _RAND_299[21:0];
  _RAND_300 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_43 = _RAND_300[21:0];
  _RAND_301 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_44 = _RAND_301[21:0];
  _RAND_302 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_45 = _RAND_302[21:0];
  _RAND_303 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_46 = _RAND_303[21:0];
  _RAND_304 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_47 = _RAND_304[21:0];
  _RAND_305 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_48 = _RAND_305[21:0];
  _RAND_306 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_49 = _RAND_306[21:0];
  _RAND_307 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_50 = _RAND_307[21:0];
  _RAND_308 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_51 = _RAND_308[21:0];
  _RAND_309 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_52 = _RAND_309[21:0];
  _RAND_310 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_53 = _RAND_310[21:0];
  _RAND_311 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_54 = _RAND_311[21:0];
  _RAND_312 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_55 = _RAND_312[21:0];
  _RAND_313 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_56 = _RAND_313[21:0];
  _RAND_314 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_57 = _RAND_314[21:0];
  _RAND_315 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_58 = _RAND_315[21:0];
  _RAND_316 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_59 = _RAND_316[21:0];
  _RAND_317 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_60 = _RAND_317[21:0];
  _RAND_318 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_61 = _RAND_318[21:0];
  _RAND_319 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_62 = _RAND_319[21:0];
  _RAND_320 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_63 = _RAND_320[21:0];
  _RAND_321 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_64 = _RAND_321[21:0];
  _RAND_322 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_65 = _RAND_322[21:0];
  _RAND_323 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_66 = _RAND_323[21:0];
  _RAND_324 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_67 = _RAND_324[21:0];
  _RAND_325 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_68 = _RAND_325[21:0];
  _RAND_326 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_69 = _RAND_326[21:0];
  _RAND_327 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_70 = _RAND_327[21:0];
  _RAND_328 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_71 = _RAND_328[21:0];
  _RAND_329 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_72 = _RAND_329[21:0];
  _RAND_330 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_73 = _RAND_330[21:0];
  _RAND_331 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_74 = _RAND_331[21:0];
  _RAND_332 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_75 = _RAND_332[21:0];
  _RAND_333 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_76 = _RAND_333[21:0];
  _RAND_334 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_77 = _RAND_334[21:0];
  _RAND_335 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_78 = _RAND_335[21:0];
  _RAND_336 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_79 = _RAND_336[21:0];
  _RAND_337 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_80 = _RAND_337[21:0];
  _RAND_338 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_81 = _RAND_338[21:0];
  _RAND_339 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_82 = _RAND_339[21:0];
  _RAND_340 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_83 = _RAND_340[21:0];
  _RAND_341 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_84 = _RAND_341[21:0];
  _RAND_342 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_85 = _RAND_342[21:0];
  _RAND_343 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_86 = _RAND_343[21:0];
  _RAND_344 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_87 = _RAND_344[21:0];
  _RAND_345 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_88 = _RAND_345[21:0];
  _RAND_346 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_89 = _RAND_346[21:0];
  _RAND_347 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_90 = _RAND_347[21:0];
  _RAND_348 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_91 = _RAND_348[21:0];
  _RAND_349 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_92 = _RAND_349[21:0];
  _RAND_350 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_93 = _RAND_350[21:0];
  _RAND_351 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_94 = _RAND_351[21:0];
  _RAND_352 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_95 = _RAND_352[21:0];
  _RAND_353 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_96 = _RAND_353[21:0];
  _RAND_354 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_97 = _RAND_354[21:0];
  _RAND_355 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_98 = _RAND_355[21:0];
  _RAND_356 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_99 = _RAND_356[21:0];
  _RAND_357 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_100 = _RAND_357[21:0];
  _RAND_358 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_101 = _RAND_358[21:0];
  _RAND_359 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_102 = _RAND_359[21:0];
  _RAND_360 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_103 = _RAND_360[21:0];
  _RAND_361 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_104 = _RAND_361[21:0];
  _RAND_362 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_105 = _RAND_362[21:0];
  _RAND_363 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_106 = _RAND_363[21:0];
  _RAND_364 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_107 = _RAND_364[21:0];
  _RAND_365 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_108 = _RAND_365[21:0];
  _RAND_366 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_109 = _RAND_366[21:0];
  _RAND_367 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_110 = _RAND_367[21:0];
  _RAND_368 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_111 = _RAND_368[21:0];
  _RAND_369 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_112 = _RAND_369[21:0];
  _RAND_370 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_113 = _RAND_370[21:0];
  _RAND_371 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_114 = _RAND_371[21:0];
  _RAND_372 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_115 = _RAND_372[21:0];
  _RAND_373 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_116 = _RAND_373[21:0];
  _RAND_374 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_117 = _RAND_374[21:0];
  _RAND_375 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_118 = _RAND_375[21:0];
  _RAND_376 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_119 = _RAND_376[21:0];
  _RAND_377 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_120 = _RAND_377[21:0];
  _RAND_378 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_121 = _RAND_378[21:0];
  _RAND_379 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_122 = _RAND_379[21:0];
  _RAND_380 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_123 = _RAND_380[21:0];
  _RAND_381 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_124 = _RAND_381[21:0];
  _RAND_382 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_125 = _RAND_382[21:0];
  _RAND_383 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_126 = _RAND_383[21:0];
  _RAND_384 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_127 = _RAND_384[21:0];
  _RAND_385 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_128 = _RAND_385[21:0];
  _RAND_386 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_129 = _RAND_386[21:0];
  _RAND_387 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_130 = _RAND_387[21:0];
  _RAND_388 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_131 = _RAND_388[21:0];
  _RAND_389 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_132 = _RAND_389[21:0];
  _RAND_390 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_133 = _RAND_390[21:0];
  _RAND_391 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_134 = _RAND_391[21:0];
  _RAND_392 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_135 = _RAND_392[21:0];
  _RAND_393 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_136 = _RAND_393[21:0];
  _RAND_394 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_137 = _RAND_394[21:0];
  _RAND_395 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_138 = _RAND_395[21:0];
  _RAND_396 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_139 = _RAND_396[21:0];
  _RAND_397 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_140 = _RAND_397[21:0];
  _RAND_398 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_141 = _RAND_398[21:0];
  _RAND_399 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_142 = _RAND_399[21:0];
  _RAND_400 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_143 = _RAND_400[21:0];
  _RAND_401 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_144 = _RAND_401[21:0];
  _RAND_402 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_145 = _RAND_402[21:0];
  _RAND_403 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_146 = _RAND_403[21:0];
  _RAND_404 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_147 = _RAND_404[21:0];
  _RAND_405 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_148 = _RAND_405[21:0];
  _RAND_406 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_149 = _RAND_406[21:0];
  _RAND_407 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_150 = _RAND_407[21:0];
  _RAND_408 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_151 = _RAND_408[21:0];
  _RAND_409 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_152 = _RAND_409[21:0];
  _RAND_410 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_153 = _RAND_410[21:0];
  _RAND_411 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_154 = _RAND_411[21:0];
  _RAND_412 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_155 = _RAND_412[21:0];
  _RAND_413 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_156 = _RAND_413[21:0];
  _RAND_414 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_157 = _RAND_414[21:0];
  _RAND_415 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_158 = _RAND_415[21:0];
  _RAND_416 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_159 = _RAND_416[21:0];
  _RAND_417 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_160 = _RAND_417[21:0];
  _RAND_418 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_161 = _RAND_418[21:0];
  _RAND_419 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_162 = _RAND_419[21:0];
  _RAND_420 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_163 = _RAND_420[21:0];
  _RAND_421 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_164 = _RAND_421[21:0];
  _RAND_422 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_165 = _RAND_422[21:0];
  _RAND_423 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_166 = _RAND_423[21:0];
  _RAND_424 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_167 = _RAND_424[21:0];
  _RAND_425 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_168 = _RAND_425[21:0];
  _RAND_426 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_169 = _RAND_426[21:0];
  _RAND_427 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_170 = _RAND_427[21:0];
  _RAND_428 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_171 = _RAND_428[21:0];
  _RAND_429 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_172 = _RAND_429[21:0];
  _RAND_430 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_173 = _RAND_430[21:0];
  _RAND_431 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_174 = _RAND_431[21:0];
  _RAND_432 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_175 = _RAND_432[21:0];
  _RAND_433 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_176 = _RAND_433[21:0];
  _RAND_434 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_177 = _RAND_434[21:0];
  _RAND_435 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_178 = _RAND_435[21:0];
  _RAND_436 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_179 = _RAND_436[21:0];
  _RAND_437 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_180 = _RAND_437[21:0];
  _RAND_438 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_181 = _RAND_438[21:0];
  _RAND_439 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_182 = _RAND_439[21:0];
  _RAND_440 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_183 = _RAND_440[21:0];
  _RAND_441 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_184 = _RAND_441[21:0];
  _RAND_442 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_185 = _RAND_442[21:0];
  _RAND_443 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_186 = _RAND_443[21:0];
  _RAND_444 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_187 = _RAND_444[21:0];
  _RAND_445 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_188 = _RAND_445[21:0];
  _RAND_446 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_189 = _RAND_446[21:0];
  _RAND_447 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_190 = _RAND_447[21:0];
  _RAND_448 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_191 = _RAND_448[21:0];
  _RAND_449 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_192 = _RAND_449[21:0];
  _RAND_450 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_193 = _RAND_450[21:0];
  _RAND_451 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_194 = _RAND_451[21:0];
  _RAND_452 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_195 = _RAND_452[21:0];
  _RAND_453 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_196 = _RAND_453[21:0];
  _RAND_454 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_197 = _RAND_454[21:0];
  _RAND_455 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_198 = _RAND_455[21:0];
  _RAND_456 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_199 = _RAND_456[21:0];
  _RAND_457 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_200 = _RAND_457[21:0];
  _RAND_458 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_201 = _RAND_458[21:0];
  _RAND_459 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_202 = _RAND_459[21:0];
  _RAND_460 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_203 = _RAND_460[21:0];
  _RAND_461 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_204 = _RAND_461[21:0];
  _RAND_462 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_205 = _RAND_462[21:0];
  _RAND_463 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_206 = _RAND_463[21:0];
  _RAND_464 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_207 = _RAND_464[21:0];
  _RAND_465 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_208 = _RAND_465[21:0];
  _RAND_466 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_209 = _RAND_466[21:0];
  _RAND_467 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_210 = _RAND_467[21:0];
  _RAND_468 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_211 = _RAND_468[21:0];
  _RAND_469 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_212 = _RAND_469[21:0];
  _RAND_470 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_213 = _RAND_470[21:0];
  _RAND_471 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_214 = _RAND_471[21:0];
  _RAND_472 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_215 = _RAND_472[21:0];
  _RAND_473 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_216 = _RAND_473[21:0];
  _RAND_474 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_217 = _RAND_474[21:0];
  _RAND_475 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_218 = _RAND_475[21:0];
  _RAND_476 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_219 = _RAND_476[21:0];
  _RAND_477 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_220 = _RAND_477[21:0];
  _RAND_478 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_221 = _RAND_478[21:0];
  _RAND_479 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_222 = _RAND_479[21:0];
  _RAND_480 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_223 = _RAND_480[21:0];
  _RAND_481 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_224 = _RAND_481[21:0];
  _RAND_482 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_225 = _RAND_482[21:0];
  _RAND_483 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_226 = _RAND_483[21:0];
  _RAND_484 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_227 = _RAND_484[21:0];
  _RAND_485 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_228 = _RAND_485[21:0];
  _RAND_486 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_229 = _RAND_486[21:0];
  _RAND_487 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_230 = _RAND_487[21:0];
  _RAND_488 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_231 = _RAND_488[21:0];
  _RAND_489 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_232 = _RAND_489[21:0];
  _RAND_490 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_233 = _RAND_490[21:0];
  _RAND_491 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_234 = _RAND_491[21:0];
  _RAND_492 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_235 = _RAND_492[21:0];
  _RAND_493 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_236 = _RAND_493[21:0];
  _RAND_494 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_237 = _RAND_494[21:0];
  _RAND_495 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_238 = _RAND_495[21:0];
  _RAND_496 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_239 = _RAND_496[21:0];
  _RAND_497 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_240 = _RAND_497[21:0];
  _RAND_498 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_241 = _RAND_498[21:0];
  _RAND_499 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_242 = _RAND_499[21:0];
  _RAND_500 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_243 = _RAND_500[21:0];
  _RAND_501 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_244 = _RAND_501[21:0];
  _RAND_502 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_245 = _RAND_502[21:0];
  _RAND_503 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_246 = _RAND_503[21:0];
  _RAND_504 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_247 = _RAND_504[21:0];
  _RAND_505 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_248 = _RAND_505[21:0];
  _RAND_506 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_249 = _RAND_506[21:0];
  _RAND_507 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_250 = _RAND_507[21:0];
  _RAND_508 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_251 = _RAND_508[21:0];
  _RAND_509 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_252 = _RAND_509[21:0];
  _RAND_510 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_253 = _RAND_510[21:0];
  _RAND_511 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_254 = _RAND_511[21:0];
  _RAND_512 = {1{`RANDOM}};
  btb_bank0_rd_data_way1_out_255 = _RAND_512[21:0];
  _RAND_513 = {1{`RANDOM}};
  fghr = _RAND_513[7:0];
  _RAND_514 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_0 = _RAND_514[1:0];
  _RAND_515 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_1 = _RAND_515[1:0];
  _RAND_516 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_2 = _RAND_516[1:0];
  _RAND_517 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_3 = _RAND_517[1:0];
  _RAND_518 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_4 = _RAND_518[1:0];
  _RAND_519 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_5 = _RAND_519[1:0];
  _RAND_520 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_6 = _RAND_520[1:0];
  _RAND_521 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_7 = _RAND_521[1:0];
  _RAND_522 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_8 = _RAND_522[1:0];
  _RAND_523 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_9 = _RAND_523[1:0];
  _RAND_524 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_10 = _RAND_524[1:0];
  _RAND_525 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_11 = _RAND_525[1:0];
  _RAND_526 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_12 = _RAND_526[1:0];
  _RAND_527 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_13 = _RAND_527[1:0];
  _RAND_528 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_14 = _RAND_528[1:0];
  _RAND_529 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_15 = _RAND_529[1:0];
  _RAND_530 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_16 = _RAND_530[1:0];
  _RAND_531 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_17 = _RAND_531[1:0];
  _RAND_532 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_18 = _RAND_532[1:0];
  _RAND_533 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_19 = _RAND_533[1:0];
  _RAND_534 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_20 = _RAND_534[1:0];
  _RAND_535 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_21 = _RAND_535[1:0];
  _RAND_536 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_22 = _RAND_536[1:0];
  _RAND_537 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_23 = _RAND_537[1:0];
  _RAND_538 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_24 = _RAND_538[1:0];
  _RAND_539 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_25 = _RAND_539[1:0];
  _RAND_540 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_26 = _RAND_540[1:0];
  _RAND_541 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_27 = _RAND_541[1:0];
  _RAND_542 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_28 = _RAND_542[1:0];
  _RAND_543 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_29 = _RAND_543[1:0];
  _RAND_544 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_30 = _RAND_544[1:0];
  _RAND_545 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_31 = _RAND_545[1:0];
  _RAND_546 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_32 = _RAND_546[1:0];
  _RAND_547 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_33 = _RAND_547[1:0];
  _RAND_548 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_34 = _RAND_548[1:0];
  _RAND_549 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_35 = _RAND_549[1:0];
  _RAND_550 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_36 = _RAND_550[1:0];
  _RAND_551 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_37 = _RAND_551[1:0];
  _RAND_552 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_38 = _RAND_552[1:0];
  _RAND_553 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_39 = _RAND_553[1:0];
  _RAND_554 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_40 = _RAND_554[1:0];
  _RAND_555 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_41 = _RAND_555[1:0];
  _RAND_556 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_42 = _RAND_556[1:0];
  _RAND_557 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_43 = _RAND_557[1:0];
  _RAND_558 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_44 = _RAND_558[1:0];
  _RAND_559 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_45 = _RAND_559[1:0];
  _RAND_560 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_46 = _RAND_560[1:0];
  _RAND_561 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_47 = _RAND_561[1:0];
  _RAND_562 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_48 = _RAND_562[1:0];
  _RAND_563 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_49 = _RAND_563[1:0];
  _RAND_564 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_50 = _RAND_564[1:0];
  _RAND_565 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_51 = _RAND_565[1:0];
  _RAND_566 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_52 = _RAND_566[1:0];
  _RAND_567 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_53 = _RAND_567[1:0];
  _RAND_568 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_54 = _RAND_568[1:0];
  _RAND_569 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_55 = _RAND_569[1:0];
  _RAND_570 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_56 = _RAND_570[1:0];
  _RAND_571 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_57 = _RAND_571[1:0];
  _RAND_572 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_58 = _RAND_572[1:0];
  _RAND_573 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_59 = _RAND_573[1:0];
  _RAND_574 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_60 = _RAND_574[1:0];
  _RAND_575 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_61 = _RAND_575[1:0];
  _RAND_576 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_62 = _RAND_576[1:0];
  _RAND_577 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_63 = _RAND_577[1:0];
  _RAND_578 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_64 = _RAND_578[1:0];
  _RAND_579 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_65 = _RAND_579[1:0];
  _RAND_580 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_66 = _RAND_580[1:0];
  _RAND_581 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_67 = _RAND_581[1:0];
  _RAND_582 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_68 = _RAND_582[1:0];
  _RAND_583 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_69 = _RAND_583[1:0];
  _RAND_584 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_70 = _RAND_584[1:0];
  _RAND_585 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_71 = _RAND_585[1:0];
  _RAND_586 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_72 = _RAND_586[1:0];
  _RAND_587 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_73 = _RAND_587[1:0];
  _RAND_588 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_74 = _RAND_588[1:0];
  _RAND_589 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_75 = _RAND_589[1:0];
  _RAND_590 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_76 = _RAND_590[1:0];
  _RAND_591 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_77 = _RAND_591[1:0];
  _RAND_592 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_78 = _RAND_592[1:0];
  _RAND_593 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_79 = _RAND_593[1:0];
  _RAND_594 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_80 = _RAND_594[1:0];
  _RAND_595 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_81 = _RAND_595[1:0];
  _RAND_596 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_82 = _RAND_596[1:0];
  _RAND_597 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_83 = _RAND_597[1:0];
  _RAND_598 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_84 = _RAND_598[1:0];
  _RAND_599 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_85 = _RAND_599[1:0];
  _RAND_600 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_86 = _RAND_600[1:0];
  _RAND_601 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_87 = _RAND_601[1:0];
  _RAND_602 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_88 = _RAND_602[1:0];
  _RAND_603 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_89 = _RAND_603[1:0];
  _RAND_604 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_90 = _RAND_604[1:0];
  _RAND_605 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_91 = _RAND_605[1:0];
  _RAND_606 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_92 = _RAND_606[1:0];
  _RAND_607 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_93 = _RAND_607[1:0];
  _RAND_608 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_94 = _RAND_608[1:0];
  _RAND_609 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_95 = _RAND_609[1:0];
  _RAND_610 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_96 = _RAND_610[1:0];
  _RAND_611 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_97 = _RAND_611[1:0];
  _RAND_612 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_98 = _RAND_612[1:0];
  _RAND_613 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_99 = _RAND_613[1:0];
  _RAND_614 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_100 = _RAND_614[1:0];
  _RAND_615 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_101 = _RAND_615[1:0];
  _RAND_616 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_102 = _RAND_616[1:0];
  _RAND_617 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_103 = _RAND_617[1:0];
  _RAND_618 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_104 = _RAND_618[1:0];
  _RAND_619 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_105 = _RAND_619[1:0];
  _RAND_620 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_106 = _RAND_620[1:0];
  _RAND_621 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_107 = _RAND_621[1:0];
  _RAND_622 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_108 = _RAND_622[1:0];
  _RAND_623 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_109 = _RAND_623[1:0];
  _RAND_624 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_110 = _RAND_624[1:0];
  _RAND_625 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_111 = _RAND_625[1:0];
  _RAND_626 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_112 = _RAND_626[1:0];
  _RAND_627 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_113 = _RAND_627[1:0];
  _RAND_628 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_114 = _RAND_628[1:0];
  _RAND_629 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_115 = _RAND_629[1:0];
  _RAND_630 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_116 = _RAND_630[1:0];
  _RAND_631 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_117 = _RAND_631[1:0];
  _RAND_632 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_118 = _RAND_632[1:0];
  _RAND_633 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_119 = _RAND_633[1:0];
  _RAND_634 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_120 = _RAND_634[1:0];
  _RAND_635 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_121 = _RAND_635[1:0];
  _RAND_636 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_122 = _RAND_636[1:0];
  _RAND_637 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_123 = _RAND_637[1:0];
  _RAND_638 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_124 = _RAND_638[1:0];
  _RAND_639 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_125 = _RAND_639[1:0];
  _RAND_640 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_126 = _RAND_640[1:0];
  _RAND_641 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_127 = _RAND_641[1:0];
  _RAND_642 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_128 = _RAND_642[1:0];
  _RAND_643 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_129 = _RAND_643[1:0];
  _RAND_644 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_130 = _RAND_644[1:0];
  _RAND_645 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_131 = _RAND_645[1:0];
  _RAND_646 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_132 = _RAND_646[1:0];
  _RAND_647 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_133 = _RAND_647[1:0];
  _RAND_648 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_134 = _RAND_648[1:0];
  _RAND_649 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_135 = _RAND_649[1:0];
  _RAND_650 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_136 = _RAND_650[1:0];
  _RAND_651 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_137 = _RAND_651[1:0];
  _RAND_652 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_138 = _RAND_652[1:0];
  _RAND_653 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_139 = _RAND_653[1:0];
  _RAND_654 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_140 = _RAND_654[1:0];
  _RAND_655 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_141 = _RAND_655[1:0];
  _RAND_656 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_142 = _RAND_656[1:0];
  _RAND_657 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_143 = _RAND_657[1:0];
  _RAND_658 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_144 = _RAND_658[1:0];
  _RAND_659 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_145 = _RAND_659[1:0];
  _RAND_660 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_146 = _RAND_660[1:0];
  _RAND_661 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_147 = _RAND_661[1:0];
  _RAND_662 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_148 = _RAND_662[1:0];
  _RAND_663 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_149 = _RAND_663[1:0];
  _RAND_664 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_150 = _RAND_664[1:0];
  _RAND_665 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_151 = _RAND_665[1:0];
  _RAND_666 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_152 = _RAND_666[1:0];
  _RAND_667 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_153 = _RAND_667[1:0];
  _RAND_668 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_154 = _RAND_668[1:0];
  _RAND_669 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_155 = _RAND_669[1:0];
  _RAND_670 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_156 = _RAND_670[1:0];
  _RAND_671 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_157 = _RAND_671[1:0];
  _RAND_672 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_158 = _RAND_672[1:0];
  _RAND_673 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_159 = _RAND_673[1:0];
  _RAND_674 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_160 = _RAND_674[1:0];
  _RAND_675 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_161 = _RAND_675[1:0];
  _RAND_676 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_162 = _RAND_676[1:0];
  _RAND_677 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_163 = _RAND_677[1:0];
  _RAND_678 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_164 = _RAND_678[1:0];
  _RAND_679 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_165 = _RAND_679[1:0];
  _RAND_680 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_166 = _RAND_680[1:0];
  _RAND_681 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_167 = _RAND_681[1:0];
  _RAND_682 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_168 = _RAND_682[1:0];
  _RAND_683 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_169 = _RAND_683[1:0];
  _RAND_684 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_170 = _RAND_684[1:0];
  _RAND_685 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_171 = _RAND_685[1:0];
  _RAND_686 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_172 = _RAND_686[1:0];
  _RAND_687 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_173 = _RAND_687[1:0];
  _RAND_688 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_174 = _RAND_688[1:0];
  _RAND_689 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_175 = _RAND_689[1:0];
  _RAND_690 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_176 = _RAND_690[1:0];
  _RAND_691 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_177 = _RAND_691[1:0];
  _RAND_692 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_178 = _RAND_692[1:0];
  _RAND_693 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_179 = _RAND_693[1:0];
  _RAND_694 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_180 = _RAND_694[1:0];
  _RAND_695 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_181 = _RAND_695[1:0];
  _RAND_696 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_182 = _RAND_696[1:0];
  _RAND_697 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_183 = _RAND_697[1:0];
  _RAND_698 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_184 = _RAND_698[1:0];
  _RAND_699 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_185 = _RAND_699[1:0];
  _RAND_700 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_186 = _RAND_700[1:0];
  _RAND_701 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_187 = _RAND_701[1:0];
  _RAND_702 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_188 = _RAND_702[1:0];
  _RAND_703 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_189 = _RAND_703[1:0];
  _RAND_704 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_190 = _RAND_704[1:0];
  _RAND_705 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_191 = _RAND_705[1:0];
  _RAND_706 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_192 = _RAND_706[1:0];
  _RAND_707 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_193 = _RAND_707[1:0];
  _RAND_708 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_194 = _RAND_708[1:0];
  _RAND_709 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_195 = _RAND_709[1:0];
  _RAND_710 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_196 = _RAND_710[1:0];
  _RAND_711 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_197 = _RAND_711[1:0];
  _RAND_712 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_198 = _RAND_712[1:0];
  _RAND_713 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_199 = _RAND_713[1:0];
  _RAND_714 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_200 = _RAND_714[1:0];
  _RAND_715 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_201 = _RAND_715[1:0];
  _RAND_716 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_202 = _RAND_716[1:0];
  _RAND_717 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_203 = _RAND_717[1:0];
  _RAND_718 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_204 = _RAND_718[1:0];
  _RAND_719 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_205 = _RAND_719[1:0];
  _RAND_720 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_206 = _RAND_720[1:0];
  _RAND_721 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_207 = _RAND_721[1:0];
  _RAND_722 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_208 = _RAND_722[1:0];
  _RAND_723 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_209 = _RAND_723[1:0];
  _RAND_724 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_210 = _RAND_724[1:0];
  _RAND_725 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_211 = _RAND_725[1:0];
  _RAND_726 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_212 = _RAND_726[1:0];
  _RAND_727 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_213 = _RAND_727[1:0];
  _RAND_728 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_214 = _RAND_728[1:0];
  _RAND_729 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_215 = _RAND_729[1:0];
  _RAND_730 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_216 = _RAND_730[1:0];
  _RAND_731 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_217 = _RAND_731[1:0];
  _RAND_732 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_218 = _RAND_732[1:0];
  _RAND_733 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_219 = _RAND_733[1:0];
  _RAND_734 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_220 = _RAND_734[1:0];
  _RAND_735 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_221 = _RAND_735[1:0];
  _RAND_736 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_222 = _RAND_736[1:0];
  _RAND_737 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_223 = _RAND_737[1:0];
  _RAND_738 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_224 = _RAND_738[1:0];
  _RAND_739 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_225 = _RAND_739[1:0];
  _RAND_740 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_226 = _RAND_740[1:0];
  _RAND_741 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_227 = _RAND_741[1:0];
  _RAND_742 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_228 = _RAND_742[1:0];
  _RAND_743 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_229 = _RAND_743[1:0];
  _RAND_744 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_230 = _RAND_744[1:0];
  _RAND_745 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_231 = _RAND_745[1:0];
  _RAND_746 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_232 = _RAND_746[1:0];
  _RAND_747 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_233 = _RAND_747[1:0];
  _RAND_748 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_234 = _RAND_748[1:0];
  _RAND_749 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_235 = _RAND_749[1:0];
  _RAND_750 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_236 = _RAND_750[1:0];
  _RAND_751 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_237 = _RAND_751[1:0];
  _RAND_752 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_238 = _RAND_752[1:0];
  _RAND_753 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_239 = _RAND_753[1:0];
  _RAND_754 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_240 = _RAND_754[1:0];
  _RAND_755 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_241 = _RAND_755[1:0];
  _RAND_756 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_242 = _RAND_756[1:0];
  _RAND_757 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_243 = _RAND_757[1:0];
  _RAND_758 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_244 = _RAND_758[1:0];
  _RAND_759 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_245 = _RAND_759[1:0];
  _RAND_760 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_246 = _RAND_760[1:0];
  _RAND_761 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_247 = _RAND_761[1:0];
  _RAND_762 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_248 = _RAND_762[1:0];
  _RAND_763 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_249 = _RAND_763[1:0];
  _RAND_764 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_250 = _RAND_764[1:0];
  _RAND_765 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_251 = _RAND_765[1:0];
  _RAND_766 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_252 = _RAND_766[1:0];
  _RAND_767 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_253 = _RAND_767[1:0];
  _RAND_768 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_254 = _RAND_768[1:0];
  _RAND_769 = {1{`RANDOM}};
  bht_bank_rd_data_out_1_255 = _RAND_769[1:0];
  _RAND_770 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_0 = _RAND_770[1:0];
  _RAND_771 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_1 = _RAND_771[1:0];
  _RAND_772 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_2 = _RAND_772[1:0];
  _RAND_773 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_3 = _RAND_773[1:0];
  _RAND_774 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_4 = _RAND_774[1:0];
  _RAND_775 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_5 = _RAND_775[1:0];
  _RAND_776 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_6 = _RAND_776[1:0];
  _RAND_777 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_7 = _RAND_777[1:0];
  _RAND_778 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_8 = _RAND_778[1:0];
  _RAND_779 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_9 = _RAND_779[1:0];
  _RAND_780 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_10 = _RAND_780[1:0];
  _RAND_781 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_11 = _RAND_781[1:0];
  _RAND_782 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_12 = _RAND_782[1:0];
  _RAND_783 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_13 = _RAND_783[1:0];
  _RAND_784 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_14 = _RAND_784[1:0];
  _RAND_785 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_15 = _RAND_785[1:0];
  _RAND_786 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_16 = _RAND_786[1:0];
  _RAND_787 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_17 = _RAND_787[1:0];
  _RAND_788 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_18 = _RAND_788[1:0];
  _RAND_789 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_19 = _RAND_789[1:0];
  _RAND_790 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_20 = _RAND_790[1:0];
  _RAND_791 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_21 = _RAND_791[1:0];
  _RAND_792 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_22 = _RAND_792[1:0];
  _RAND_793 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_23 = _RAND_793[1:0];
  _RAND_794 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_24 = _RAND_794[1:0];
  _RAND_795 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_25 = _RAND_795[1:0];
  _RAND_796 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_26 = _RAND_796[1:0];
  _RAND_797 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_27 = _RAND_797[1:0];
  _RAND_798 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_28 = _RAND_798[1:0];
  _RAND_799 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_29 = _RAND_799[1:0];
  _RAND_800 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_30 = _RAND_800[1:0];
  _RAND_801 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_31 = _RAND_801[1:0];
  _RAND_802 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_32 = _RAND_802[1:0];
  _RAND_803 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_33 = _RAND_803[1:0];
  _RAND_804 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_34 = _RAND_804[1:0];
  _RAND_805 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_35 = _RAND_805[1:0];
  _RAND_806 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_36 = _RAND_806[1:0];
  _RAND_807 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_37 = _RAND_807[1:0];
  _RAND_808 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_38 = _RAND_808[1:0];
  _RAND_809 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_39 = _RAND_809[1:0];
  _RAND_810 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_40 = _RAND_810[1:0];
  _RAND_811 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_41 = _RAND_811[1:0];
  _RAND_812 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_42 = _RAND_812[1:0];
  _RAND_813 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_43 = _RAND_813[1:0];
  _RAND_814 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_44 = _RAND_814[1:0];
  _RAND_815 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_45 = _RAND_815[1:0];
  _RAND_816 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_46 = _RAND_816[1:0];
  _RAND_817 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_47 = _RAND_817[1:0];
  _RAND_818 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_48 = _RAND_818[1:0];
  _RAND_819 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_49 = _RAND_819[1:0];
  _RAND_820 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_50 = _RAND_820[1:0];
  _RAND_821 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_51 = _RAND_821[1:0];
  _RAND_822 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_52 = _RAND_822[1:0];
  _RAND_823 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_53 = _RAND_823[1:0];
  _RAND_824 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_54 = _RAND_824[1:0];
  _RAND_825 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_55 = _RAND_825[1:0];
  _RAND_826 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_56 = _RAND_826[1:0];
  _RAND_827 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_57 = _RAND_827[1:0];
  _RAND_828 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_58 = _RAND_828[1:0];
  _RAND_829 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_59 = _RAND_829[1:0];
  _RAND_830 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_60 = _RAND_830[1:0];
  _RAND_831 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_61 = _RAND_831[1:0];
  _RAND_832 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_62 = _RAND_832[1:0];
  _RAND_833 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_63 = _RAND_833[1:0];
  _RAND_834 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_64 = _RAND_834[1:0];
  _RAND_835 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_65 = _RAND_835[1:0];
  _RAND_836 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_66 = _RAND_836[1:0];
  _RAND_837 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_67 = _RAND_837[1:0];
  _RAND_838 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_68 = _RAND_838[1:0];
  _RAND_839 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_69 = _RAND_839[1:0];
  _RAND_840 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_70 = _RAND_840[1:0];
  _RAND_841 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_71 = _RAND_841[1:0];
  _RAND_842 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_72 = _RAND_842[1:0];
  _RAND_843 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_73 = _RAND_843[1:0];
  _RAND_844 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_74 = _RAND_844[1:0];
  _RAND_845 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_75 = _RAND_845[1:0];
  _RAND_846 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_76 = _RAND_846[1:0];
  _RAND_847 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_77 = _RAND_847[1:0];
  _RAND_848 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_78 = _RAND_848[1:0];
  _RAND_849 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_79 = _RAND_849[1:0];
  _RAND_850 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_80 = _RAND_850[1:0];
  _RAND_851 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_81 = _RAND_851[1:0];
  _RAND_852 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_82 = _RAND_852[1:0];
  _RAND_853 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_83 = _RAND_853[1:0];
  _RAND_854 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_84 = _RAND_854[1:0];
  _RAND_855 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_85 = _RAND_855[1:0];
  _RAND_856 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_86 = _RAND_856[1:0];
  _RAND_857 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_87 = _RAND_857[1:0];
  _RAND_858 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_88 = _RAND_858[1:0];
  _RAND_859 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_89 = _RAND_859[1:0];
  _RAND_860 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_90 = _RAND_860[1:0];
  _RAND_861 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_91 = _RAND_861[1:0];
  _RAND_862 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_92 = _RAND_862[1:0];
  _RAND_863 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_93 = _RAND_863[1:0];
  _RAND_864 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_94 = _RAND_864[1:0];
  _RAND_865 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_95 = _RAND_865[1:0];
  _RAND_866 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_96 = _RAND_866[1:0];
  _RAND_867 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_97 = _RAND_867[1:0];
  _RAND_868 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_98 = _RAND_868[1:0];
  _RAND_869 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_99 = _RAND_869[1:0];
  _RAND_870 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_100 = _RAND_870[1:0];
  _RAND_871 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_101 = _RAND_871[1:0];
  _RAND_872 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_102 = _RAND_872[1:0];
  _RAND_873 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_103 = _RAND_873[1:0];
  _RAND_874 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_104 = _RAND_874[1:0];
  _RAND_875 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_105 = _RAND_875[1:0];
  _RAND_876 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_106 = _RAND_876[1:0];
  _RAND_877 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_107 = _RAND_877[1:0];
  _RAND_878 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_108 = _RAND_878[1:0];
  _RAND_879 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_109 = _RAND_879[1:0];
  _RAND_880 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_110 = _RAND_880[1:0];
  _RAND_881 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_111 = _RAND_881[1:0];
  _RAND_882 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_112 = _RAND_882[1:0];
  _RAND_883 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_113 = _RAND_883[1:0];
  _RAND_884 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_114 = _RAND_884[1:0];
  _RAND_885 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_115 = _RAND_885[1:0];
  _RAND_886 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_116 = _RAND_886[1:0];
  _RAND_887 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_117 = _RAND_887[1:0];
  _RAND_888 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_118 = _RAND_888[1:0];
  _RAND_889 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_119 = _RAND_889[1:0];
  _RAND_890 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_120 = _RAND_890[1:0];
  _RAND_891 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_121 = _RAND_891[1:0];
  _RAND_892 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_122 = _RAND_892[1:0];
  _RAND_893 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_123 = _RAND_893[1:0];
  _RAND_894 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_124 = _RAND_894[1:0];
  _RAND_895 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_125 = _RAND_895[1:0];
  _RAND_896 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_126 = _RAND_896[1:0];
  _RAND_897 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_127 = _RAND_897[1:0];
  _RAND_898 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_128 = _RAND_898[1:0];
  _RAND_899 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_129 = _RAND_899[1:0];
  _RAND_900 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_130 = _RAND_900[1:0];
  _RAND_901 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_131 = _RAND_901[1:0];
  _RAND_902 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_132 = _RAND_902[1:0];
  _RAND_903 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_133 = _RAND_903[1:0];
  _RAND_904 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_134 = _RAND_904[1:0];
  _RAND_905 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_135 = _RAND_905[1:0];
  _RAND_906 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_136 = _RAND_906[1:0];
  _RAND_907 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_137 = _RAND_907[1:0];
  _RAND_908 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_138 = _RAND_908[1:0];
  _RAND_909 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_139 = _RAND_909[1:0];
  _RAND_910 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_140 = _RAND_910[1:0];
  _RAND_911 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_141 = _RAND_911[1:0];
  _RAND_912 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_142 = _RAND_912[1:0];
  _RAND_913 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_143 = _RAND_913[1:0];
  _RAND_914 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_144 = _RAND_914[1:0];
  _RAND_915 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_145 = _RAND_915[1:0];
  _RAND_916 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_146 = _RAND_916[1:0];
  _RAND_917 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_147 = _RAND_917[1:0];
  _RAND_918 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_148 = _RAND_918[1:0];
  _RAND_919 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_149 = _RAND_919[1:0];
  _RAND_920 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_150 = _RAND_920[1:0];
  _RAND_921 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_151 = _RAND_921[1:0];
  _RAND_922 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_152 = _RAND_922[1:0];
  _RAND_923 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_153 = _RAND_923[1:0];
  _RAND_924 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_154 = _RAND_924[1:0];
  _RAND_925 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_155 = _RAND_925[1:0];
  _RAND_926 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_156 = _RAND_926[1:0];
  _RAND_927 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_157 = _RAND_927[1:0];
  _RAND_928 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_158 = _RAND_928[1:0];
  _RAND_929 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_159 = _RAND_929[1:0];
  _RAND_930 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_160 = _RAND_930[1:0];
  _RAND_931 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_161 = _RAND_931[1:0];
  _RAND_932 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_162 = _RAND_932[1:0];
  _RAND_933 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_163 = _RAND_933[1:0];
  _RAND_934 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_164 = _RAND_934[1:0];
  _RAND_935 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_165 = _RAND_935[1:0];
  _RAND_936 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_166 = _RAND_936[1:0];
  _RAND_937 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_167 = _RAND_937[1:0];
  _RAND_938 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_168 = _RAND_938[1:0];
  _RAND_939 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_169 = _RAND_939[1:0];
  _RAND_940 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_170 = _RAND_940[1:0];
  _RAND_941 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_171 = _RAND_941[1:0];
  _RAND_942 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_172 = _RAND_942[1:0];
  _RAND_943 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_173 = _RAND_943[1:0];
  _RAND_944 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_174 = _RAND_944[1:0];
  _RAND_945 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_175 = _RAND_945[1:0];
  _RAND_946 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_176 = _RAND_946[1:0];
  _RAND_947 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_177 = _RAND_947[1:0];
  _RAND_948 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_178 = _RAND_948[1:0];
  _RAND_949 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_179 = _RAND_949[1:0];
  _RAND_950 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_180 = _RAND_950[1:0];
  _RAND_951 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_181 = _RAND_951[1:0];
  _RAND_952 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_182 = _RAND_952[1:0];
  _RAND_953 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_183 = _RAND_953[1:0];
  _RAND_954 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_184 = _RAND_954[1:0];
  _RAND_955 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_185 = _RAND_955[1:0];
  _RAND_956 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_186 = _RAND_956[1:0];
  _RAND_957 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_187 = _RAND_957[1:0];
  _RAND_958 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_188 = _RAND_958[1:0];
  _RAND_959 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_189 = _RAND_959[1:0];
  _RAND_960 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_190 = _RAND_960[1:0];
  _RAND_961 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_191 = _RAND_961[1:0];
  _RAND_962 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_192 = _RAND_962[1:0];
  _RAND_963 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_193 = _RAND_963[1:0];
  _RAND_964 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_194 = _RAND_964[1:0];
  _RAND_965 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_195 = _RAND_965[1:0];
  _RAND_966 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_196 = _RAND_966[1:0];
  _RAND_967 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_197 = _RAND_967[1:0];
  _RAND_968 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_198 = _RAND_968[1:0];
  _RAND_969 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_199 = _RAND_969[1:0];
  _RAND_970 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_200 = _RAND_970[1:0];
  _RAND_971 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_201 = _RAND_971[1:0];
  _RAND_972 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_202 = _RAND_972[1:0];
  _RAND_973 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_203 = _RAND_973[1:0];
  _RAND_974 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_204 = _RAND_974[1:0];
  _RAND_975 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_205 = _RAND_975[1:0];
  _RAND_976 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_206 = _RAND_976[1:0];
  _RAND_977 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_207 = _RAND_977[1:0];
  _RAND_978 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_208 = _RAND_978[1:0];
  _RAND_979 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_209 = _RAND_979[1:0];
  _RAND_980 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_210 = _RAND_980[1:0];
  _RAND_981 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_211 = _RAND_981[1:0];
  _RAND_982 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_212 = _RAND_982[1:0];
  _RAND_983 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_213 = _RAND_983[1:0];
  _RAND_984 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_214 = _RAND_984[1:0];
  _RAND_985 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_215 = _RAND_985[1:0];
  _RAND_986 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_216 = _RAND_986[1:0];
  _RAND_987 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_217 = _RAND_987[1:0];
  _RAND_988 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_218 = _RAND_988[1:0];
  _RAND_989 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_219 = _RAND_989[1:0];
  _RAND_990 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_220 = _RAND_990[1:0];
  _RAND_991 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_221 = _RAND_991[1:0];
  _RAND_992 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_222 = _RAND_992[1:0];
  _RAND_993 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_223 = _RAND_993[1:0];
  _RAND_994 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_224 = _RAND_994[1:0];
  _RAND_995 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_225 = _RAND_995[1:0];
  _RAND_996 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_226 = _RAND_996[1:0];
  _RAND_997 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_227 = _RAND_997[1:0];
  _RAND_998 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_228 = _RAND_998[1:0];
  _RAND_999 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_229 = _RAND_999[1:0];
  _RAND_1000 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_230 = _RAND_1000[1:0];
  _RAND_1001 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_231 = _RAND_1001[1:0];
  _RAND_1002 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_232 = _RAND_1002[1:0];
  _RAND_1003 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_233 = _RAND_1003[1:0];
  _RAND_1004 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_234 = _RAND_1004[1:0];
  _RAND_1005 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_235 = _RAND_1005[1:0];
  _RAND_1006 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_236 = _RAND_1006[1:0];
  _RAND_1007 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_237 = _RAND_1007[1:0];
  _RAND_1008 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_238 = _RAND_1008[1:0];
  _RAND_1009 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_239 = _RAND_1009[1:0];
  _RAND_1010 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_240 = _RAND_1010[1:0];
  _RAND_1011 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_241 = _RAND_1011[1:0];
  _RAND_1012 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_242 = _RAND_1012[1:0];
  _RAND_1013 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_243 = _RAND_1013[1:0];
  _RAND_1014 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_244 = _RAND_1014[1:0];
  _RAND_1015 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_245 = _RAND_1015[1:0];
  _RAND_1016 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_246 = _RAND_1016[1:0];
  _RAND_1017 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_247 = _RAND_1017[1:0];
  _RAND_1018 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_248 = _RAND_1018[1:0];
  _RAND_1019 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_249 = _RAND_1019[1:0];
  _RAND_1020 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_250 = _RAND_1020[1:0];
  _RAND_1021 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_251 = _RAND_1021[1:0];
  _RAND_1022 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_252 = _RAND_1022[1:0];
  _RAND_1023 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_253 = _RAND_1023[1:0];
  _RAND_1024 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_254 = _RAND_1024[1:0];
  _RAND_1025 = {1{`RANDOM}};
  bht_bank_rd_data_out_0_255 = _RAND_1025[1:0];
  _RAND_1026 = {1{`RANDOM}};
  exu_mp_way_f = _RAND_1026[0:0];
  _RAND_1027 = {8{`RANDOM}};
  btb_lru_b0_f = _RAND_1027[255:0];
  _RAND_1028 = {1{`RANDOM}};
  exu_flush_final_d1 = _RAND_1028[0:0];
  _RAND_1029 = {1{`RANDOM}};
  ifc_fetch_adder_prior = _RAND_1029[29:0];
  _RAND_1030 = {1{`RANDOM}};
  rets_out_0 = _RAND_1030[31:0];
  _RAND_1031 = {1{`RANDOM}};
  rets_out_1 = _RAND_1031[31:0];
  _RAND_1032 = {1{`RANDOM}};
  rets_out_2 = _RAND_1032[31:0];
  _RAND_1033 = {1{`RANDOM}};
  rets_out_3 = _RAND_1033[31:0];
  _RAND_1034 = {1{`RANDOM}};
  rets_out_4 = _RAND_1034[31:0];
  _RAND_1035 = {1{`RANDOM}};
  rets_out_5 = _RAND_1035[31:0];
  _RAND_1036 = {1{`RANDOM}};
  rets_out_6 = _RAND_1036[31:0];
  _RAND_1037 = {1{`RANDOM}};
  rets_out_7 = _RAND_1037[31:0];
`endif // RANDOMIZE_REG_INIT
  if (reset) begin
    leak_one_f_d1 = 1'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way0_out_255 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_0 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_1 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_2 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_3 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_4 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_5 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_6 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_7 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_8 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_9 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_10 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_11 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_12 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_13 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_14 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_15 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_16 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_17 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_18 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_19 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_20 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_21 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_22 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_23 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_24 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_25 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_26 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_27 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_28 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_29 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_30 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_31 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_32 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_33 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_34 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_35 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_36 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_37 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_38 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_39 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_40 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_41 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_42 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_43 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_44 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_45 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_46 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_47 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_48 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_49 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_50 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_51 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_52 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_53 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_54 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_55 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_56 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_57 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_58 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_59 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_60 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_61 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_62 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_63 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_64 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_65 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_66 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_67 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_68 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_69 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_70 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_71 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_72 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_73 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_74 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_75 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_76 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_77 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_78 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_79 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_80 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_81 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_82 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_83 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_84 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_85 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_86 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_87 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_88 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_89 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_90 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_91 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_92 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_93 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_94 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_95 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_96 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_97 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_98 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_99 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_100 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_101 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_102 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_103 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_104 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_105 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_106 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_107 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_108 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_109 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_110 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_111 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_112 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_113 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_114 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_115 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_116 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_117 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_118 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_119 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_120 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_121 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_122 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_123 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_124 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_125 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_126 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_127 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_128 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_129 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_130 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_131 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_132 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_133 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_134 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_135 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_136 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_137 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_138 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_139 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_140 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_141 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_142 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_143 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_144 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_145 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_146 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_147 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_148 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_149 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_150 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_151 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_152 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_153 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_154 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_155 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_156 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_157 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_158 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_159 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_160 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_161 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_162 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_163 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_164 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_165 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_166 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_167 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_168 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_169 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_170 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_171 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_172 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_173 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_174 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_175 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_176 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_177 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_178 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_179 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_180 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_181 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_182 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_183 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_184 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_185 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_186 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_187 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_188 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_189 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_190 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_191 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_192 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_193 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_194 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_195 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_196 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_197 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_198 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_199 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_200 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_201 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_202 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_203 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_204 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_205 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_206 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_207 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_208 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_209 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_210 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_211 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_212 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_213 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_214 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_215 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_216 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_217 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_218 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_219 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_220 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_221 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_222 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_223 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_224 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_225 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_226 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_227 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_228 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_229 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_230 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_231 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_232 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_233 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_234 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_235 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_236 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_237 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_238 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_239 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_240 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_241 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_242 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_243 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_244 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_245 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_246 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_247 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_248 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_249 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_250 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_251 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_252 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_253 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_254 = 22'h0;
  end
  if (reset) begin
    btb_bank0_rd_data_way1_out_255 = 22'h0;
  end
  if (reset) begin
    fghr = 8'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_1_255 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_0 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_1 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_2 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_3 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_4 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_5 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_6 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_7 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_8 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_9 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_10 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_11 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_12 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_13 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_14 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_15 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_16 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_17 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_18 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_19 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_20 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_21 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_22 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_23 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_24 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_25 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_26 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_27 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_28 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_29 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_30 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_31 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_32 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_33 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_34 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_35 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_36 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_37 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_38 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_39 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_40 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_41 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_42 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_43 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_44 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_45 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_46 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_47 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_48 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_49 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_50 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_51 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_52 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_53 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_54 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_55 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_56 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_57 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_58 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_59 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_60 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_61 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_62 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_63 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_64 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_65 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_66 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_67 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_68 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_69 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_70 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_71 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_72 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_73 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_74 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_75 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_76 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_77 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_78 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_79 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_80 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_81 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_82 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_83 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_84 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_85 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_86 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_87 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_88 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_89 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_90 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_91 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_92 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_93 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_94 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_95 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_96 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_97 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_98 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_99 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_100 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_101 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_102 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_103 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_104 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_105 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_106 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_107 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_108 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_109 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_110 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_111 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_112 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_113 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_114 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_115 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_116 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_117 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_118 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_119 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_120 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_121 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_122 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_123 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_124 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_125 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_126 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_127 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_128 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_129 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_130 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_131 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_132 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_133 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_134 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_135 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_136 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_137 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_138 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_139 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_140 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_141 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_142 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_143 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_144 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_145 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_146 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_147 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_148 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_149 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_150 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_151 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_152 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_153 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_154 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_155 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_156 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_157 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_158 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_159 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_160 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_161 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_162 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_163 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_164 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_165 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_166 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_167 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_168 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_169 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_170 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_171 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_172 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_173 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_174 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_175 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_176 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_177 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_178 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_179 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_180 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_181 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_182 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_183 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_184 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_185 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_186 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_187 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_188 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_189 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_190 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_191 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_192 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_193 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_194 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_195 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_196 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_197 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_198 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_199 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_200 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_201 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_202 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_203 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_204 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_205 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_206 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_207 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_208 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_209 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_210 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_211 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_212 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_213 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_214 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_215 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_216 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_217 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_218 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_219 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_220 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_221 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_222 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_223 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_224 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_225 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_226 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_227 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_228 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_229 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_230 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_231 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_232 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_233 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_234 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_235 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_236 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_237 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_238 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_239 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_240 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_241 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_242 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_243 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_244 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_245 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_246 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_247 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_248 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_249 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_250 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_251 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_252 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_253 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_254 = 2'h0;
  end
  if (reset) begin
    bht_bank_rd_data_out_0_255 = 2'h0;
  end
  if (reset) begin
    exu_mp_way_f = 1'h0;
  end
  if (reset) begin
    btb_lru_b0_f = 256'h0;
  end
  if (reset) begin
    exu_flush_final_d1 = 1'h0;
  end
  if (reset) begin
    ifc_fetch_adder_prior = 30'h0;
  end
  if (reset) begin
    rets_out_0 = 32'h0;
  end
  if (reset) begin
    rets_out_1 = 32'h0;
  end
  if (reset) begin
    rets_out_2 = 32'h0;
  end
  if (reset) begin
    rets_out_3 = 32'h0;
  end
  if (reset) begin
    rets_out_4 = 32'h0;
  end
  if (reset) begin
    rets_out_5 = 32'h0;
  end
  if (reset) begin
    rets_out_6 = 32'h0;
  end
  if (reset) begin
    rets_out_7 = 32'h0;
  end
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      leak_one_f_d1 <= 1'h0;
    end else if (_T_337) begin
      leak_one_f_d1 <= leak_one_f;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_0 <= 22'h0;
    end else if (_T_614) begin
      btb_bank0_rd_data_way0_out_0 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_1 <= 22'h0;
    end else if (_T_618) begin
      btb_bank0_rd_data_way0_out_1 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_2 <= 22'h0;
    end else if (_T_622) begin
      btb_bank0_rd_data_way0_out_2 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_3 <= 22'h0;
    end else if (_T_626) begin
      btb_bank0_rd_data_way0_out_3 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_4 <= 22'h0;
    end else if (_T_630) begin
      btb_bank0_rd_data_way0_out_4 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_5 <= 22'h0;
    end else if (_T_634) begin
      btb_bank0_rd_data_way0_out_5 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_6 <= 22'h0;
    end else if (_T_638) begin
      btb_bank0_rd_data_way0_out_6 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_7 <= 22'h0;
    end else if (_T_642) begin
      btb_bank0_rd_data_way0_out_7 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_8 <= 22'h0;
    end else if (_T_646) begin
      btb_bank0_rd_data_way0_out_8 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_9 <= 22'h0;
    end else if (_T_650) begin
      btb_bank0_rd_data_way0_out_9 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_10 <= 22'h0;
    end else if (_T_654) begin
      btb_bank0_rd_data_way0_out_10 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_11 <= 22'h0;
    end else if (_T_658) begin
      btb_bank0_rd_data_way0_out_11 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_12 <= 22'h0;
    end else if (_T_662) begin
      btb_bank0_rd_data_way0_out_12 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_13 <= 22'h0;
    end else if (_T_666) begin
      btb_bank0_rd_data_way0_out_13 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_14 <= 22'h0;
    end else if (_T_670) begin
      btb_bank0_rd_data_way0_out_14 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_15 <= 22'h0;
    end else if (_T_674) begin
      btb_bank0_rd_data_way0_out_15 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_16 <= 22'h0;
    end else if (_T_678) begin
      btb_bank0_rd_data_way0_out_16 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_17 <= 22'h0;
    end else if (_T_682) begin
      btb_bank0_rd_data_way0_out_17 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_18 <= 22'h0;
    end else if (_T_686) begin
      btb_bank0_rd_data_way0_out_18 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_19 <= 22'h0;
    end else if (_T_690) begin
      btb_bank0_rd_data_way0_out_19 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_20 <= 22'h0;
    end else if (_T_694) begin
      btb_bank0_rd_data_way0_out_20 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_21 <= 22'h0;
    end else if (_T_698) begin
      btb_bank0_rd_data_way0_out_21 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_22 <= 22'h0;
    end else if (_T_702) begin
      btb_bank0_rd_data_way0_out_22 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_23 <= 22'h0;
    end else if (_T_706) begin
      btb_bank0_rd_data_way0_out_23 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_24 <= 22'h0;
    end else if (_T_710) begin
      btb_bank0_rd_data_way0_out_24 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_25 <= 22'h0;
    end else if (_T_714) begin
      btb_bank0_rd_data_way0_out_25 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_26 <= 22'h0;
    end else if (_T_718) begin
      btb_bank0_rd_data_way0_out_26 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_27 <= 22'h0;
    end else if (_T_722) begin
      btb_bank0_rd_data_way0_out_27 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_28 <= 22'h0;
    end else if (_T_726) begin
      btb_bank0_rd_data_way0_out_28 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_29 <= 22'h0;
    end else if (_T_730) begin
      btb_bank0_rd_data_way0_out_29 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_30 <= 22'h0;
    end else if (_T_734) begin
      btb_bank0_rd_data_way0_out_30 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_31 <= 22'h0;
    end else if (_T_738) begin
      btb_bank0_rd_data_way0_out_31 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_32 <= 22'h0;
    end else if (_T_742) begin
      btb_bank0_rd_data_way0_out_32 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_33 <= 22'h0;
    end else if (_T_746) begin
      btb_bank0_rd_data_way0_out_33 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_34 <= 22'h0;
    end else if (_T_750) begin
      btb_bank0_rd_data_way0_out_34 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_35 <= 22'h0;
    end else if (_T_754) begin
      btb_bank0_rd_data_way0_out_35 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_36 <= 22'h0;
    end else if (_T_758) begin
      btb_bank0_rd_data_way0_out_36 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_37 <= 22'h0;
    end else if (_T_762) begin
      btb_bank0_rd_data_way0_out_37 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_38 <= 22'h0;
    end else if (_T_766) begin
      btb_bank0_rd_data_way0_out_38 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_39 <= 22'h0;
    end else if (_T_770) begin
      btb_bank0_rd_data_way0_out_39 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_40 <= 22'h0;
    end else if (_T_774) begin
      btb_bank0_rd_data_way0_out_40 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_41 <= 22'h0;
    end else if (_T_778) begin
      btb_bank0_rd_data_way0_out_41 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_42 <= 22'h0;
    end else if (_T_782) begin
      btb_bank0_rd_data_way0_out_42 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_43 <= 22'h0;
    end else if (_T_786) begin
      btb_bank0_rd_data_way0_out_43 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_44 <= 22'h0;
    end else if (_T_790) begin
      btb_bank0_rd_data_way0_out_44 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_45 <= 22'h0;
    end else if (_T_794) begin
      btb_bank0_rd_data_way0_out_45 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_46 <= 22'h0;
    end else if (_T_798) begin
      btb_bank0_rd_data_way0_out_46 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_47 <= 22'h0;
    end else if (_T_802) begin
      btb_bank0_rd_data_way0_out_47 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_48 <= 22'h0;
    end else if (_T_806) begin
      btb_bank0_rd_data_way0_out_48 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_49 <= 22'h0;
    end else if (_T_810) begin
      btb_bank0_rd_data_way0_out_49 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_50 <= 22'h0;
    end else if (_T_814) begin
      btb_bank0_rd_data_way0_out_50 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_51 <= 22'h0;
    end else if (_T_818) begin
      btb_bank0_rd_data_way0_out_51 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_52 <= 22'h0;
    end else if (_T_822) begin
      btb_bank0_rd_data_way0_out_52 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_53 <= 22'h0;
    end else if (_T_826) begin
      btb_bank0_rd_data_way0_out_53 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_54 <= 22'h0;
    end else if (_T_830) begin
      btb_bank0_rd_data_way0_out_54 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_55 <= 22'h0;
    end else if (_T_834) begin
      btb_bank0_rd_data_way0_out_55 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_56 <= 22'h0;
    end else if (_T_838) begin
      btb_bank0_rd_data_way0_out_56 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_57 <= 22'h0;
    end else if (_T_842) begin
      btb_bank0_rd_data_way0_out_57 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_58 <= 22'h0;
    end else if (_T_846) begin
      btb_bank0_rd_data_way0_out_58 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_59 <= 22'h0;
    end else if (_T_850) begin
      btb_bank0_rd_data_way0_out_59 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_60 <= 22'h0;
    end else if (_T_854) begin
      btb_bank0_rd_data_way0_out_60 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_61 <= 22'h0;
    end else if (_T_858) begin
      btb_bank0_rd_data_way0_out_61 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_62 <= 22'h0;
    end else if (_T_862) begin
      btb_bank0_rd_data_way0_out_62 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_63 <= 22'h0;
    end else if (_T_866) begin
      btb_bank0_rd_data_way0_out_63 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_64 <= 22'h0;
    end else if (_T_870) begin
      btb_bank0_rd_data_way0_out_64 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_65 <= 22'h0;
    end else if (_T_874) begin
      btb_bank0_rd_data_way0_out_65 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_66 <= 22'h0;
    end else if (_T_878) begin
      btb_bank0_rd_data_way0_out_66 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_67 <= 22'h0;
    end else if (_T_882) begin
      btb_bank0_rd_data_way0_out_67 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_68 <= 22'h0;
    end else if (_T_886) begin
      btb_bank0_rd_data_way0_out_68 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_69 <= 22'h0;
    end else if (_T_890) begin
      btb_bank0_rd_data_way0_out_69 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_70 <= 22'h0;
    end else if (_T_894) begin
      btb_bank0_rd_data_way0_out_70 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_71 <= 22'h0;
    end else if (_T_898) begin
      btb_bank0_rd_data_way0_out_71 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_72 <= 22'h0;
    end else if (_T_902) begin
      btb_bank0_rd_data_way0_out_72 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_73 <= 22'h0;
    end else if (_T_906) begin
      btb_bank0_rd_data_way0_out_73 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_74 <= 22'h0;
    end else if (_T_910) begin
      btb_bank0_rd_data_way0_out_74 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_75 <= 22'h0;
    end else if (_T_914) begin
      btb_bank0_rd_data_way0_out_75 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_76 <= 22'h0;
    end else if (_T_918) begin
      btb_bank0_rd_data_way0_out_76 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_77 <= 22'h0;
    end else if (_T_922) begin
      btb_bank0_rd_data_way0_out_77 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_78 <= 22'h0;
    end else if (_T_926) begin
      btb_bank0_rd_data_way0_out_78 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_79 <= 22'h0;
    end else if (_T_930) begin
      btb_bank0_rd_data_way0_out_79 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_80 <= 22'h0;
    end else if (_T_934) begin
      btb_bank0_rd_data_way0_out_80 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_81 <= 22'h0;
    end else if (_T_938) begin
      btb_bank0_rd_data_way0_out_81 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_82 <= 22'h0;
    end else if (_T_942) begin
      btb_bank0_rd_data_way0_out_82 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_83 <= 22'h0;
    end else if (_T_946) begin
      btb_bank0_rd_data_way0_out_83 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_84 <= 22'h0;
    end else if (_T_950) begin
      btb_bank0_rd_data_way0_out_84 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_85 <= 22'h0;
    end else if (_T_954) begin
      btb_bank0_rd_data_way0_out_85 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_86 <= 22'h0;
    end else if (_T_958) begin
      btb_bank0_rd_data_way0_out_86 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_87 <= 22'h0;
    end else if (_T_962) begin
      btb_bank0_rd_data_way0_out_87 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_88 <= 22'h0;
    end else if (_T_966) begin
      btb_bank0_rd_data_way0_out_88 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_89 <= 22'h0;
    end else if (_T_970) begin
      btb_bank0_rd_data_way0_out_89 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_90 <= 22'h0;
    end else if (_T_974) begin
      btb_bank0_rd_data_way0_out_90 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_91 <= 22'h0;
    end else if (_T_978) begin
      btb_bank0_rd_data_way0_out_91 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_92 <= 22'h0;
    end else if (_T_982) begin
      btb_bank0_rd_data_way0_out_92 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_93 <= 22'h0;
    end else if (_T_986) begin
      btb_bank0_rd_data_way0_out_93 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_94 <= 22'h0;
    end else if (_T_990) begin
      btb_bank0_rd_data_way0_out_94 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_95 <= 22'h0;
    end else if (_T_994) begin
      btb_bank0_rd_data_way0_out_95 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_96 <= 22'h0;
    end else if (_T_998) begin
      btb_bank0_rd_data_way0_out_96 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_97 <= 22'h0;
    end else if (_T_1002) begin
      btb_bank0_rd_data_way0_out_97 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_98 <= 22'h0;
    end else if (_T_1006) begin
      btb_bank0_rd_data_way0_out_98 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_99 <= 22'h0;
    end else if (_T_1010) begin
      btb_bank0_rd_data_way0_out_99 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_100 <= 22'h0;
    end else if (_T_1014) begin
      btb_bank0_rd_data_way0_out_100 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_101 <= 22'h0;
    end else if (_T_1018) begin
      btb_bank0_rd_data_way0_out_101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_102 <= 22'h0;
    end else if (_T_1022) begin
      btb_bank0_rd_data_way0_out_102 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_103 <= 22'h0;
    end else if (_T_1026) begin
      btb_bank0_rd_data_way0_out_103 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_104 <= 22'h0;
    end else if (_T_1030) begin
      btb_bank0_rd_data_way0_out_104 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_105 <= 22'h0;
    end else if (_T_1034) begin
      btb_bank0_rd_data_way0_out_105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_106 <= 22'h0;
    end else if (_T_1038) begin
      btb_bank0_rd_data_way0_out_106 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_107 <= 22'h0;
    end else if (_T_1042) begin
      btb_bank0_rd_data_way0_out_107 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_108 <= 22'h0;
    end else if (_T_1046) begin
      btb_bank0_rd_data_way0_out_108 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_109 <= 22'h0;
    end else if (_T_1050) begin
      btb_bank0_rd_data_way0_out_109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_110 <= 22'h0;
    end else if (_T_1054) begin
      btb_bank0_rd_data_way0_out_110 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_111 <= 22'h0;
    end else if (_T_1058) begin
      btb_bank0_rd_data_way0_out_111 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_112 <= 22'h0;
    end else if (_T_1062) begin
      btb_bank0_rd_data_way0_out_112 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_113 <= 22'h0;
    end else if (_T_1066) begin
      btb_bank0_rd_data_way0_out_113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_114 <= 22'h0;
    end else if (_T_1070) begin
      btb_bank0_rd_data_way0_out_114 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_115 <= 22'h0;
    end else if (_T_1074) begin
      btb_bank0_rd_data_way0_out_115 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_116 <= 22'h0;
    end else if (_T_1078) begin
      btb_bank0_rd_data_way0_out_116 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_117 <= 22'h0;
    end else if (_T_1082) begin
      btb_bank0_rd_data_way0_out_117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_118 <= 22'h0;
    end else if (_T_1086) begin
      btb_bank0_rd_data_way0_out_118 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_119 <= 22'h0;
    end else if (_T_1090) begin
      btb_bank0_rd_data_way0_out_119 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_120 <= 22'h0;
    end else if (_T_1094) begin
      btb_bank0_rd_data_way0_out_120 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_121 <= 22'h0;
    end else if (_T_1098) begin
      btb_bank0_rd_data_way0_out_121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_122 <= 22'h0;
    end else if (_T_1102) begin
      btb_bank0_rd_data_way0_out_122 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_123 <= 22'h0;
    end else if (_T_1106) begin
      btb_bank0_rd_data_way0_out_123 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_124 <= 22'h0;
    end else if (_T_1110) begin
      btb_bank0_rd_data_way0_out_124 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_125 <= 22'h0;
    end else if (_T_1114) begin
      btb_bank0_rd_data_way0_out_125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_126 <= 22'h0;
    end else if (_T_1118) begin
      btb_bank0_rd_data_way0_out_126 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_127 <= 22'h0;
    end else if (_T_1122) begin
      btb_bank0_rd_data_way0_out_127 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_128 <= 22'h0;
    end else if (_T_1126) begin
      btb_bank0_rd_data_way0_out_128 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_129 <= 22'h0;
    end else if (_T_1130) begin
      btb_bank0_rd_data_way0_out_129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_130 <= 22'h0;
    end else if (_T_1134) begin
      btb_bank0_rd_data_way0_out_130 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_131 <= 22'h0;
    end else if (_T_1138) begin
      btb_bank0_rd_data_way0_out_131 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_132 <= 22'h0;
    end else if (_T_1142) begin
      btb_bank0_rd_data_way0_out_132 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_133 <= 22'h0;
    end else if (_T_1146) begin
      btb_bank0_rd_data_way0_out_133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_134 <= 22'h0;
    end else if (_T_1150) begin
      btb_bank0_rd_data_way0_out_134 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_135 <= 22'h0;
    end else if (_T_1154) begin
      btb_bank0_rd_data_way0_out_135 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_136 <= 22'h0;
    end else if (_T_1158) begin
      btb_bank0_rd_data_way0_out_136 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_137 <= 22'h0;
    end else if (_T_1162) begin
      btb_bank0_rd_data_way0_out_137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_138 <= 22'h0;
    end else if (_T_1166) begin
      btb_bank0_rd_data_way0_out_138 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_139 <= 22'h0;
    end else if (_T_1170) begin
      btb_bank0_rd_data_way0_out_139 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_140 <= 22'h0;
    end else if (_T_1174) begin
      btb_bank0_rd_data_way0_out_140 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_141 <= 22'h0;
    end else if (_T_1178) begin
      btb_bank0_rd_data_way0_out_141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_142 <= 22'h0;
    end else if (_T_1182) begin
      btb_bank0_rd_data_way0_out_142 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_143 <= 22'h0;
    end else if (_T_1186) begin
      btb_bank0_rd_data_way0_out_143 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_144 <= 22'h0;
    end else if (_T_1190) begin
      btb_bank0_rd_data_way0_out_144 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_145 <= 22'h0;
    end else if (_T_1194) begin
      btb_bank0_rd_data_way0_out_145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_146 <= 22'h0;
    end else if (_T_1198) begin
      btb_bank0_rd_data_way0_out_146 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_147 <= 22'h0;
    end else if (_T_1202) begin
      btb_bank0_rd_data_way0_out_147 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_148 <= 22'h0;
    end else if (_T_1206) begin
      btb_bank0_rd_data_way0_out_148 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_149 <= 22'h0;
    end else if (_T_1210) begin
      btb_bank0_rd_data_way0_out_149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_150 <= 22'h0;
    end else if (_T_1214) begin
      btb_bank0_rd_data_way0_out_150 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_151 <= 22'h0;
    end else if (_T_1218) begin
      btb_bank0_rd_data_way0_out_151 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_152 <= 22'h0;
    end else if (_T_1222) begin
      btb_bank0_rd_data_way0_out_152 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_153 <= 22'h0;
    end else if (_T_1226) begin
      btb_bank0_rd_data_way0_out_153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_154 <= 22'h0;
    end else if (_T_1230) begin
      btb_bank0_rd_data_way0_out_154 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_155 <= 22'h0;
    end else if (_T_1234) begin
      btb_bank0_rd_data_way0_out_155 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_156 <= 22'h0;
    end else if (_T_1238) begin
      btb_bank0_rd_data_way0_out_156 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_157 <= 22'h0;
    end else if (_T_1242) begin
      btb_bank0_rd_data_way0_out_157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_158 <= 22'h0;
    end else if (_T_1246) begin
      btb_bank0_rd_data_way0_out_158 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_159 <= 22'h0;
    end else if (_T_1250) begin
      btb_bank0_rd_data_way0_out_159 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_160 <= 22'h0;
    end else if (_T_1254) begin
      btb_bank0_rd_data_way0_out_160 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_161 <= 22'h0;
    end else if (_T_1258) begin
      btb_bank0_rd_data_way0_out_161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_162 <= 22'h0;
    end else if (_T_1262) begin
      btb_bank0_rd_data_way0_out_162 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_163 <= 22'h0;
    end else if (_T_1266) begin
      btb_bank0_rd_data_way0_out_163 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_164 <= 22'h0;
    end else if (_T_1270) begin
      btb_bank0_rd_data_way0_out_164 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_165 <= 22'h0;
    end else if (_T_1274) begin
      btb_bank0_rd_data_way0_out_165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_166 <= 22'h0;
    end else if (_T_1278) begin
      btb_bank0_rd_data_way0_out_166 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_167 <= 22'h0;
    end else if (_T_1282) begin
      btb_bank0_rd_data_way0_out_167 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_168 <= 22'h0;
    end else if (_T_1286) begin
      btb_bank0_rd_data_way0_out_168 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_169 <= 22'h0;
    end else if (_T_1290) begin
      btb_bank0_rd_data_way0_out_169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_170 <= 22'h0;
    end else if (_T_1294) begin
      btb_bank0_rd_data_way0_out_170 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_171 <= 22'h0;
    end else if (_T_1298) begin
      btb_bank0_rd_data_way0_out_171 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_172 <= 22'h0;
    end else if (_T_1302) begin
      btb_bank0_rd_data_way0_out_172 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_173 <= 22'h0;
    end else if (_T_1306) begin
      btb_bank0_rd_data_way0_out_173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_174 <= 22'h0;
    end else if (_T_1310) begin
      btb_bank0_rd_data_way0_out_174 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_175 <= 22'h0;
    end else if (_T_1314) begin
      btb_bank0_rd_data_way0_out_175 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_176 <= 22'h0;
    end else if (_T_1318) begin
      btb_bank0_rd_data_way0_out_176 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_177 <= 22'h0;
    end else if (_T_1322) begin
      btb_bank0_rd_data_way0_out_177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_178 <= 22'h0;
    end else if (_T_1326) begin
      btb_bank0_rd_data_way0_out_178 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_179 <= 22'h0;
    end else if (_T_1330) begin
      btb_bank0_rd_data_way0_out_179 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_180 <= 22'h0;
    end else if (_T_1334) begin
      btb_bank0_rd_data_way0_out_180 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_181 <= 22'h0;
    end else if (_T_1338) begin
      btb_bank0_rd_data_way0_out_181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_182 <= 22'h0;
    end else if (_T_1342) begin
      btb_bank0_rd_data_way0_out_182 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_183 <= 22'h0;
    end else if (_T_1346) begin
      btb_bank0_rd_data_way0_out_183 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_184 <= 22'h0;
    end else if (_T_1350) begin
      btb_bank0_rd_data_way0_out_184 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_185 <= 22'h0;
    end else if (_T_1354) begin
      btb_bank0_rd_data_way0_out_185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_186 <= 22'h0;
    end else if (_T_1358) begin
      btb_bank0_rd_data_way0_out_186 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_187 <= 22'h0;
    end else if (_T_1362) begin
      btb_bank0_rd_data_way0_out_187 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_188 <= 22'h0;
    end else if (_T_1366) begin
      btb_bank0_rd_data_way0_out_188 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_189 <= 22'h0;
    end else if (_T_1370) begin
      btb_bank0_rd_data_way0_out_189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_190 <= 22'h0;
    end else if (_T_1374) begin
      btb_bank0_rd_data_way0_out_190 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_191 <= 22'h0;
    end else if (_T_1378) begin
      btb_bank0_rd_data_way0_out_191 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_192 <= 22'h0;
    end else if (_T_1382) begin
      btb_bank0_rd_data_way0_out_192 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_193 <= 22'h0;
    end else if (_T_1386) begin
      btb_bank0_rd_data_way0_out_193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_194 <= 22'h0;
    end else if (_T_1390) begin
      btb_bank0_rd_data_way0_out_194 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_195 <= 22'h0;
    end else if (_T_1394) begin
      btb_bank0_rd_data_way0_out_195 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_196 <= 22'h0;
    end else if (_T_1398) begin
      btb_bank0_rd_data_way0_out_196 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_197 <= 22'h0;
    end else if (_T_1402) begin
      btb_bank0_rd_data_way0_out_197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_198 <= 22'h0;
    end else if (_T_1406) begin
      btb_bank0_rd_data_way0_out_198 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_199 <= 22'h0;
    end else if (_T_1410) begin
      btb_bank0_rd_data_way0_out_199 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_200 <= 22'h0;
    end else if (_T_1414) begin
      btb_bank0_rd_data_way0_out_200 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_201 <= 22'h0;
    end else if (_T_1418) begin
      btb_bank0_rd_data_way0_out_201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_202 <= 22'h0;
    end else if (_T_1422) begin
      btb_bank0_rd_data_way0_out_202 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_203 <= 22'h0;
    end else if (_T_1426) begin
      btb_bank0_rd_data_way0_out_203 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_204 <= 22'h0;
    end else if (_T_1430) begin
      btb_bank0_rd_data_way0_out_204 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_205 <= 22'h0;
    end else if (_T_1434) begin
      btb_bank0_rd_data_way0_out_205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_206 <= 22'h0;
    end else if (_T_1438) begin
      btb_bank0_rd_data_way0_out_206 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_207 <= 22'h0;
    end else if (_T_1442) begin
      btb_bank0_rd_data_way0_out_207 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_208 <= 22'h0;
    end else if (_T_1446) begin
      btb_bank0_rd_data_way0_out_208 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_209 <= 22'h0;
    end else if (_T_1450) begin
      btb_bank0_rd_data_way0_out_209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_210 <= 22'h0;
    end else if (_T_1454) begin
      btb_bank0_rd_data_way0_out_210 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_211 <= 22'h0;
    end else if (_T_1458) begin
      btb_bank0_rd_data_way0_out_211 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_212 <= 22'h0;
    end else if (_T_1462) begin
      btb_bank0_rd_data_way0_out_212 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_213 <= 22'h0;
    end else if (_T_1466) begin
      btb_bank0_rd_data_way0_out_213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_214 <= 22'h0;
    end else if (_T_1470) begin
      btb_bank0_rd_data_way0_out_214 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_215 <= 22'h0;
    end else if (_T_1474) begin
      btb_bank0_rd_data_way0_out_215 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_216 <= 22'h0;
    end else if (_T_1478) begin
      btb_bank0_rd_data_way0_out_216 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_217 <= 22'h0;
    end else if (_T_1482) begin
      btb_bank0_rd_data_way0_out_217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_218 <= 22'h0;
    end else if (_T_1486) begin
      btb_bank0_rd_data_way0_out_218 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_219 <= 22'h0;
    end else if (_T_1490) begin
      btb_bank0_rd_data_way0_out_219 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_220 <= 22'h0;
    end else if (_T_1494) begin
      btb_bank0_rd_data_way0_out_220 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_221 <= 22'h0;
    end else if (_T_1498) begin
      btb_bank0_rd_data_way0_out_221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_222 <= 22'h0;
    end else if (_T_1502) begin
      btb_bank0_rd_data_way0_out_222 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_223 <= 22'h0;
    end else if (_T_1506) begin
      btb_bank0_rd_data_way0_out_223 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_224 <= 22'h0;
    end else if (_T_1510) begin
      btb_bank0_rd_data_way0_out_224 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_225 <= 22'h0;
    end else if (_T_1514) begin
      btb_bank0_rd_data_way0_out_225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_226 <= 22'h0;
    end else if (_T_1518) begin
      btb_bank0_rd_data_way0_out_226 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_227 <= 22'h0;
    end else if (_T_1522) begin
      btb_bank0_rd_data_way0_out_227 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_228 <= 22'h0;
    end else if (_T_1526) begin
      btb_bank0_rd_data_way0_out_228 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_229 <= 22'h0;
    end else if (_T_1530) begin
      btb_bank0_rd_data_way0_out_229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_230 <= 22'h0;
    end else if (_T_1534) begin
      btb_bank0_rd_data_way0_out_230 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_231 <= 22'h0;
    end else if (_T_1538) begin
      btb_bank0_rd_data_way0_out_231 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_232 <= 22'h0;
    end else if (_T_1542) begin
      btb_bank0_rd_data_way0_out_232 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_233 <= 22'h0;
    end else if (_T_1546) begin
      btb_bank0_rd_data_way0_out_233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_234 <= 22'h0;
    end else if (_T_1550) begin
      btb_bank0_rd_data_way0_out_234 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_235 <= 22'h0;
    end else if (_T_1554) begin
      btb_bank0_rd_data_way0_out_235 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_236 <= 22'h0;
    end else if (_T_1558) begin
      btb_bank0_rd_data_way0_out_236 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_237 <= 22'h0;
    end else if (_T_1562) begin
      btb_bank0_rd_data_way0_out_237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_238 <= 22'h0;
    end else if (_T_1566) begin
      btb_bank0_rd_data_way0_out_238 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_239 <= 22'h0;
    end else if (_T_1570) begin
      btb_bank0_rd_data_way0_out_239 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_240 <= 22'h0;
    end else if (_T_1574) begin
      btb_bank0_rd_data_way0_out_240 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_241 <= 22'h0;
    end else if (_T_1578) begin
      btb_bank0_rd_data_way0_out_241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_242 <= 22'h0;
    end else if (_T_1582) begin
      btb_bank0_rd_data_way0_out_242 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_243 <= 22'h0;
    end else if (_T_1586) begin
      btb_bank0_rd_data_way0_out_243 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_244 <= 22'h0;
    end else if (_T_1590) begin
      btb_bank0_rd_data_way0_out_244 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_245 <= 22'h0;
    end else if (_T_1594) begin
      btb_bank0_rd_data_way0_out_245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_246 <= 22'h0;
    end else if (_T_1598) begin
      btb_bank0_rd_data_way0_out_246 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_247 <= 22'h0;
    end else if (_T_1602) begin
      btb_bank0_rd_data_way0_out_247 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_248 <= 22'h0;
    end else if (_T_1606) begin
      btb_bank0_rd_data_way0_out_248 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_249 <= 22'h0;
    end else if (_T_1610) begin
      btb_bank0_rd_data_way0_out_249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_250 <= 22'h0;
    end else if (_T_1614) begin
      btb_bank0_rd_data_way0_out_250 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_251 <= 22'h0;
    end else if (_T_1618) begin
      btb_bank0_rd_data_way0_out_251 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_252 <= 22'h0;
    end else if (_T_1622) begin
      btb_bank0_rd_data_way0_out_252 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_253 <= 22'h0;
    end else if (_T_1626) begin
      btb_bank0_rd_data_way0_out_253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_254 <= 22'h0;
    end else if (_T_1630) begin
      btb_bank0_rd_data_way0_out_254 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way0_out_255 <= 22'h0;
    end else if (_T_1634) begin
      btb_bank0_rd_data_way0_out_255 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_0 <= 22'h0;
    end else if (_T_1638) begin
      btb_bank0_rd_data_way1_out_0 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_1 <= 22'h0;
    end else if (_T_1642) begin
      btb_bank0_rd_data_way1_out_1 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_2 <= 22'h0;
    end else if (_T_1646) begin
      btb_bank0_rd_data_way1_out_2 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_3 <= 22'h0;
    end else if (_T_1650) begin
      btb_bank0_rd_data_way1_out_3 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_4 <= 22'h0;
    end else if (_T_1654) begin
      btb_bank0_rd_data_way1_out_4 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_5 <= 22'h0;
    end else if (_T_1658) begin
      btb_bank0_rd_data_way1_out_5 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_6 <= 22'h0;
    end else if (_T_1662) begin
      btb_bank0_rd_data_way1_out_6 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_7 <= 22'h0;
    end else if (_T_1666) begin
      btb_bank0_rd_data_way1_out_7 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_8 <= 22'h0;
    end else if (_T_1670) begin
      btb_bank0_rd_data_way1_out_8 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_9 <= 22'h0;
    end else if (_T_1674) begin
      btb_bank0_rd_data_way1_out_9 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_10 <= 22'h0;
    end else if (_T_1678) begin
      btb_bank0_rd_data_way1_out_10 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_11 <= 22'h0;
    end else if (_T_1682) begin
      btb_bank0_rd_data_way1_out_11 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_12 <= 22'h0;
    end else if (_T_1686) begin
      btb_bank0_rd_data_way1_out_12 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_13 <= 22'h0;
    end else if (_T_1690) begin
      btb_bank0_rd_data_way1_out_13 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_14 <= 22'h0;
    end else if (_T_1694) begin
      btb_bank0_rd_data_way1_out_14 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_15 <= 22'h0;
    end else if (_T_1698) begin
      btb_bank0_rd_data_way1_out_15 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_16 <= 22'h0;
    end else if (_T_1702) begin
      btb_bank0_rd_data_way1_out_16 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_17 <= 22'h0;
    end else if (_T_1706) begin
      btb_bank0_rd_data_way1_out_17 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_18 <= 22'h0;
    end else if (_T_1710) begin
      btb_bank0_rd_data_way1_out_18 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_19 <= 22'h0;
    end else if (_T_1714) begin
      btb_bank0_rd_data_way1_out_19 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_20 <= 22'h0;
    end else if (_T_1718) begin
      btb_bank0_rd_data_way1_out_20 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_21 <= 22'h0;
    end else if (_T_1722) begin
      btb_bank0_rd_data_way1_out_21 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_22 <= 22'h0;
    end else if (_T_1726) begin
      btb_bank0_rd_data_way1_out_22 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_23 <= 22'h0;
    end else if (_T_1730) begin
      btb_bank0_rd_data_way1_out_23 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_24 <= 22'h0;
    end else if (_T_1734) begin
      btb_bank0_rd_data_way1_out_24 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_25 <= 22'h0;
    end else if (_T_1738) begin
      btb_bank0_rd_data_way1_out_25 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_26 <= 22'h0;
    end else if (_T_1742) begin
      btb_bank0_rd_data_way1_out_26 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_27 <= 22'h0;
    end else if (_T_1746) begin
      btb_bank0_rd_data_way1_out_27 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_28 <= 22'h0;
    end else if (_T_1750) begin
      btb_bank0_rd_data_way1_out_28 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_29 <= 22'h0;
    end else if (_T_1754) begin
      btb_bank0_rd_data_way1_out_29 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_30 <= 22'h0;
    end else if (_T_1758) begin
      btb_bank0_rd_data_way1_out_30 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_31 <= 22'h0;
    end else if (_T_1762) begin
      btb_bank0_rd_data_way1_out_31 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_32 <= 22'h0;
    end else if (_T_1766) begin
      btb_bank0_rd_data_way1_out_32 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_33 <= 22'h0;
    end else if (_T_1770) begin
      btb_bank0_rd_data_way1_out_33 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_34 <= 22'h0;
    end else if (_T_1774) begin
      btb_bank0_rd_data_way1_out_34 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_35 <= 22'h0;
    end else if (_T_1778) begin
      btb_bank0_rd_data_way1_out_35 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_36 <= 22'h0;
    end else if (_T_1782) begin
      btb_bank0_rd_data_way1_out_36 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_37 <= 22'h0;
    end else if (_T_1786) begin
      btb_bank0_rd_data_way1_out_37 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_38 <= 22'h0;
    end else if (_T_1790) begin
      btb_bank0_rd_data_way1_out_38 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_39 <= 22'h0;
    end else if (_T_1794) begin
      btb_bank0_rd_data_way1_out_39 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_40 <= 22'h0;
    end else if (_T_1798) begin
      btb_bank0_rd_data_way1_out_40 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_41 <= 22'h0;
    end else if (_T_1802) begin
      btb_bank0_rd_data_way1_out_41 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_42 <= 22'h0;
    end else if (_T_1806) begin
      btb_bank0_rd_data_way1_out_42 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_43 <= 22'h0;
    end else if (_T_1810) begin
      btb_bank0_rd_data_way1_out_43 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_44 <= 22'h0;
    end else if (_T_1814) begin
      btb_bank0_rd_data_way1_out_44 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_45 <= 22'h0;
    end else if (_T_1818) begin
      btb_bank0_rd_data_way1_out_45 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_46 <= 22'h0;
    end else if (_T_1822) begin
      btb_bank0_rd_data_way1_out_46 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_47 <= 22'h0;
    end else if (_T_1826) begin
      btb_bank0_rd_data_way1_out_47 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_48 <= 22'h0;
    end else if (_T_1830) begin
      btb_bank0_rd_data_way1_out_48 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_49 <= 22'h0;
    end else if (_T_1834) begin
      btb_bank0_rd_data_way1_out_49 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_50 <= 22'h0;
    end else if (_T_1838) begin
      btb_bank0_rd_data_way1_out_50 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_51 <= 22'h0;
    end else if (_T_1842) begin
      btb_bank0_rd_data_way1_out_51 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_52 <= 22'h0;
    end else if (_T_1846) begin
      btb_bank0_rd_data_way1_out_52 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_53 <= 22'h0;
    end else if (_T_1850) begin
      btb_bank0_rd_data_way1_out_53 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_54 <= 22'h0;
    end else if (_T_1854) begin
      btb_bank0_rd_data_way1_out_54 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_55 <= 22'h0;
    end else if (_T_1858) begin
      btb_bank0_rd_data_way1_out_55 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_56 <= 22'h0;
    end else if (_T_1862) begin
      btb_bank0_rd_data_way1_out_56 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_57 <= 22'h0;
    end else if (_T_1866) begin
      btb_bank0_rd_data_way1_out_57 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_58 <= 22'h0;
    end else if (_T_1870) begin
      btb_bank0_rd_data_way1_out_58 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_59 <= 22'h0;
    end else if (_T_1874) begin
      btb_bank0_rd_data_way1_out_59 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_60 <= 22'h0;
    end else if (_T_1878) begin
      btb_bank0_rd_data_way1_out_60 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_61 <= 22'h0;
    end else if (_T_1882) begin
      btb_bank0_rd_data_way1_out_61 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_62 <= 22'h0;
    end else if (_T_1886) begin
      btb_bank0_rd_data_way1_out_62 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_63 <= 22'h0;
    end else if (_T_1890) begin
      btb_bank0_rd_data_way1_out_63 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_64 <= 22'h0;
    end else if (_T_1894) begin
      btb_bank0_rd_data_way1_out_64 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_65 <= 22'h0;
    end else if (_T_1898) begin
      btb_bank0_rd_data_way1_out_65 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_66 <= 22'h0;
    end else if (_T_1902) begin
      btb_bank0_rd_data_way1_out_66 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_67 <= 22'h0;
    end else if (_T_1906) begin
      btb_bank0_rd_data_way1_out_67 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_68 <= 22'h0;
    end else if (_T_1910) begin
      btb_bank0_rd_data_way1_out_68 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_69 <= 22'h0;
    end else if (_T_1914) begin
      btb_bank0_rd_data_way1_out_69 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_70 <= 22'h0;
    end else if (_T_1918) begin
      btb_bank0_rd_data_way1_out_70 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_71 <= 22'h0;
    end else if (_T_1922) begin
      btb_bank0_rd_data_way1_out_71 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_72 <= 22'h0;
    end else if (_T_1926) begin
      btb_bank0_rd_data_way1_out_72 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_73 <= 22'h0;
    end else if (_T_1930) begin
      btb_bank0_rd_data_way1_out_73 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_74 <= 22'h0;
    end else if (_T_1934) begin
      btb_bank0_rd_data_way1_out_74 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_75 <= 22'h0;
    end else if (_T_1938) begin
      btb_bank0_rd_data_way1_out_75 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_76 <= 22'h0;
    end else if (_T_1942) begin
      btb_bank0_rd_data_way1_out_76 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_77 <= 22'h0;
    end else if (_T_1946) begin
      btb_bank0_rd_data_way1_out_77 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_78 <= 22'h0;
    end else if (_T_1950) begin
      btb_bank0_rd_data_way1_out_78 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_79 <= 22'h0;
    end else if (_T_1954) begin
      btb_bank0_rd_data_way1_out_79 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_80 <= 22'h0;
    end else if (_T_1958) begin
      btb_bank0_rd_data_way1_out_80 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_81 <= 22'h0;
    end else if (_T_1962) begin
      btb_bank0_rd_data_way1_out_81 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_82 <= 22'h0;
    end else if (_T_1966) begin
      btb_bank0_rd_data_way1_out_82 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_83 <= 22'h0;
    end else if (_T_1970) begin
      btb_bank0_rd_data_way1_out_83 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_84 <= 22'h0;
    end else if (_T_1974) begin
      btb_bank0_rd_data_way1_out_84 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_85 <= 22'h0;
    end else if (_T_1978) begin
      btb_bank0_rd_data_way1_out_85 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_86 <= 22'h0;
    end else if (_T_1982) begin
      btb_bank0_rd_data_way1_out_86 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_87 <= 22'h0;
    end else if (_T_1986) begin
      btb_bank0_rd_data_way1_out_87 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_88 <= 22'h0;
    end else if (_T_1990) begin
      btb_bank0_rd_data_way1_out_88 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_89 <= 22'h0;
    end else if (_T_1994) begin
      btb_bank0_rd_data_way1_out_89 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_90 <= 22'h0;
    end else if (_T_1998) begin
      btb_bank0_rd_data_way1_out_90 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_91 <= 22'h0;
    end else if (_T_2002) begin
      btb_bank0_rd_data_way1_out_91 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_92 <= 22'h0;
    end else if (_T_2006) begin
      btb_bank0_rd_data_way1_out_92 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_93 <= 22'h0;
    end else if (_T_2010) begin
      btb_bank0_rd_data_way1_out_93 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_94 <= 22'h0;
    end else if (_T_2014) begin
      btb_bank0_rd_data_way1_out_94 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_95 <= 22'h0;
    end else if (_T_2018) begin
      btb_bank0_rd_data_way1_out_95 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_96 <= 22'h0;
    end else if (_T_2022) begin
      btb_bank0_rd_data_way1_out_96 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_97 <= 22'h0;
    end else if (_T_2026) begin
      btb_bank0_rd_data_way1_out_97 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_98 <= 22'h0;
    end else if (_T_2030) begin
      btb_bank0_rd_data_way1_out_98 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_99 <= 22'h0;
    end else if (_T_2034) begin
      btb_bank0_rd_data_way1_out_99 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_100 <= 22'h0;
    end else if (_T_2038) begin
      btb_bank0_rd_data_way1_out_100 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_101 <= 22'h0;
    end else if (_T_2042) begin
      btb_bank0_rd_data_way1_out_101 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_102 <= 22'h0;
    end else if (_T_2046) begin
      btb_bank0_rd_data_way1_out_102 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_103 <= 22'h0;
    end else if (_T_2050) begin
      btb_bank0_rd_data_way1_out_103 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_104 <= 22'h0;
    end else if (_T_2054) begin
      btb_bank0_rd_data_way1_out_104 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_105 <= 22'h0;
    end else if (_T_2058) begin
      btb_bank0_rd_data_way1_out_105 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_106 <= 22'h0;
    end else if (_T_2062) begin
      btb_bank0_rd_data_way1_out_106 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_107 <= 22'h0;
    end else if (_T_2066) begin
      btb_bank0_rd_data_way1_out_107 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_108 <= 22'h0;
    end else if (_T_2070) begin
      btb_bank0_rd_data_way1_out_108 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_109 <= 22'h0;
    end else if (_T_2074) begin
      btb_bank0_rd_data_way1_out_109 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_110 <= 22'h0;
    end else if (_T_2078) begin
      btb_bank0_rd_data_way1_out_110 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_111 <= 22'h0;
    end else if (_T_2082) begin
      btb_bank0_rd_data_way1_out_111 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_112 <= 22'h0;
    end else if (_T_2086) begin
      btb_bank0_rd_data_way1_out_112 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_113 <= 22'h0;
    end else if (_T_2090) begin
      btb_bank0_rd_data_way1_out_113 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_114 <= 22'h0;
    end else if (_T_2094) begin
      btb_bank0_rd_data_way1_out_114 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_115 <= 22'h0;
    end else if (_T_2098) begin
      btb_bank0_rd_data_way1_out_115 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_116 <= 22'h0;
    end else if (_T_2102) begin
      btb_bank0_rd_data_way1_out_116 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_117 <= 22'h0;
    end else if (_T_2106) begin
      btb_bank0_rd_data_way1_out_117 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_118 <= 22'h0;
    end else if (_T_2110) begin
      btb_bank0_rd_data_way1_out_118 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_119 <= 22'h0;
    end else if (_T_2114) begin
      btb_bank0_rd_data_way1_out_119 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_120 <= 22'h0;
    end else if (_T_2118) begin
      btb_bank0_rd_data_way1_out_120 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_121 <= 22'h0;
    end else if (_T_2122) begin
      btb_bank0_rd_data_way1_out_121 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_122 <= 22'h0;
    end else if (_T_2126) begin
      btb_bank0_rd_data_way1_out_122 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_123 <= 22'h0;
    end else if (_T_2130) begin
      btb_bank0_rd_data_way1_out_123 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_124 <= 22'h0;
    end else if (_T_2134) begin
      btb_bank0_rd_data_way1_out_124 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_125 <= 22'h0;
    end else if (_T_2138) begin
      btb_bank0_rd_data_way1_out_125 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_126 <= 22'h0;
    end else if (_T_2142) begin
      btb_bank0_rd_data_way1_out_126 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_127 <= 22'h0;
    end else if (_T_2146) begin
      btb_bank0_rd_data_way1_out_127 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_128 <= 22'h0;
    end else if (_T_2150) begin
      btb_bank0_rd_data_way1_out_128 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_129 <= 22'h0;
    end else if (_T_2154) begin
      btb_bank0_rd_data_way1_out_129 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_130 <= 22'h0;
    end else if (_T_2158) begin
      btb_bank0_rd_data_way1_out_130 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_131 <= 22'h0;
    end else if (_T_2162) begin
      btb_bank0_rd_data_way1_out_131 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_132 <= 22'h0;
    end else if (_T_2166) begin
      btb_bank0_rd_data_way1_out_132 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_133 <= 22'h0;
    end else if (_T_2170) begin
      btb_bank0_rd_data_way1_out_133 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_134 <= 22'h0;
    end else if (_T_2174) begin
      btb_bank0_rd_data_way1_out_134 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_135 <= 22'h0;
    end else if (_T_2178) begin
      btb_bank0_rd_data_way1_out_135 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_136 <= 22'h0;
    end else if (_T_2182) begin
      btb_bank0_rd_data_way1_out_136 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_137 <= 22'h0;
    end else if (_T_2186) begin
      btb_bank0_rd_data_way1_out_137 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_138 <= 22'h0;
    end else if (_T_2190) begin
      btb_bank0_rd_data_way1_out_138 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_139 <= 22'h0;
    end else if (_T_2194) begin
      btb_bank0_rd_data_way1_out_139 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_140 <= 22'h0;
    end else if (_T_2198) begin
      btb_bank0_rd_data_way1_out_140 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_141 <= 22'h0;
    end else if (_T_2202) begin
      btb_bank0_rd_data_way1_out_141 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_142 <= 22'h0;
    end else if (_T_2206) begin
      btb_bank0_rd_data_way1_out_142 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_143 <= 22'h0;
    end else if (_T_2210) begin
      btb_bank0_rd_data_way1_out_143 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_144 <= 22'h0;
    end else if (_T_2214) begin
      btb_bank0_rd_data_way1_out_144 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_145 <= 22'h0;
    end else if (_T_2218) begin
      btb_bank0_rd_data_way1_out_145 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_146 <= 22'h0;
    end else if (_T_2222) begin
      btb_bank0_rd_data_way1_out_146 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_147 <= 22'h0;
    end else if (_T_2226) begin
      btb_bank0_rd_data_way1_out_147 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_148 <= 22'h0;
    end else if (_T_2230) begin
      btb_bank0_rd_data_way1_out_148 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_149 <= 22'h0;
    end else if (_T_2234) begin
      btb_bank0_rd_data_way1_out_149 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_150 <= 22'h0;
    end else if (_T_2238) begin
      btb_bank0_rd_data_way1_out_150 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_151 <= 22'h0;
    end else if (_T_2242) begin
      btb_bank0_rd_data_way1_out_151 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_152 <= 22'h0;
    end else if (_T_2246) begin
      btb_bank0_rd_data_way1_out_152 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_153 <= 22'h0;
    end else if (_T_2250) begin
      btb_bank0_rd_data_way1_out_153 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_154 <= 22'h0;
    end else if (_T_2254) begin
      btb_bank0_rd_data_way1_out_154 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_155 <= 22'h0;
    end else if (_T_2258) begin
      btb_bank0_rd_data_way1_out_155 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_156 <= 22'h0;
    end else if (_T_2262) begin
      btb_bank0_rd_data_way1_out_156 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_157 <= 22'h0;
    end else if (_T_2266) begin
      btb_bank0_rd_data_way1_out_157 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_158 <= 22'h0;
    end else if (_T_2270) begin
      btb_bank0_rd_data_way1_out_158 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_159 <= 22'h0;
    end else if (_T_2274) begin
      btb_bank0_rd_data_way1_out_159 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_160 <= 22'h0;
    end else if (_T_2278) begin
      btb_bank0_rd_data_way1_out_160 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_161 <= 22'h0;
    end else if (_T_2282) begin
      btb_bank0_rd_data_way1_out_161 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_162 <= 22'h0;
    end else if (_T_2286) begin
      btb_bank0_rd_data_way1_out_162 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_163 <= 22'h0;
    end else if (_T_2290) begin
      btb_bank0_rd_data_way1_out_163 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_164 <= 22'h0;
    end else if (_T_2294) begin
      btb_bank0_rd_data_way1_out_164 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_165 <= 22'h0;
    end else if (_T_2298) begin
      btb_bank0_rd_data_way1_out_165 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_166 <= 22'h0;
    end else if (_T_2302) begin
      btb_bank0_rd_data_way1_out_166 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_167 <= 22'h0;
    end else if (_T_2306) begin
      btb_bank0_rd_data_way1_out_167 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_168 <= 22'h0;
    end else if (_T_2310) begin
      btb_bank0_rd_data_way1_out_168 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_169 <= 22'h0;
    end else if (_T_2314) begin
      btb_bank0_rd_data_way1_out_169 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_170 <= 22'h0;
    end else if (_T_2318) begin
      btb_bank0_rd_data_way1_out_170 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_171 <= 22'h0;
    end else if (_T_2322) begin
      btb_bank0_rd_data_way1_out_171 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_172 <= 22'h0;
    end else if (_T_2326) begin
      btb_bank0_rd_data_way1_out_172 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_173 <= 22'h0;
    end else if (_T_2330) begin
      btb_bank0_rd_data_way1_out_173 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_174 <= 22'h0;
    end else if (_T_2334) begin
      btb_bank0_rd_data_way1_out_174 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_175 <= 22'h0;
    end else if (_T_2338) begin
      btb_bank0_rd_data_way1_out_175 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_176 <= 22'h0;
    end else if (_T_2342) begin
      btb_bank0_rd_data_way1_out_176 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_177 <= 22'h0;
    end else if (_T_2346) begin
      btb_bank0_rd_data_way1_out_177 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_178 <= 22'h0;
    end else if (_T_2350) begin
      btb_bank0_rd_data_way1_out_178 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_179 <= 22'h0;
    end else if (_T_2354) begin
      btb_bank0_rd_data_way1_out_179 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_180 <= 22'h0;
    end else if (_T_2358) begin
      btb_bank0_rd_data_way1_out_180 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_181 <= 22'h0;
    end else if (_T_2362) begin
      btb_bank0_rd_data_way1_out_181 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_182 <= 22'h0;
    end else if (_T_2366) begin
      btb_bank0_rd_data_way1_out_182 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_183 <= 22'h0;
    end else if (_T_2370) begin
      btb_bank0_rd_data_way1_out_183 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_184 <= 22'h0;
    end else if (_T_2374) begin
      btb_bank0_rd_data_way1_out_184 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_185 <= 22'h0;
    end else if (_T_2378) begin
      btb_bank0_rd_data_way1_out_185 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_186 <= 22'h0;
    end else if (_T_2382) begin
      btb_bank0_rd_data_way1_out_186 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_187 <= 22'h0;
    end else if (_T_2386) begin
      btb_bank0_rd_data_way1_out_187 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_188 <= 22'h0;
    end else if (_T_2390) begin
      btb_bank0_rd_data_way1_out_188 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_189 <= 22'h0;
    end else if (_T_2394) begin
      btb_bank0_rd_data_way1_out_189 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_190 <= 22'h0;
    end else if (_T_2398) begin
      btb_bank0_rd_data_way1_out_190 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_191 <= 22'h0;
    end else if (_T_2402) begin
      btb_bank0_rd_data_way1_out_191 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_192 <= 22'h0;
    end else if (_T_2406) begin
      btb_bank0_rd_data_way1_out_192 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_193 <= 22'h0;
    end else if (_T_2410) begin
      btb_bank0_rd_data_way1_out_193 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_194 <= 22'h0;
    end else if (_T_2414) begin
      btb_bank0_rd_data_way1_out_194 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_195 <= 22'h0;
    end else if (_T_2418) begin
      btb_bank0_rd_data_way1_out_195 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_196 <= 22'h0;
    end else if (_T_2422) begin
      btb_bank0_rd_data_way1_out_196 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_197 <= 22'h0;
    end else if (_T_2426) begin
      btb_bank0_rd_data_way1_out_197 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_198 <= 22'h0;
    end else if (_T_2430) begin
      btb_bank0_rd_data_way1_out_198 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_199 <= 22'h0;
    end else if (_T_2434) begin
      btb_bank0_rd_data_way1_out_199 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_200 <= 22'h0;
    end else if (_T_2438) begin
      btb_bank0_rd_data_way1_out_200 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_201 <= 22'h0;
    end else if (_T_2442) begin
      btb_bank0_rd_data_way1_out_201 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_202 <= 22'h0;
    end else if (_T_2446) begin
      btb_bank0_rd_data_way1_out_202 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_203 <= 22'h0;
    end else if (_T_2450) begin
      btb_bank0_rd_data_way1_out_203 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_204 <= 22'h0;
    end else if (_T_2454) begin
      btb_bank0_rd_data_way1_out_204 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_205 <= 22'h0;
    end else if (_T_2458) begin
      btb_bank0_rd_data_way1_out_205 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_206 <= 22'h0;
    end else if (_T_2462) begin
      btb_bank0_rd_data_way1_out_206 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_207 <= 22'h0;
    end else if (_T_2466) begin
      btb_bank0_rd_data_way1_out_207 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_208 <= 22'h0;
    end else if (_T_2470) begin
      btb_bank0_rd_data_way1_out_208 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_209 <= 22'h0;
    end else if (_T_2474) begin
      btb_bank0_rd_data_way1_out_209 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_210 <= 22'h0;
    end else if (_T_2478) begin
      btb_bank0_rd_data_way1_out_210 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_211 <= 22'h0;
    end else if (_T_2482) begin
      btb_bank0_rd_data_way1_out_211 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_212 <= 22'h0;
    end else if (_T_2486) begin
      btb_bank0_rd_data_way1_out_212 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_213 <= 22'h0;
    end else if (_T_2490) begin
      btb_bank0_rd_data_way1_out_213 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_214 <= 22'h0;
    end else if (_T_2494) begin
      btb_bank0_rd_data_way1_out_214 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_215 <= 22'h0;
    end else if (_T_2498) begin
      btb_bank0_rd_data_way1_out_215 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_216 <= 22'h0;
    end else if (_T_2502) begin
      btb_bank0_rd_data_way1_out_216 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_217 <= 22'h0;
    end else if (_T_2506) begin
      btb_bank0_rd_data_way1_out_217 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_218 <= 22'h0;
    end else if (_T_2510) begin
      btb_bank0_rd_data_way1_out_218 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_219 <= 22'h0;
    end else if (_T_2514) begin
      btb_bank0_rd_data_way1_out_219 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_220 <= 22'h0;
    end else if (_T_2518) begin
      btb_bank0_rd_data_way1_out_220 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_221 <= 22'h0;
    end else if (_T_2522) begin
      btb_bank0_rd_data_way1_out_221 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_222 <= 22'h0;
    end else if (_T_2526) begin
      btb_bank0_rd_data_way1_out_222 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_223 <= 22'h0;
    end else if (_T_2530) begin
      btb_bank0_rd_data_way1_out_223 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_224 <= 22'h0;
    end else if (_T_2534) begin
      btb_bank0_rd_data_way1_out_224 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_225 <= 22'h0;
    end else if (_T_2538) begin
      btb_bank0_rd_data_way1_out_225 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_226 <= 22'h0;
    end else if (_T_2542) begin
      btb_bank0_rd_data_way1_out_226 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_227 <= 22'h0;
    end else if (_T_2546) begin
      btb_bank0_rd_data_way1_out_227 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_228 <= 22'h0;
    end else if (_T_2550) begin
      btb_bank0_rd_data_way1_out_228 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_229 <= 22'h0;
    end else if (_T_2554) begin
      btb_bank0_rd_data_way1_out_229 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_230 <= 22'h0;
    end else if (_T_2558) begin
      btb_bank0_rd_data_way1_out_230 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_231 <= 22'h0;
    end else if (_T_2562) begin
      btb_bank0_rd_data_way1_out_231 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_232 <= 22'h0;
    end else if (_T_2566) begin
      btb_bank0_rd_data_way1_out_232 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_233 <= 22'h0;
    end else if (_T_2570) begin
      btb_bank0_rd_data_way1_out_233 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_234 <= 22'h0;
    end else if (_T_2574) begin
      btb_bank0_rd_data_way1_out_234 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_235 <= 22'h0;
    end else if (_T_2578) begin
      btb_bank0_rd_data_way1_out_235 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_236 <= 22'h0;
    end else if (_T_2582) begin
      btb_bank0_rd_data_way1_out_236 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_237 <= 22'h0;
    end else if (_T_2586) begin
      btb_bank0_rd_data_way1_out_237 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_238 <= 22'h0;
    end else if (_T_2590) begin
      btb_bank0_rd_data_way1_out_238 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_239 <= 22'h0;
    end else if (_T_2594) begin
      btb_bank0_rd_data_way1_out_239 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_240 <= 22'h0;
    end else if (_T_2598) begin
      btb_bank0_rd_data_way1_out_240 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_241 <= 22'h0;
    end else if (_T_2602) begin
      btb_bank0_rd_data_way1_out_241 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_242 <= 22'h0;
    end else if (_T_2606) begin
      btb_bank0_rd_data_way1_out_242 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_243 <= 22'h0;
    end else if (_T_2610) begin
      btb_bank0_rd_data_way1_out_243 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_244 <= 22'h0;
    end else if (_T_2614) begin
      btb_bank0_rd_data_way1_out_244 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_245 <= 22'h0;
    end else if (_T_2618) begin
      btb_bank0_rd_data_way1_out_245 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_246 <= 22'h0;
    end else if (_T_2622) begin
      btb_bank0_rd_data_way1_out_246 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_247 <= 22'h0;
    end else if (_T_2626) begin
      btb_bank0_rd_data_way1_out_247 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_248 <= 22'h0;
    end else if (_T_2630) begin
      btb_bank0_rd_data_way1_out_248 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_249 <= 22'h0;
    end else if (_T_2634) begin
      btb_bank0_rd_data_way1_out_249 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_250 <= 22'h0;
    end else if (_T_2638) begin
      btb_bank0_rd_data_way1_out_250 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_251 <= 22'h0;
    end else if (_T_2642) begin
      btb_bank0_rd_data_way1_out_251 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_252 <= 22'h0;
    end else if (_T_2646) begin
      btb_bank0_rd_data_way1_out_252 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_253 <= 22'h0;
    end else if (_T_2650) begin
      btb_bank0_rd_data_way1_out_253 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_254 <= 22'h0;
    end else if (_T_2654) begin
      btb_bank0_rd_data_way1_out_254 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_bank0_rd_data_way1_out_255 <= 22'h0;
    end else if (_T_2658) begin
      btb_bank0_rd_data_way1_out_255 <= btb_wr_data;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      fghr <= 8'h0;
    end else if (_T_349) begin
      fghr <= fghr_ns;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_0 <= 2'h0;
    end else if (bht_bank_sel_1_0_0) begin
      if (_T_9420) begin
        bht_bank_rd_data_out_1_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_1 <= 2'h0;
    end else if (bht_bank_sel_1_0_1) begin
      if (_T_9429) begin
        bht_bank_rd_data_out_1_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_2 <= 2'h0;
    end else if (bht_bank_sel_1_0_2) begin
      if (_T_9438) begin
        bht_bank_rd_data_out_1_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_3 <= 2'h0;
    end else if (bht_bank_sel_1_0_3) begin
      if (_T_9447) begin
        bht_bank_rd_data_out_1_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_4 <= 2'h0;
    end else if (bht_bank_sel_1_0_4) begin
      if (_T_9456) begin
        bht_bank_rd_data_out_1_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_5 <= 2'h0;
    end else if (bht_bank_sel_1_0_5) begin
      if (_T_9465) begin
        bht_bank_rd_data_out_1_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_6 <= 2'h0;
    end else if (bht_bank_sel_1_0_6) begin
      if (_T_9474) begin
        bht_bank_rd_data_out_1_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_7 <= 2'h0;
    end else if (bht_bank_sel_1_0_7) begin
      if (_T_9483) begin
        bht_bank_rd_data_out_1_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_8 <= 2'h0;
    end else if (bht_bank_sel_1_0_8) begin
      if (_T_9492) begin
        bht_bank_rd_data_out_1_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_9 <= 2'h0;
    end else if (bht_bank_sel_1_0_9) begin
      if (_T_9501) begin
        bht_bank_rd_data_out_1_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_10 <= 2'h0;
    end else if (bht_bank_sel_1_0_10) begin
      if (_T_9510) begin
        bht_bank_rd_data_out_1_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_11 <= 2'h0;
    end else if (bht_bank_sel_1_0_11) begin
      if (_T_9519) begin
        bht_bank_rd_data_out_1_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_12 <= 2'h0;
    end else if (bht_bank_sel_1_0_12) begin
      if (_T_9528) begin
        bht_bank_rd_data_out_1_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_13 <= 2'h0;
    end else if (bht_bank_sel_1_0_13) begin
      if (_T_9537) begin
        bht_bank_rd_data_out_1_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_14 <= 2'h0;
    end else if (bht_bank_sel_1_0_14) begin
      if (_T_9546) begin
        bht_bank_rd_data_out_1_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_15 <= 2'h0;
    end else if (bht_bank_sel_1_0_15) begin
      if (_T_9555) begin
        bht_bank_rd_data_out_1_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_16 <= 2'h0;
    end else if (bht_bank_sel_1_1_0) begin
      if (_T_9564) begin
        bht_bank_rd_data_out_1_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_17 <= 2'h0;
    end else if (bht_bank_sel_1_1_1) begin
      if (_T_9573) begin
        bht_bank_rd_data_out_1_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_18 <= 2'h0;
    end else if (bht_bank_sel_1_1_2) begin
      if (_T_9582) begin
        bht_bank_rd_data_out_1_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_19 <= 2'h0;
    end else if (bht_bank_sel_1_1_3) begin
      if (_T_9591) begin
        bht_bank_rd_data_out_1_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_20 <= 2'h0;
    end else if (bht_bank_sel_1_1_4) begin
      if (_T_9600) begin
        bht_bank_rd_data_out_1_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_21 <= 2'h0;
    end else if (bht_bank_sel_1_1_5) begin
      if (_T_9609) begin
        bht_bank_rd_data_out_1_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_22 <= 2'h0;
    end else if (bht_bank_sel_1_1_6) begin
      if (_T_9618) begin
        bht_bank_rd_data_out_1_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_23 <= 2'h0;
    end else if (bht_bank_sel_1_1_7) begin
      if (_T_9627) begin
        bht_bank_rd_data_out_1_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_24 <= 2'h0;
    end else if (bht_bank_sel_1_1_8) begin
      if (_T_9636) begin
        bht_bank_rd_data_out_1_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_25 <= 2'h0;
    end else if (bht_bank_sel_1_1_9) begin
      if (_T_9645) begin
        bht_bank_rd_data_out_1_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_26 <= 2'h0;
    end else if (bht_bank_sel_1_1_10) begin
      if (_T_9654) begin
        bht_bank_rd_data_out_1_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_27 <= 2'h0;
    end else if (bht_bank_sel_1_1_11) begin
      if (_T_9663) begin
        bht_bank_rd_data_out_1_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_28 <= 2'h0;
    end else if (bht_bank_sel_1_1_12) begin
      if (_T_9672) begin
        bht_bank_rd_data_out_1_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_29 <= 2'h0;
    end else if (bht_bank_sel_1_1_13) begin
      if (_T_9681) begin
        bht_bank_rd_data_out_1_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_30 <= 2'h0;
    end else if (bht_bank_sel_1_1_14) begin
      if (_T_9690) begin
        bht_bank_rd_data_out_1_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_31 <= 2'h0;
    end else if (bht_bank_sel_1_1_15) begin
      if (_T_9699) begin
        bht_bank_rd_data_out_1_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_32 <= 2'h0;
    end else if (bht_bank_sel_1_2_0) begin
      if (_T_9708) begin
        bht_bank_rd_data_out_1_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_33 <= 2'h0;
    end else if (bht_bank_sel_1_2_1) begin
      if (_T_9717) begin
        bht_bank_rd_data_out_1_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_34 <= 2'h0;
    end else if (bht_bank_sel_1_2_2) begin
      if (_T_9726) begin
        bht_bank_rd_data_out_1_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_35 <= 2'h0;
    end else if (bht_bank_sel_1_2_3) begin
      if (_T_9735) begin
        bht_bank_rd_data_out_1_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_36 <= 2'h0;
    end else if (bht_bank_sel_1_2_4) begin
      if (_T_9744) begin
        bht_bank_rd_data_out_1_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_37 <= 2'h0;
    end else if (bht_bank_sel_1_2_5) begin
      if (_T_9753) begin
        bht_bank_rd_data_out_1_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_38 <= 2'h0;
    end else if (bht_bank_sel_1_2_6) begin
      if (_T_9762) begin
        bht_bank_rd_data_out_1_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_39 <= 2'h0;
    end else if (bht_bank_sel_1_2_7) begin
      if (_T_9771) begin
        bht_bank_rd_data_out_1_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_40 <= 2'h0;
    end else if (bht_bank_sel_1_2_8) begin
      if (_T_9780) begin
        bht_bank_rd_data_out_1_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_41 <= 2'h0;
    end else if (bht_bank_sel_1_2_9) begin
      if (_T_9789) begin
        bht_bank_rd_data_out_1_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_42 <= 2'h0;
    end else if (bht_bank_sel_1_2_10) begin
      if (_T_9798) begin
        bht_bank_rd_data_out_1_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_43 <= 2'h0;
    end else if (bht_bank_sel_1_2_11) begin
      if (_T_9807) begin
        bht_bank_rd_data_out_1_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_44 <= 2'h0;
    end else if (bht_bank_sel_1_2_12) begin
      if (_T_9816) begin
        bht_bank_rd_data_out_1_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_45 <= 2'h0;
    end else if (bht_bank_sel_1_2_13) begin
      if (_T_9825) begin
        bht_bank_rd_data_out_1_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_46 <= 2'h0;
    end else if (bht_bank_sel_1_2_14) begin
      if (_T_9834) begin
        bht_bank_rd_data_out_1_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_47 <= 2'h0;
    end else if (bht_bank_sel_1_2_15) begin
      if (_T_9843) begin
        bht_bank_rd_data_out_1_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_48 <= 2'h0;
    end else if (bht_bank_sel_1_3_0) begin
      if (_T_9852) begin
        bht_bank_rd_data_out_1_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_49 <= 2'h0;
    end else if (bht_bank_sel_1_3_1) begin
      if (_T_9861) begin
        bht_bank_rd_data_out_1_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_50 <= 2'h0;
    end else if (bht_bank_sel_1_3_2) begin
      if (_T_9870) begin
        bht_bank_rd_data_out_1_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_51 <= 2'h0;
    end else if (bht_bank_sel_1_3_3) begin
      if (_T_9879) begin
        bht_bank_rd_data_out_1_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_52 <= 2'h0;
    end else if (bht_bank_sel_1_3_4) begin
      if (_T_9888) begin
        bht_bank_rd_data_out_1_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_53 <= 2'h0;
    end else if (bht_bank_sel_1_3_5) begin
      if (_T_9897) begin
        bht_bank_rd_data_out_1_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_54 <= 2'h0;
    end else if (bht_bank_sel_1_3_6) begin
      if (_T_9906) begin
        bht_bank_rd_data_out_1_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_55 <= 2'h0;
    end else if (bht_bank_sel_1_3_7) begin
      if (_T_9915) begin
        bht_bank_rd_data_out_1_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_56 <= 2'h0;
    end else if (bht_bank_sel_1_3_8) begin
      if (_T_9924) begin
        bht_bank_rd_data_out_1_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_57 <= 2'h0;
    end else if (bht_bank_sel_1_3_9) begin
      if (_T_9933) begin
        bht_bank_rd_data_out_1_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_58 <= 2'h0;
    end else if (bht_bank_sel_1_3_10) begin
      if (_T_9942) begin
        bht_bank_rd_data_out_1_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_59 <= 2'h0;
    end else if (bht_bank_sel_1_3_11) begin
      if (_T_9951) begin
        bht_bank_rd_data_out_1_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_60 <= 2'h0;
    end else if (bht_bank_sel_1_3_12) begin
      if (_T_9960) begin
        bht_bank_rd_data_out_1_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_61 <= 2'h0;
    end else if (bht_bank_sel_1_3_13) begin
      if (_T_9969) begin
        bht_bank_rd_data_out_1_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_62 <= 2'h0;
    end else if (bht_bank_sel_1_3_14) begin
      if (_T_9978) begin
        bht_bank_rd_data_out_1_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_63 <= 2'h0;
    end else if (bht_bank_sel_1_3_15) begin
      if (_T_9987) begin
        bht_bank_rd_data_out_1_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_64 <= 2'h0;
    end else if (bht_bank_sel_1_4_0) begin
      if (_T_9996) begin
        bht_bank_rd_data_out_1_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_65 <= 2'h0;
    end else if (bht_bank_sel_1_4_1) begin
      if (_T_10005) begin
        bht_bank_rd_data_out_1_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_66 <= 2'h0;
    end else if (bht_bank_sel_1_4_2) begin
      if (_T_10014) begin
        bht_bank_rd_data_out_1_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_67 <= 2'h0;
    end else if (bht_bank_sel_1_4_3) begin
      if (_T_10023) begin
        bht_bank_rd_data_out_1_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_68 <= 2'h0;
    end else if (bht_bank_sel_1_4_4) begin
      if (_T_10032) begin
        bht_bank_rd_data_out_1_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_69 <= 2'h0;
    end else if (bht_bank_sel_1_4_5) begin
      if (_T_10041) begin
        bht_bank_rd_data_out_1_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_70 <= 2'h0;
    end else if (bht_bank_sel_1_4_6) begin
      if (_T_10050) begin
        bht_bank_rd_data_out_1_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_71 <= 2'h0;
    end else if (bht_bank_sel_1_4_7) begin
      if (_T_10059) begin
        bht_bank_rd_data_out_1_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_72 <= 2'h0;
    end else if (bht_bank_sel_1_4_8) begin
      if (_T_10068) begin
        bht_bank_rd_data_out_1_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_73 <= 2'h0;
    end else if (bht_bank_sel_1_4_9) begin
      if (_T_10077) begin
        bht_bank_rd_data_out_1_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_74 <= 2'h0;
    end else if (bht_bank_sel_1_4_10) begin
      if (_T_10086) begin
        bht_bank_rd_data_out_1_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_75 <= 2'h0;
    end else if (bht_bank_sel_1_4_11) begin
      if (_T_10095) begin
        bht_bank_rd_data_out_1_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_76 <= 2'h0;
    end else if (bht_bank_sel_1_4_12) begin
      if (_T_10104) begin
        bht_bank_rd_data_out_1_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_77 <= 2'h0;
    end else if (bht_bank_sel_1_4_13) begin
      if (_T_10113) begin
        bht_bank_rd_data_out_1_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_78 <= 2'h0;
    end else if (bht_bank_sel_1_4_14) begin
      if (_T_10122) begin
        bht_bank_rd_data_out_1_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_79 <= 2'h0;
    end else if (bht_bank_sel_1_4_15) begin
      if (_T_10131) begin
        bht_bank_rd_data_out_1_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_80 <= 2'h0;
    end else if (bht_bank_sel_1_5_0) begin
      if (_T_10140) begin
        bht_bank_rd_data_out_1_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_81 <= 2'h0;
    end else if (bht_bank_sel_1_5_1) begin
      if (_T_10149) begin
        bht_bank_rd_data_out_1_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_82 <= 2'h0;
    end else if (bht_bank_sel_1_5_2) begin
      if (_T_10158) begin
        bht_bank_rd_data_out_1_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_83 <= 2'h0;
    end else if (bht_bank_sel_1_5_3) begin
      if (_T_10167) begin
        bht_bank_rd_data_out_1_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_84 <= 2'h0;
    end else if (bht_bank_sel_1_5_4) begin
      if (_T_10176) begin
        bht_bank_rd_data_out_1_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_85 <= 2'h0;
    end else if (bht_bank_sel_1_5_5) begin
      if (_T_10185) begin
        bht_bank_rd_data_out_1_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_86 <= 2'h0;
    end else if (bht_bank_sel_1_5_6) begin
      if (_T_10194) begin
        bht_bank_rd_data_out_1_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_87 <= 2'h0;
    end else if (bht_bank_sel_1_5_7) begin
      if (_T_10203) begin
        bht_bank_rd_data_out_1_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_88 <= 2'h0;
    end else if (bht_bank_sel_1_5_8) begin
      if (_T_10212) begin
        bht_bank_rd_data_out_1_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_89 <= 2'h0;
    end else if (bht_bank_sel_1_5_9) begin
      if (_T_10221) begin
        bht_bank_rd_data_out_1_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_90 <= 2'h0;
    end else if (bht_bank_sel_1_5_10) begin
      if (_T_10230) begin
        bht_bank_rd_data_out_1_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_91 <= 2'h0;
    end else if (bht_bank_sel_1_5_11) begin
      if (_T_10239) begin
        bht_bank_rd_data_out_1_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_92 <= 2'h0;
    end else if (bht_bank_sel_1_5_12) begin
      if (_T_10248) begin
        bht_bank_rd_data_out_1_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_93 <= 2'h0;
    end else if (bht_bank_sel_1_5_13) begin
      if (_T_10257) begin
        bht_bank_rd_data_out_1_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_94 <= 2'h0;
    end else if (bht_bank_sel_1_5_14) begin
      if (_T_10266) begin
        bht_bank_rd_data_out_1_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_95 <= 2'h0;
    end else if (bht_bank_sel_1_5_15) begin
      if (_T_10275) begin
        bht_bank_rd_data_out_1_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_96 <= 2'h0;
    end else if (bht_bank_sel_1_6_0) begin
      if (_T_10284) begin
        bht_bank_rd_data_out_1_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_97 <= 2'h0;
    end else if (bht_bank_sel_1_6_1) begin
      if (_T_10293) begin
        bht_bank_rd_data_out_1_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_98 <= 2'h0;
    end else if (bht_bank_sel_1_6_2) begin
      if (_T_10302) begin
        bht_bank_rd_data_out_1_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_99 <= 2'h0;
    end else if (bht_bank_sel_1_6_3) begin
      if (_T_10311) begin
        bht_bank_rd_data_out_1_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_100 <= 2'h0;
    end else if (bht_bank_sel_1_6_4) begin
      if (_T_10320) begin
        bht_bank_rd_data_out_1_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_101 <= 2'h0;
    end else if (bht_bank_sel_1_6_5) begin
      if (_T_10329) begin
        bht_bank_rd_data_out_1_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_102 <= 2'h0;
    end else if (bht_bank_sel_1_6_6) begin
      if (_T_10338) begin
        bht_bank_rd_data_out_1_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_103 <= 2'h0;
    end else if (bht_bank_sel_1_6_7) begin
      if (_T_10347) begin
        bht_bank_rd_data_out_1_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_104 <= 2'h0;
    end else if (bht_bank_sel_1_6_8) begin
      if (_T_10356) begin
        bht_bank_rd_data_out_1_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_105 <= 2'h0;
    end else if (bht_bank_sel_1_6_9) begin
      if (_T_10365) begin
        bht_bank_rd_data_out_1_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_106 <= 2'h0;
    end else if (bht_bank_sel_1_6_10) begin
      if (_T_10374) begin
        bht_bank_rd_data_out_1_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_107 <= 2'h0;
    end else if (bht_bank_sel_1_6_11) begin
      if (_T_10383) begin
        bht_bank_rd_data_out_1_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_108 <= 2'h0;
    end else if (bht_bank_sel_1_6_12) begin
      if (_T_10392) begin
        bht_bank_rd_data_out_1_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_109 <= 2'h0;
    end else if (bht_bank_sel_1_6_13) begin
      if (_T_10401) begin
        bht_bank_rd_data_out_1_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_110 <= 2'h0;
    end else if (bht_bank_sel_1_6_14) begin
      if (_T_10410) begin
        bht_bank_rd_data_out_1_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_111 <= 2'h0;
    end else if (bht_bank_sel_1_6_15) begin
      if (_T_10419) begin
        bht_bank_rd_data_out_1_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_112 <= 2'h0;
    end else if (bht_bank_sel_1_7_0) begin
      if (_T_10428) begin
        bht_bank_rd_data_out_1_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_113 <= 2'h0;
    end else if (bht_bank_sel_1_7_1) begin
      if (_T_10437) begin
        bht_bank_rd_data_out_1_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_114 <= 2'h0;
    end else if (bht_bank_sel_1_7_2) begin
      if (_T_10446) begin
        bht_bank_rd_data_out_1_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_115 <= 2'h0;
    end else if (bht_bank_sel_1_7_3) begin
      if (_T_10455) begin
        bht_bank_rd_data_out_1_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_116 <= 2'h0;
    end else if (bht_bank_sel_1_7_4) begin
      if (_T_10464) begin
        bht_bank_rd_data_out_1_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_117 <= 2'h0;
    end else if (bht_bank_sel_1_7_5) begin
      if (_T_10473) begin
        bht_bank_rd_data_out_1_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_118 <= 2'h0;
    end else if (bht_bank_sel_1_7_6) begin
      if (_T_10482) begin
        bht_bank_rd_data_out_1_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_119 <= 2'h0;
    end else if (bht_bank_sel_1_7_7) begin
      if (_T_10491) begin
        bht_bank_rd_data_out_1_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_120 <= 2'h0;
    end else if (bht_bank_sel_1_7_8) begin
      if (_T_10500) begin
        bht_bank_rd_data_out_1_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_121 <= 2'h0;
    end else if (bht_bank_sel_1_7_9) begin
      if (_T_10509) begin
        bht_bank_rd_data_out_1_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_122 <= 2'h0;
    end else if (bht_bank_sel_1_7_10) begin
      if (_T_10518) begin
        bht_bank_rd_data_out_1_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_123 <= 2'h0;
    end else if (bht_bank_sel_1_7_11) begin
      if (_T_10527) begin
        bht_bank_rd_data_out_1_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_124 <= 2'h0;
    end else if (bht_bank_sel_1_7_12) begin
      if (_T_10536) begin
        bht_bank_rd_data_out_1_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_125 <= 2'h0;
    end else if (bht_bank_sel_1_7_13) begin
      if (_T_10545) begin
        bht_bank_rd_data_out_1_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_126 <= 2'h0;
    end else if (bht_bank_sel_1_7_14) begin
      if (_T_10554) begin
        bht_bank_rd_data_out_1_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_127 <= 2'h0;
    end else if (bht_bank_sel_1_7_15) begin
      if (_T_10563) begin
        bht_bank_rd_data_out_1_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_128 <= 2'h0;
    end else if (bht_bank_sel_1_8_0) begin
      if (_T_10572) begin
        bht_bank_rd_data_out_1_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_129 <= 2'h0;
    end else if (bht_bank_sel_1_8_1) begin
      if (_T_10581) begin
        bht_bank_rd_data_out_1_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_130 <= 2'h0;
    end else if (bht_bank_sel_1_8_2) begin
      if (_T_10590) begin
        bht_bank_rd_data_out_1_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_131 <= 2'h0;
    end else if (bht_bank_sel_1_8_3) begin
      if (_T_10599) begin
        bht_bank_rd_data_out_1_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_132 <= 2'h0;
    end else if (bht_bank_sel_1_8_4) begin
      if (_T_10608) begin
        bht_bank_rd_data_out_1_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_133 <= 2'h0;
    end else if (bht_bank_sel_1_8_5) begin
      if (_T_10617) begin
        bht_bank_rd_data_out_1_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_134 <= 2'h0;
    end else if (bht_bank_sel_1_8_6) begin
      if (_T_10626) begin
        bht_bank_rd_data_out_1_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_135 <= 2'h0;
    end else if (bht_bank_sel_1_8_7) begin
      if (_T_10635) begin
        bht_bank_rd_data_out_1_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_136 <= 2'h0;
    end else if (bht_bank_sel_1_8_8) begin
      if (_T_10644) begin
        bht_bank_rd_data_out_1_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_137 <= 2'h0;
    end else if (bht_bank_sel_1_8_9) begin
      if (_T_10653) begin
        bht_bank_rd_data_out_1_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_138 <= 2'h0;
    end else if (bht_bank_sel_1_8_10) begin
      if (_T_10662) begin
        bht_bank_rd_data_out_1_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_139 <= 2'h0;
    end else if (bht_bank_sel_1_8_11) begin
      if (_T_10671) begin
        bht_bank_rd_data_out_1_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_140 <= 2'h0;
    end else if (bht_bank_sel_1_8_12) begin
      if (_T_10680) begin
        bht_bank_rd_data_out_1_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_141 <= 2'h0;
    end else if (bht_bank_sel_1_8_13) begin
      if (_T_10689) begin
        bht_bank_rd_data_out_1_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_142 <= 2'h0;
    end else if (bht_bank_sel_1_8_14) begin
      if (_T_10698) begin
        bht_bank_rd_data_out_1_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_143 <= 2'h0;
    end else if (bht_bank_sel_1_8_15) begin
      if (_T_10707) begin
        bht_bank_rd_data_out_1_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_144 <= 2'h0;
    end else if (bht_bank_sel_1_9_0) begin
      if (_T_10716) begin
        bht_bank_rd_data_out_1_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_145 <= 2'h0;
    end else if (bht_bank_sel_1_9_1) begin
      if (_T_10725) begin
        bht_bank_rd_data_out_1_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_146 <= 2'h0;
    end else if (bht_bank_sel_1_9_2) begin
      if (_T_10734) begin
        bht_bank_rd_data_out_1_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_147 <= 2'h0;
    end else if (bht_bank_sel_1_9_3) begin
      if (_T_10743) begin
        bht_bank_rd_data_out_1_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_148 <= 2'h0;
    end else if (bht_bank_sel_1_9_4) begin
      if (_T_10752) begin
        bht_bank_rd_data_out_1_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_149 <= 2'h0;
    end else if (bht_bank_sel_1_9_5) begin
      if (_T_10761) begin
        bht_bank_rd_data_out_1_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_150 <= 2'h0;
    end else if (bht_bank_sel_1_9_6) begin
      if (_T_10770) begin
        bht_bank_rd_data_out_1_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_151 <= 2'h0;
    end else if (bht_bank_sel_1_9_7) begin
      if (_T_10779) begin
        bht_bank_rd_data_out_1_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_152 <= 2'h0;
    end else if (bht_bank_sel_1_9_8) begin
      if (_T_10788) begin
        bht_bank_rd_data_out_1_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_153 <= 2'h0;
    end else if (bht_bank_sel_1_9_9) begin
      if (_T_10797) begin
        bht_bank_rd_data_out_1_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_154 <= 2'h0;
    end else if (bht_bank_sel_1_9_10) begin
      if (_T_10806) begin
        bht_bank_rd_data_out_1_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_155 <= 2'h0;
    end else if (bht_bank_sel_1_9_11) begin
      if (_T_10815) begin
        bht_bank_rd_data_out_1_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_156 <= 2'h0;
    end else if (bht_bank_sel_1_9_12) begin
      if (_T_10824) begin
        bht_bank_rd_data_out_1_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_157 <= 2'h0;
    end else if (bht_bank_sel_1_9_13) begin
      if (_T_10833) begin
        bht_bank_rd_data_out_1_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_158 <= 2'h0;
    end else if (bht_bank_sel_1_9_14) begin
      if (_T_10842) begin
        bht_bank_rd_data_out_1_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_159 <= 2'h0;
    end else if (bht_bank_sel_1_9_15) begin
      if (_T_10851) begin
        bht_bank_rd_data_out_1_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_160 <= 2'h0;
    end else if (bht_bank_sel_1_10_0) begin
      if (_T_10860) begin
        bht_bank_rd_data_out_1_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_161 <= 2'h0;
    end else if (bht_bank_sel_1_10_1) begin
      if (_T_10869) begin
        bht_bank_rd_data_out_1_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_162 <= 2'h0;
    end else if (bht_bank_sel_1_10_2) begin
      if (_T_10878) begin
        bht_bank_rd_data_out_1_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_163 <= 2'h0;
    end else if (bht_bank_sel_1_10_3) begin
      if (_T_10887) begin
        bht_bank_rd_data_out_1_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_164 <= 2'h0;
    end else if (bht_bank_sel_1_10_4) begin
      if (_T_10896) begin
        bht_bank_rd_data_out_1_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_165 <= 2'h0;
    end else if (bht_bank_sel_1_10_5) begin
      if (_T_10905) begin
        bht_bank_rd_data_out_1_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_166 <= 2'h0;
    end else if (bht_bank_sel_1_10_6) begin
      if (_T_10914) begin
        bht_bank_rd_data_out_1_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_167 <= 2'h0;
    end else if (bht_bank_sel_1_10_7) begin
      if (_T_10923) begin
        bht_bank_rd_data_out_1_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_168 <= 2'h0;
    end else if (bht_bank_sel_1_10_8) begin
      if (_T_10932) begin
        bht_bank_rd_data_out_1_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_169 <= 2'h0;
    end else if (bht_bank_sel_1_10_9) begin
      if (_T_10941) begin
        bht_bank_rd_data_out_1_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_170 <= 2'h0;
    end else if (bht_bank_sel_1_10_10) begin
      if (_T_10950) begin
        bht_bank_rd_data_out_1_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_171 <= 2'h0;
    end else if (bht_bank_sel_1_10_11) begin
      if (_T_10959) begin
        bht_bank_rd_data_out_1_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_172 <= 2'h0;
    end else if (bht_bank_sel_1_10_12) begin
      if (_T_10968) begin
        bht_bank_rd_data_out_1_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_173 <= 2'h0;
    end else if (bht_bank_sel_1_10_13) begin
      if (_T_10977) begin
        bht_bank_rd_data_out_1_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_174 <= 2'h0;
    end else if (bht_bank_sel_1_10_14) begin
      if (_T_10986) begin
        bht_bank_rd_data_out_1_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_175 <= 2'h0;
    end else if (bht_bank_sel_1_10_15) begin
      if (_T_10995) begin
        bht_bank_rd_data_out_1_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_176 <= 2'h0;
    end else if (bht_bank_sel_1_11_0) begin
      if (_T_11004) begin
        bht_bank_rd_data_out_1_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_177 <= 2'h0;
    end else if (bht_bank_sel_1_11_1) begin
      if (_T_11013) begin
        bht_bank_rd_data_out_1_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_178 <= 2'h0;
    end else if (bht_bank_sel_1_11_2) begin
      if (_T_11022) begin
        bht_bank_rd_data_out_1_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_179 <= 2'h0;
    end else if (bht_bank_sel_1_11_3) begin
      if (_T_11031) begin
        bht_bank_rd_data_out_1_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_180 <= 2'h0;
    end else if (bht_bank_sel_1_11_4) begin
      if (_T_11040) begin
        bht_bank_rd_data_out_1_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_181 <= 2'h0;
    end else if (bht_bank_sel_1_11_5) begin
      if (_T_11049) begin
        bht_bank_rd_data_out_1_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_182 <= 2'h0;
    end else if (bht_bank_sel_1_11_6) begin
      if (_T_11058) begin
        bht_bank_rd_data_out_1_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_183 <= 2'h0;
    end else if (bht_bank_sel_1_11_7) begin
      if (_T_11067) begin
        bht_bank_rd_data_out_1_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_184 <= 2'h0;
    end else if (bht_bank_sel_1_11_8) begin
      if (_T_11076) begin
        bht_bank_rd_data_out_1_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_185 <= 2'h0;
    end else if (bht_bank_sel_1_11_9) begin
      if (_T_11085) begin
        bht_bank_rd_data_out_1_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_186 <= 2'h0;
    end else if (bht_bank_sel_1_11_10) begin
      if (_T_11094) begin
        bht_bank_rd_data_out_1_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_187 <= 2'h0;
    end else if (bht_bank_sel_1_11_11) begin
      if (_T_11103) begin
        bht_bank_rd_data_out_1_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_188 <= 2'h0;
    end else if (bht_bank_sel_1_11_12) begin
      if (_T_11112) begin
        bht_bank_rd_data_out_1_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_189 <= 2'h0;
    end else if (bht_bank_sel_1_11_13) begin
      if (_T_11121) begin
        bht_bank_rd_data_out_1_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_190 <= 2'h0;
    end else if (bht_bank_sel_1_11_14) begin
      if (_T_11130) begin
        bht_bank_rd_data_out_1_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_191 <= 2'h0;
    end else if (bht_bank_sel_1_11_15) begin
      if (_T_11139) begin
        bht_bank_rd_data_out_1_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_192 <= 2'h0;
    end else if (bht_bank_sel_1_12_0) begin
      if (_T_11148) begin
        bht_bank_rd_data_out_1_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_193 <= 2'h0;
    end else if (bht_bank_sel_1_12_1) begin
      if (_T_11157) begin
        bht_bank_rd_data_out_1_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_194 <= 2'h0;
    end else if (bht_bank_sel_1_12_2) begin
      if (_T_11166) begin
        bht_bank_rd_data_out_1_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_195 <= 2'h0;
    end else if (bht_bank_sel_1_12_3) begin
      if (_T_11175) begin
        bht_bank_rd_data_out_1_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_196 <= 2'h0;
    end else if (bht_bank_sel_1_12_4) begin
      if (_T_11184) begin
        bht_bank_rd_data_out_1_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_197 <= 2'h0;
    end else if (bht_bank_sel_1_12_5) begin
      if (_T_11193) begin
        bht_bank_rd_data_out_1_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_198 <= 2'h0;
    end else if (bht_bank_sel_1_12_6) begin
      if (_T_11202) begin
        bht_bank_rd_data_out_1_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_199 <= 2'h0;
    end else if (bht_bank_sel_1_12_7) begin
      if (_T_11211) begin
        bht_bank_rd_data_out_1_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_200 <= 2'h0;
    end else if (bht_bank_sel_1_12_8) begin
      if (_T_11220) begin
        bht_bank_rd_data_out_1_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_201 <= 2'h0;
    end else if (bht_bank_sel_1_12_9) begin
      if (_T_11229) begin
        bht_bank_rd_data_out_1_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_202 <= 2'h0;
    end else if (bht_bank_sel_1_12_10) begin
      if (_T_11238) begin
        bht_bank_rd_data_out_1_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_203 <= 2'h0;
    end else if (bht_bank_sel_1_12_11) begin
      if (_T_11247) begin
        bht_bank_rd_data_out_1_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_204 <= 2'h0;
    end else if (bht_bank_sel_1_12_12) begin
      if (_T_11256) begin
        bht_bank_rd_data_out_1_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_205 <= 2'h0;
    end else if (bht_bank_sel_1_12_13) begin
      if (_T_11265) begin
        bht_bank_rd_data_out_1_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_206 <= 2'h0;
    end else if (bht_bank_sel_1_12_14) begin
      if (_T_11274) begin
        bht_bank_rd_data_out_1_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_207 <= 2'h0;
    end else if (bht_bank_sel_1_12_15) begin
      if (_T_11283) begin
        bht_bank_rd_data_out_1_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_208 <= 2'h0;
    end else if (bht_bank_sel_1_13_0) begin
      if (_T_11292) begin
        bht_bank_rd_data_out_1_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_209 <= 2'h0;
    end else if (bht_bank_sel_1_13_1) begin
      if (_T_11301) begin
        bht_bank_rd_data_out_1_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_210 <= 2'h0;
    end else if (bht_bank_sel_1_13_2) begin
      if (_T_11310) begin
        bht_bank_rd_data_out_1_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_211 <= 2'h0;
    end else if (bht_bank_sel_1_13_3) begin
      if (_T_11319) begin
        bht_bank_rd_data_out_1_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_212 <= 2'h0;
    end else if (bht_bank_sel_1_13_4) begin
      if (_T_11328) begin
        bht_bank_rd_data_out_1_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_213 <= 2'h0;
    end else if (bht_bank_sel_1_13_5) begin
      if (_T_11337) begin
        bht_bank_rd_data_out_1_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_214 <= 2'h0;
    end else if (bht_bank_sel_1_13_6) begin
      if (_T_11346) begin
        bht_bank_rd_data_out_1_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_215 <= 2'h0;
    end else if (bht_bank_sel_1_13_7) begin
      if (_T_11355) begin
        bht_bank_rd_data_out_1_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_216 <= 2'h0;
    end else if (bht_bank_sel_1_13_8) begin
      if (_T_11364) begin
        bht_bank_rd_data_out_1_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_217 <= 2'h0;
    end else if (bht_bank_sel_1_13_9) begin
      if (_T_11373) begin
        bht_bank_rd_data_out_1_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_218 <= 2'h0;
    end else if (bht_bank_sel_1_13_10) begin
      if (_T_11382) begin
        bht_bank_rd_data_out_1_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_219 <= 2'h0;
    end else if (bht_bank_sel_1_13_11) begin
      if (_T_11391) begin
        bht_bank_rd_data_out_1_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_220 <= 2'h0;
    end else if (bht_bank_sel_1_13_12) begin
      if (_T_11400) begin
        bht_bank_rd_data_out_1_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_221 <= 2'h0;
    end else if (bht_bank_sel_1_13_13) begin
      if (_T_11409) begin
        bht_bank_rd_data_out_1_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_222 <= 2'h0;
    end else if (bht_bank_sel_1_13_14) begin
      if (_T_11418) begin
        bht_bank_rd_data_out_1_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_223 <= 2'h0;
    end else if (bht_bank_sel_1_13_15) begin
      if (_T_11427) begin
        bht_bank_rd_data_out_1_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_224 <= 2'h0;
    end else if (bht_bank_sel_1_14_0) begin
      if (_T_11436) begin
        bht_bank_rd_data_out_1_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_225 <= 2'h0;
    end else if (bht_bank_sel_1_14_1) begin
      if (_T_11445) begin
        bht_bank_rd_data_out_1_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_226 <= 2'h0;
    end else if (bht_bank_sel_1_14_2) begin
      if (_T_11454) begin
        bht_bank_rd_data_out_1_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_227 <= 2'h0;
    end else if (bht_bank_sel_1_14_3) begin
      if (_T_11463) begin
        bht_bank_rd_data_out_1_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_228 <= 2'h0;
    end else if (bht_bank_sel_1_14_4) begin
      if (_T_11472) begin
        bht_bank_rd_data_out_1_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_229 <= 2'h0;
    end else if (bht_bank_sel_1_14_5) begin
      if (_T_11481) begin
        bht_bank_rd_data_out_1_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_230 <= 2'h0;
    end else if (bht_bank_sel_1_14_6) begin
      if (_T_11490) begin
        bht_bank_rd_data_out_1_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_231 <= 2'h0;
    end else if (bht_bank_sel_1_14_7) begin
      if (_T_11499) begin
        bht_bank_rd_data_out_1_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_232 <= 2'h0;
    end else if (bht_bank_sel_1_14_8) begin
      if (_T_11508) begin
        bht_bank_rd_data_out_1_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_233 <= 2'h0;
    end else if (bht_bank_sel_1_14_9) begin
      if (_T_11517) begin
        bht_bank_rd_data_out_1_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_234 <= 2'h0;
    end else if (bht_bank_sel_1_14_10) begin
      if (_T_11526) begin
        bht_bank_rd_data_out_1_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_235 <= 2'h0;
    end else if (bht_bank_sel_1_14_11) begin
      if (_T_11535) begin
        bht_bank_rd_data_out_1_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_236 <= 2'h0;
    end else if (bht_bank_sel_1_14_12) begin
      if (_T_11544) begin
        bht_bank_rd_data_out_1_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_237 <= 2'h0;
    end else if (bht_bank_sel_1_14_13) begin
      if (_T_11553) begin
        bht_bank_rd_data_out_1_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_238 <= 2'h0;
    end else if (bht_bank_sel_1_14_14) begin
      if (_T_11562) begin
        bht_bank_rd_data_out_1_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_239 <= 2'h0;
    end else if (bht_bank_sel_1_14_15) begin
      if (_T_11571) begin
        bht_bank_rd_data_out_1_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_240 <= 2'h0;
    end else if (bht_bank_sel_1_15_0) begin
      if (_T_11580) begin
        bht_bank_rd_data_out_1_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_241 <= 2'h0;
    end else if (bht_bank_sel_1_15_1) begin
      if (_T_11589) begin
        bht_bank_rd_data_out_1_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_242 <= 2'h0;
    end else if (bht_bank_sel_1_15_2) begin
      if (_T_11598) begin
        bht_bank_rd_data_out_1_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_243 <= 2'h0;
    end else if (bht_bank_sel_1_15_3) begin
      if (_T_11607) begin
        bht_bank_rd_data_out_1_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_244 <= 2'h0;
    end else if (bht_bank_sel_1_15_4) begin
      if (_T_11616) begin
        bht_bank_rd_data_out_1_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_245 <= 2'h0;
    end else if (bht_bank_sel_1_15_5) begin
      if (_T_11625) begin
        bht_bank_rd_data_out_1_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_246 <= 2'h0;
    end else if (bht_bank_sel_1_15_6) begin
      if (_T_11634) begin
        bht_bank_rd_data_out_1_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_247 <= 2'h0;
    end else if (bht_bank_sel_1_15_7) begin
      if (_T_11643) begin
        bht_bank_rd_data_out_1_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_248 <= 2'h0;
    end else if (bht_bank_sel_1_15_8) begin
      if (_T_11652) begin
        bht_bank_rd_data_out_1_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_249 <= 2'h0;
    end else if (bht_bank_sel_1_15_9) begin
      if (_T_11661) begin
        bht_bank_rd_data_out_1_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_250 <= 2'h0;
    end else if (bht_bank_sel_1_15_10) begin
      if (_T_11670) begin
        bht_bank_rd_data_out_1_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_251 <= 2'h0;
    end else if (bht_bank_sel_1_15_11) begin
      if (_T_11679) begin
        bht_bank_rd_data_out_1_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_252 <= 2'h0;
    end else if (bht_bank_sel_1_15_12) begin
      if (_T_11688) begin
        bht_bank_rd_data_out_1_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_253 <= 2'h0;
    end else if (bht_bank_sel_1_15_13) begin
      if (_T_11697) begin
        bht_bank_rd_data_out_1_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_254 <= 2'h0;
    end else if (bht_bank_sel_1_15_14) begin
      if (_T_11706) begin
        bht_bank_rd_data_out_1_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_1_255 <= 2'h0;
    end else if (bht_bank_sel_1_15_15) begin
      if (_T_11715) begin
        bht_bank_rd_data_out_1_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_1_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_0 <= 2'h0;
    end else if (bht_bank_sel_0_0_0) begin
      if (_T_7116) begin
        bht_bank_rd_data_out_0_0 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_0 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_1 <= 2'h0;
    end else if (bht_bank_sel_0_0_1) begin
      if (_T_7125) begin
        bht_bank_rd_data_out_0_1 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_1 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_2 <= 2'h0;
    end else if (bht_bank_sel_0_0_2) begin
      if (_T_7134) begin
        bht_bank_rd_data_out_0_2 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_2 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_3 <= 2'h0;
    end else if (bht_bank_sel_0_0_3) begin
      if (_T_7143) begin
        bht_bank_rd_data_out_0_3 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_3 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_4 <= 2'h0;
    end else if (bht_bank_sel_0_0_4) begin
      if (_T_7152) begin
        bht_bank_rd_data_out_0_4 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_4 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_5 <= 2'h0;
    end else if (bht_bank_sel_0_0_5) begin
      if (_T_7161) begin
        bht_bank_rd_data_out_0_5 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_5 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_6 <= 2'h0;
    end else if (bht_bank_sel_0_0_6) begin
      if (_T_7170) begin
        bht_bank_rd_data_out_0_6 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_6 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_7 <= 2'h0;
    end else if (bht_bank_sel_0_0_7) begin
      if (_T_7179) begin
        bht_bank_rd_data_out_0_7 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_7 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_8 <= 2'h0;
    end else if (bht_bank_sel_0_0_8) begin
      if (_T_7188) begin
        bht_bank_rd_data_out_0_8 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_8 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_9 <= 2'h0;
    end else if (bht_bank_sel_0_0_9) begin
      if (_T_7197) begin
        bht_bank_rd_data_out_0_9 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_9 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_10 <= 2'h0;
    end else if (bht_bank_sel_0_0_10) begin
      if (_T_7206) begin
        bht_bank_rd_data_out_0_10 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_10 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_11 <= 2'h0;
    end else if (bht_bank_sel_0_0_11) begin
      if (_T_7215) begin
        bht_bank_rd_data_out_0_11 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_11 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_12 <= 2'h0;
    end else if (bht_bank_sel_0_0_12) begin
      if (_T_7224) begin
        bht_bank_rd_data_out_0_12 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_12 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_13 <= 2'h0;
    end else if (bht_bank_sel_0_0_13) begin
      if (_T_7233) begin
        bht_bank_rd_data_out_0_13 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_13 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_14 <= 2'h0;
    end else if (bht_bank_sel_0_0_14) begin
      if (_T_7242) begin
        bht_bank_rd_data_out_0_14 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_14 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_15 <= 2'h0;
    end else if (bht_bank_sel_0_0_15) begin
      if (_T_7251) begin
        bht_bank_rd_data_out_0_15 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_15 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_16 <= 2'h0;
    end else if (bht_bank_sel_0_1_0) begin
      if (_T_7260) begin
        bht_bank_rd_data_out_0_16 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_16 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_17 <= 2'h0;
    end else if (bht_bank_sel_0_1_1) begin
      if (_T_7269) begin
        bht_bank_rd_data_out_0_17 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_17 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_18 <= 2'h0;
    end else if (bht_bank_sel_0_1_2) begin
      if (_T_7278) begin
        bht_bank_rd_data_out_0_18 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_18 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_19 <= 2'h0;
    end else if (bht_bank_sel_0_1_3) begin
      if (_T_7287) begin
        bht_bank_rd_data_out_0_19 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_19 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_20 <= 2'h0;
    end else if (bht_bank_sel_0_1_4) begin
      if (_T_7296) begin
        bht_bank_rd_data_out_0_20 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_20 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_21 <= 2'h0;
    end else if (bht_bank_sel_0_1_5) begin
      if (_T_7305) begin
        bht_bank_rd_data_out_0_21 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_21 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_22 <= 2'h0;
    end else if (bht_bank_sel_0_1_6) begin
      if (_T_7314) begin
        bht_bank_rd_data_out_0_22 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_22 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_23 <= 2'h0;
    end else if (bht_bank_sel_0_1_7) begin
      if (_T_7323) begin
        bht_bank_rd_data_out_0_23 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_23 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_24 <= 2'h0;
    end else if (bht_bank_sel_0_1_8) begin
      if (_T_7332) begin
        bht_bank_rd_data_out_0_24 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_24 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_25 <= 2'h0;
    end else if (bht_bank_sel_0_1_9) begin
      if (_T_7341) begin
        bht_bank_rd_data_out_0_25 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_25 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_26 <= 2'h0;
    end else if (bht_bank_sel_0_1_10) begin
      if (_T_7350) begin
        bht_bank_rd_data_out_0_26 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_26 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_27 <= 2'h0;
    end else if (bht_bank_sel_0_1_11) begin
      if (_T_7359) begin
        bht_bank_rd_data_out_0_27 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_27 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_28 <= 2'h0;
    end else if (bht_bank_sel_0_1_12) begin
      if (_T_7368) begin
        bht_bank_rd_data_out_0_28 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_28 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_29 <= 2'h0;
    end else if (bht_bank_sel_0_1_13) begin
      if (_T_7377) begin
        bht_bank_rd_data_out_0_29 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_29 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_30 <= 2'h0;
    end else if (bht_bank_sel_0_1_14) begin
      if (_T_7386) begin
        bht_bank_rd_data_out_0_30 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_30 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_31 <= 2'h0;
    end else if (bht_bank_sel_0_1_15) begin
      if (_T_7395) begin
        bht_bank_rd_data_out_0_31 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_31 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_32 <= 2'h0;
    end else if (bht_bank_sel_0_2_0) begin
      if (_T_7404) begin
        bht_bank_rd_data_out_0_32 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_32 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_33 <= 2'h0;
    end else if (bht_bank_sel_0_2_1) begin
      if (_T_7413) begin
        bht_bank_rd_data_out_0_33 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_33 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_34 <= 2'h0;
    end else if (bht_bank_sel_0_2_2) begin
      if (_T_7422) begin
        bht_bank_rd_data_out_0_34 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_34 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_35 <= 2'h0;
    end else if (bht_bank_sel_0_2_3) begin
      if (_T_7431) begin
        bht_bank_rd_data_out_0_35 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_35 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_36 <= 2'h0;
    end else if (bht_bank_sel_0_2_4) begin
      if (_T_7440) begin
        bht_bank_rd_data_out_0_36 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_36 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_37 <= 2'h0;
    end else if (bht_bank_sel_0_2_5) begin
      if (_T_7449) begin
        bht_bank_rd_data_out_0_37 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_37 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_38 <= 2'h0;
    end else if (bht_bank_sel_0_2_6) begin
      if (_T_7458) begin
        bht_bank_rd_data_out_0_38 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_38 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_39 <= 2'h0;
    end else if (bht_bank_sel_0_2_7) begin
      if (_T_7467) begin
        bht_bank_rd_data_out_0_39 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_39 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_40 <= 2'h0;
    end else if (bht_bank_sel_0_2_8) begin
      if (_T_7476) begin
        bht_bank_rd_data_out_0_40 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_40 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_41 <= 2'h0;
    end else if (bht_bank_sel_0_2_9) begin
      if (_T_7485) begin
        bht_bank_rd_data_out_0_41 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_41 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_42 <= 2'h0;
    end else if (bht_bank_sel_0_2_10) begin
      if (_T_7494) begin
        bht_bank_rd_data_out_0_42 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_42 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_43 <= 2'h0;
    end else if (bht_bank_sel_0_2_11) begin
      if (_T_7503) begin
        bht_bank_rd_data_out_0_43 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_43 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_44 <= 2'h0;
    end else if (bht_bank_sel_0_2_12) begin
      if (_T_7512) begin
        bht_bank_rd_data_out_0_44 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_44 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_45 <= 2'h0;
    end else if (bht_bank_sel_0_2_13) begin
      if (_T_7521) begin
        bht_bank_rd_data_out_0_45 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_45 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_46 <= 2'h0;
    end else if (bht_bank_sel_0_2_14) begin
      if (_T_7530) begin
        bht_bank_rd_data_out_0_46 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_46 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_47 <= 2'h0;
    end else if (bht_bank_sel_0_2_15) begin
      if (_T_7539) begin
        bht_bank_rd_data_out_0_47 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_47 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_48 <= 2'h0;
    end else if (bht_bank_sel_0_3_0) begin
      if (_T_7548) begin
        bht_bank_rd_data_out_0_48 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_48 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_49 <= 2'h0;
    end else if (bht_bank_sel_0_3_1) begin
      if (_T_7557) begin
        bht_bank_rd_data_out_0_49 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_49 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_50 <= 2'h0;
    end else if (bht_bank_sel_0_3_2) begin
      if (_T_7566) begin
        bht_bank_rd_data_out_0_50 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_50 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_51 <= 2'h0;
    end else if (bht_bank_sel_0_3_3) begin
      if (_T_7575) begin
        bht_bank_rd_data_out_0_51 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_51 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_52 <= 2'h0;
    end else if (bht_bank_sel_0_3_4) begin
      if (_T_7584) begin
        bht_bank_rd_data_out_0_52 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_52 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_53 <= 2'h0;
    end else if (bht_bank_sel_0_3_5) begin
      if (_T_7593) begin
        bht_bank_rd_data_out_0_53 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_53 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_54 <= 2'h0;
    end else if (bht_bank_sel_0_3_6) begin
      if (_T_7602) begin
        bht_bank_rd_data_out_0_54 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_54 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_55 <= 2'h0;
    end else if (bht_bank_sel_0_3_7) begin
      if (_T_7611) begin
        bht_bank_rd_data_out_0_55 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_55 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_56 <= 2'h0;
    end else if (bht_bank_sel_0_3_8) begin
      if (_T_7620) begin
        bht_bank_rd_data_out_0_56 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_56 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_57 <= 2'h0;
    end else if (bht_bank_sel_0_3_9) begin
      if (_T_7629) begin
        bht_bank_rd_data_out_0_57 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_57 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_58 <= 2'h0;
    end else if (bht_bank_sel_0_3_10) begin
      if (_T_7638) begin
        bht_bank_rd_data_out_0_58 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_58 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_59 <= 2'h0;
    end else if (bht_bank_sel_0_3_11) begin
      if (_T_7647) begin
        bht_bank_rd_data_out_0_59 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_59 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_60 <= 2'h0;
    end else if (bht_bank_sel_0_3_12) begin
      if (_T_7656) begin
        bht_bank_rd_data_out_0_60 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_60 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_61 <= 2'h0;
    end else if (bht_bank_sel_0_3_13) begin
      if (_T_7665) begin
        bht_bank_rd_data_out_0_61 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_61 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_62 <= 2'h0;
    end else if (bht_bank_sel_0_3_14) begin
      if (_T_7674) begin
        bht_bank_rd_data_out_0_62 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_62 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_63 <= 2'h0;
    end else if (bht_bank_sel_0_3_15) begin
      if (_T_7683) begin
        bht_bank_rd_data_out_0_63 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_63 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_64 <= 2'h0;
    end else if (bht_bank_sel_0_4_0) begin
      if (_T_7692) begin
        bht_bank_rd_data_out_0_64 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_64 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_65 <= 2'h0;
    end else if (bht_bank_sel_0_4_1) begin
      if (_T_7701) begin
        bht_bank_rd_data_out_0_65 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_65 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_66 <= 2'h0;
    end else if (bht_bank_sel_0_4_2) begin
      if (_T_7710) begin
        bht_bank_rd_data_out_0_66 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_66 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_67 <= 2'h0;
    end else if (bht_bank_sel_0_4_3) begin
      if (_T_7719) begin
        bht_bank_rd_data_out_0_67 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_67 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_68 <= 2'h0;
    end else if (bht_bank_sel_0_4_4) begin
      if (_T_7728) begin
        bht_bank_rd_data_out_0_68 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_68 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_69 <= 2'h0;
    end else if (bht_bank_sel_0_4_5) begin
      if (_T_7737) begin
        bht_bank_rd_data_out_0_69 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_69 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_70 <= 2'h0;
    end else if (bht_bank_sel_0_4_6) begin
      if (_T_7746) begin
        bht_bank_rd_data_out_0_70 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_70 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_71 <= 2'h0;
    end else if (bht_bank_sel_0_4_7) begin
      if (_T_7755) begin
        bht_bank_rd_data_out_0_71 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_71 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_72 <= 2'h0;
    end else if (bht_bank_sel_0_4_8) begin
      if (_T_7764) begin
        bht_bank_rd_data_out_0_72 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_72 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_73 <= 2'h0;
    end else if (bht_bank_sel_0_4_9) begin
      if (_T_7773) begin
        bht_bank_rd_data_out_0_73 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_73 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_74 <= 2'h0;
    end else if (bht_bank_sel_0_4_10) begin
      if (_T_7782) begin
        bht_bank_rd_data_out_0_74 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_74 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_75 <= 2'h0;
    end else if (bht_bank_sel_0_4_11) begin
      if (_T_7791) begin
        bht_bank_rd_data_out_0_75 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_75 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_76 <= 2'h0;
    end else if (bht_bank_sel_0_4_12) begin
      if (_T_7800) begin
        bht_bank_rd_data_out_0_76 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_76 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_77 <= 2'h0;
    end else if (bht_bank_sel_0_4_13) begin
      if (_T_7809) begin
        bht_bank_rd_data_out_0_77 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_77 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_78 <= 2'h0;
    end else if (bht_bank_sel_0_4_14) begin
      if (_T_7818) begin
        bht_bank_rd_data_out_0_78 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_78 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_79 <= 2'h0;
    end else if (bht_bank_sel_0_4_15) begin
      if (_T_7827) begin
        bht_bank_rd_data_out_0_79 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_79 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_80 <= 2'h0;
    end else if (bht_bank_sel_0_5_0) begin
      if (_T_7836) begin
        bht_bank_rd_data_out_0_80 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_80 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_81 <= 2'h0;
    end else if (bht_bank_sel_0_5_1) begin
      if (_T_7845) begin
        bht_bank_rd_data_out_0_81 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_81 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_82 <= 2'h0;
    end else if (bht_bank_sel_0_5_2) begin
      if (_T_7854) begin
        bht_bank_rd_data_out_0_82 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_82 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_83 <= 2'h0;
    end else if (bht_bank_sel_0_5_3) begin
      if (_T_7863) begin
        bht_bank_rd_data_out_0_83 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_83 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_84 <= 2'h0;
    end else if (bht_bank_sel_0_5_4) begin
      if (_T_7872) begin
        bht_bank_rd_data_out_0_84 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_84 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_85 <= 2'h0;
    end else if (bht_bank_sel_0_5_5) begin
      if (_T_7881) begin
        bht_bank_rd_data_out_0_85 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_85 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_86 <= 2'h0;
    end else if (bht_bank_sel_0_5_6) begin
      if (_T_7890) begin
        bht_bank_rd_data_out_0_86 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_86 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_87 <= 2'h0;
    end else if (bht_bank_sel_0_5_7) begin
      if (_T_7899) begin
        bht_bank_rd_data_out_0_87 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_87 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_88 <= 2'h0;
    end else if (bht_bank_sel_0_5_8) begin
      if (_T_7908) begin
        bht_bank_rd_data_out_0_88 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_88 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_89 <= 2'h0;
    end else if (bht_bank_sel_0_5_9) begin
      if (_T_7917) begin
        bht_bank_rd_data_out_0_89 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_89 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_90 <= 2'h0;
    end else if (bht_bank_sel_0_5_10) begin
      if (_T_7926) begin
        bht_bank_rd_data_out_0_90 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_90 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_91 <= 2'h0;
    end else if (bht_bank_sel_0_5_11) begin
      if (_T_7935) begin
        bht_bank_rd_data_out_0_91 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_91 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_92 <= 2'h0;
    end else if (bht_bank_sel_0_5_12) begin
      if (_T_7944) begin
        bht_bank_rd_data_out_0_92 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_92 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_93 <= 2'h0;
    end else if (bht_bank_sel_0_5_13) begin
      if (_T_7953) begin
        bht_bank_rd_data_out_0_93 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_93 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_94 <= 2'h0;
    end else if (bht_bank_sel_0_5_14) begin
      if (_T_7962) begin
        bht_bank_rd_data_out_0_94 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_94 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_95 <= 2'h0;
    end else if (bht_bank_sel_0_5_15) begin
      if (_T_7971) begin
        bht_bank_rd_data_out_0_95 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_95 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_96 <= 2'h0;
    end else if (bht_bank_sel_0_6_0) begin
      if (_T_7980) begin
        bht_bank_rd_data_out_0_96 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_96 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_97 <= 2'h0;
    end else if (bht_bank_sel_0_6_1) begin
      if (_T_7989) begin
        bht_bank_rd_data_out_0_97 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_97 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_98 <= 2'h0;
    end else if (bht_bank_sel_0_6_2) begin
      if (_T_7998) begin
        bht_bank_rd_data_out_0_98 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_98 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_99 <= 2'h0;
    end else if (bht_bank_sel_0_6_3) begin
      if (_T_8007) begin
        bht_bank_rd_data_out_0_99 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_99 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_100 <= 2'h0;
    end else if (bht_bank_sel_0_6_4) begin
      if (_T_8016) begin
        bht_bank_rd_data_out_0_100 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_100 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_101 <= 2'h0;
    end else if (bht_bank_sel_0_6_5) begin
      if (_T_8025) begin
        bht_bank_rd_data_out_0_101 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_101 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_102 <= 2'h0;
    end else if (bht_bank_sel_0_6_6) begin
      if (_T_8034) begin
        bht_bank_rd_data_out_0_102 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_102 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_103 <= 2'h0;
    end else if (bht_bank_sel_0_6_7) begin
      if (_T_8043) begin
        bht_bank_rd_data_out_0_103 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_103 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_104 <= 2'h0;
    end else if (bht_bank_sel_0_6_8) begin
      if (_T_8052) begin
        bht_bank_rd_data_out_0_104 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_104 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_105 <= 2'h0;
    end else if (bht_bank_sel_0_6_9) begin
      if (_T_8061) begin
        bht_bank_rd_data_out_0_105 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_105 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_106 <= 2'h0;
    end else if (bht_bank_sel_0_6_10) begin
      if (_T_8070) begin
        bht_bank_rd_data_out_0_106 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_106 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_107 <= 2'h0;
    end else if (bht_bank_sel_0_6_11) begin
      if (_T_8079) begin
        bht_bank_rd_data_out_0_107 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_107 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_108 <= 2'h0;
    end else if (bht_bank_sel_0_6_12) begin
      if (_T_8088) begin
        bht_bank_rd_data_out_0_108 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_108 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_109 <= 2'h0;
    end else if (bht_bank_sel_0_6_13) begin
      if (_T_8097) begin
        bht_bank_rd_data_out_0_109 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_109 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_110 <= 2'h0;
    end else if (bht_bank_sel_0_6_14) begin
      if (_T_8106) begin
        bht_bank_rd_data_out_0_110 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_110 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_111 <= 2'h0;
    end else if (bht_bank_sel_0_6_15) begin
      if (_T_8115) begin
        bht_bank_rd_data_out_0_111 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_111 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_112 <= 2'h0;
    end else if (bht_bank_sel_0_7_0) begin
      if (_T_8124) begin
        bht_bank_rd_data_out_0_112 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_112 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_113 <= 2'h0;
    end else if (bht_bank_sel_0_7_1) begin
      if (_T_8133) begin
        bht_bank_rd_data_out_0_113 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_113 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_114 <= 2'h0;
    end else if (bht_bank_sel_0_7_2) begin
      if (_T_8142) begin
        bht_bank_rd_data_out_0_114 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_114 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_115 <= 2'h0;
    end else if (bht_bank_sel_0_7_3) begin
      if (_T_8151) begin
        bht_bank_rd_data_out_0_115 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_115 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_116 <= 2'h0;
    end else if (bht_bank_sel_0_7_4) begin
      if (_T_8160) begin
        bht_bank_rd_data_out_0_116 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_116 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_117 <= 2'h0;
    end else if (bht_bank_sel_0_7_5) begin
      if (_T_8169) begin
        bht_bank_rd_data_out_0_117 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_117 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_118 <= 2'h0;
    end else if (bht_bank_sel_0_7_6) begin
      if (_T_8178) begin
        bht_bank_rd_data_out_0_118 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_118 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_119 <= 2'h0;
    end else if (bht_bank_sel_0_7_7) begin
      if (_T_8187) begin
        bht_bank_rd_data_out_0_119 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_119 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_120 <= 2'h0;
    end else if (bht_bank_sel_0_7_8) begin
      if (_T_8196) begin
        bht_bank_rd_data_out_0_120 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_120 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_121 <= 2'h0;
    end else if (bht_bank_sel_0_7_9) begin
      if (_T_8205) begin
        bht_bank_rd_data_out_0_121 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_121 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_122 <= 2'h0;
    end else if (bht_bank_sel_0_7_10) begin
      if (_T_8214) begin
        bht_bank_rd_data_out_0_122 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_122 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_123 <= 2'h0;
    end else if (bht_bank_sel_0_7_11) begin
      if (_T_8223) begin
        bht_bank_rd_data_out_0_123 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_123 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_124 <= 2'h0;
    end else if (bht_bank_sel_0_7_12) begin
      if (_T_8232) begin
        bht_bank_rd_data_out_0_124 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_124 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_125 <= 2'h0;
    end else if (bht_bank_sel_0_7_13) begin
      if (_T_8241) begin
        bht_bank_rd_data_out_0_125 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_125 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_126 <= 2'h0;
    end else if (bht_bank_sel_0_7_14) begin
      if (_T_8250) begin
        bht_bank_rd_data_out_0_126 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_126 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_127 <= 2'h0;
    end else if (bht_bank_sel_0_7_15) begin
      if (_T_8259) begin
        bht_bank_rd_data_out_0_127 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_127 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_128 <= 2'h0;
    end else if (bht_bank_sel_0_8_0) begin
      if (_T_8268) begin
        bht_bank_rd_data_out_0_128 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_128 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_129 <= 2'h0;
    end else if (bht_bank_sel_0_8_1) begin
      if (_T_8277) begin
        bht_bank_rd_data_out_0_129 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_129 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_130 <= 2'h0;
    end else if (bht_bank_sel_0_8_2) begin
      if (_T_8286) begin
        bht_bank_rd_data_out_0_130 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_130 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_131 <= 2'h0;
    end else if (bht_bank_sel_0_8_3) begin
      if (_T_8295) begin
        bht_bank_rd_data_out_0_131 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_131 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_132 <= 2'h0;
    end else if (bht_bank_sel_0_8_4) begin
      if (_T_8304) begin
        bht_bank_rd_data_out_0_132 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_132 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_133 <= 2'h0;
    end else if (bht_bank_sel_0_8_5) begin
      if (_T_8313) begin
        bht_bank_rd_data_out_0_133 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_133 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_134 <= 2'h0;
    end else if (bht_bank_sel_0_8_6) begin
      if (_T_8322) begin
        bht_bank_rd_data_out_0_134 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_134 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_135 <= 2'h0;
    end else if (bht_bank_sel_0_8_7) begin
      if (_T_8331) begin
        bht_bank_rd_data_out_0_135 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_135 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_136 <= 2'h0;
    end else if (bht_bank_sel_0_8_8) begin
      if (_T_8340) begin
        bht_bank_rd_data_out_0_136 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_136 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_137 <= 2'h0;
    end else if (bht_bank_sel_0_8_9) begin
      if (_T_8349) begin
        bht_bank_rd_data_out_0_137 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_137 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_138 <= 2'h0;
    end else if (bht_bank_sel_0_8_10) begin
      if (_T_8358) begin
        bht_bank_rd_data_out_0_138 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_138 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_139 <= 2'h0;
    end else if (bht_bank_sel_0_8_11) begin
      if (_T_8367) begin
        bht_bank_rd_data_out_0_139 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_139 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_140 <= 2'h0;
    end else if (bht_bank_sel_0_8_12) begin
      if (_T_8376) begin
        bht_bank_rd_data_out_0_140 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_140 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_141 <= 2'h0;
    end else if (bht_bank_sel_0_8_13) begin
      if (_T_8385) begin
        bht_bank_rd_data_out_0_141 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_141 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_142 <= 2'h0;
    end else if (bht_bank_sel_0_8_14) begin
      if (_T_8394) begin
        bht_bank_rd_data_out_0_142 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_142 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_143 <= 2'h0;
    end else if (bht_bank_sel_0_8_15) begin
      if (_T_8403) begin
        bht_bank_rd_data_out_0_143 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_143 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_144 <= 2'h0;
    end else if (bht_bank_sel_0_9_0) begin
      if (_T_8412) begin
        bht_bank_rd_data_out_0_144 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_144 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_145 <= 2'h0;
    end else if (bht_bank_sel_0_9_1) begin
      if (_T_8421) begin
        bht_bank_rd_data_out_0_145 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_145 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_146 <= 2'h0;
    end else if (bht_bank_sel_0_9_2) begin
      if (_T_8430) begin
        bht_bank_rd_data_out_0_146 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_146 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_147 <= 2'h0;
    end else if (bht_bank_sel_0_9_3) begin
      if (_T_8439) begin
        bht_bank_rd_data_out_0_147 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_147 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_148 <= 2'h0;
    end else if (bht_bank_sel_0_9_4) begin
      if (_T_8448) begin
        bht_bank_rd_data_out_0_148 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_148 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_149 <= 2'h0;
    end else if (bht_bank_sel_0_9_5) begin
      if (_T_8457) begin
        bht_bank_rd_data_out_0_149 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_149 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_150 <= 2'h0;
    end else if (bht_bank_sel_0_9_6) begin
      if (_T_8466) begin
        bht_bank_rd_data_out_0_150 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_150 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_151 <= 2'h0;
    end else if (bht_bank_sel_0_9_7) begin
      if (_T_8475) begin
        bht_bank_rd_data_out_0_151 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_151 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_152 <= 2'h0;
    end else if (bht_bank_sel_0_9_8) begin
      if (_T_8484) begin
        bht_bank_rd_data_out_0_152 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_152 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_153 <= 2'h0;
    end else if (bht_bank_sel_0_9_9) begin
      if (_T_8493) begin
        bht_bank_rd_data_out_0_153 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_153 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_154 <= 2'h0;
    end else if (bht_bank_sel_0_9_10) begin
      if (_T_8502) begin
        bht_bank_rd_data_out_0_154 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_154 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_155 <= 2'h0;
    end else if (bht_bank_sel_0_9_11) begin
      if (_T_8511) begin
        bht_bank_rd_data_out_0_155 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_155 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_156 <= 2'h0;
    end else if (bht_bank_sel_0_9_12) begin
      if (_T_8520) begin
        bht_bank_rd_data_out_0_156 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_156 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_157 <= 2'h0;
    end else if (bht_bank_sel_0_9_13) begin
      if (_T_8529) begin
        bht_bank_rd_data_out_0_157 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_157 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_158 <= 2'h0;
    end else if (bht_bank_sel_0_9_14) begin
      if (_T_8538) begin
        bht_bank_rd_data_out_0_158 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_158 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_159 <= 2'h0;
    end else if (bht_bank_sel_0_9_15) begin
      if (_T_8547) begin
        bht_bank_rd_data_out_0_159 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_159 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_160 <= 2'h0;
    end else if (bht_bank_sel_0_10_0) begin
      if (_T_8556) begin
        bht_bank_rd_data_out_0_160 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_160 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_161 <= 2'h0;
    end else if (bht_bank_sel_0_10_1) begin
      if (_T_8565) begin
        bht_bank_rd_data_out_0_161 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_161 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_162 <= 2'h0;
    end else if (bht_bank_sel_0_10_2) begin
      if (_T_8574) begin
        bht_bank_rd_data_out_0_162 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_162 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_163 <= 2'h0;
    end else if (bht_bank_sel_0_10_3) begin
      if (_T_8583) begin
        bht_bank_rd_data_out_0_163 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_163 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_164 <= 2'h0;
    end else if (bht_bank_sel_0_10_4) begin
      if (_T_8592) begin
        bht_bank_rd_data_out_0_164 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_164 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_165 <= 2'h0;
    end else if (bht_bank_sel_0_10_5) begin
      if (_T_8601) begin
        bht_bank_rd_data_out_0_165 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_165 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_166 <= 2'h0;
    end else if (bht_bank_sel_0_10_6) begin
      if (_T_8610) begin
        bht_bank_rd_data_out_0_166 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_166 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_167 <= 2'h0;
    end else if (bht_bank_sel_0_10_7) begin
      if (_T_8619) begin
        bht_bank_rd_data_out_0_167 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_167 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_168 <= 2'h0;
    end else if (bht_bank_sel_0_10_8) begin
      if (_T_8628) begin
        bht_bank_rd_data_out_0_168 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_168 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_169 <= 2'h0;
    end else if (bht_bank_sel_0_10_9) begin
      if (_T_8637) begin
        bht_bank_rd_data_out_0_169 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_169 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_170 <= 2'h0;
    end else if (bht_bank_sel_0_10_10) begin
      if (_T_8646) begin
        bht_bank_rd_data_out_0_170 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_170 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_171 <= 2'h0;
    end else if (bht_bank_sel_0_10_11) begin
      if (_T_8655) begin
        bht_bank_rd_data_out_0_171 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_171 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_172 <= 2'h0;
    end else if (bht_bank_sel_0_10_12) begin
      if (_T_8664) begin
        bht_bank_rd_data_out_0_172 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_172 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_173 <= 2'h0;
    end else if (bht_bank_sel_0_10_13) begin
      if (_T_8673) begin
        bht_bank_rd_data_out_0_173 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_173 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_174 <= 2'h0;
    end else if (bht_bank_sel_0_10_14) begin
      if (_T_8682) begin
        bht_bank_rd_data_out_0_174 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_174 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_175 <= 2'h0;
    end else if (bht_bank_sel_0_10_15) begin
      if (_T_8691) begin
        bht_bank_rd_data_out_0_175 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_175 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_176 <= 2'h0;
    end else if (bht_bank_sel_0_11_0) begin
      if (_T_8700) begin
        bht_bank_rd_data_out_0_176 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_176 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_177 <= 2'h0;
    end else if (bht_bank_sel_0_11_1) begin
      if (_T_8709) begin
        bht_bank_rd_data_out_0_177 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_177 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_178 <= 2'h0;
    end else if (bht_bank_sel_0_11_2) begin
      if (_T_8718) begin
        bht_bank_rd_data_out_0_178 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_178 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_179 <= 2'h0;
    end else if (bht_bank_sel_0_11_3) begin
      if (_T_8727) begin
        bht_bank_rd_data_out_0_179 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_179 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_180 <= 2'h0;
    end else if (bht_bank_sel_0_11_4) begin
      if (_T_8736) begin
        bht_bank_rd_data_out_0_180 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_180 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_181 <= 2'h0;
    end else if (bht_bank_sel_0_11_5) begin
      if (_T_8745) begin
        bht_bank_rd_data_out_0_181 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_181 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_182 <= 2'h0;
    end else if (bht_bank_sel_0_11_6) begin
      if (_T_8754) begin
        bht_bank_rd_data_out_0_182 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_182 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_183 <= 2'h0;
    end else if (bht_bank_sel_0_11_7) begin
      if (_T_8763) begin
        bht_bank_rd_data_out_0_183 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_183 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_184 <= 2'h0;
    end else if (bht_bank_sel_0_11_8) begin
      if (_T_8772) begin
        bht_bank_rd_data_out_0_184 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_184 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_185 <= 2'h0;
    end else if (bht_bank_sel_0_11_9) begin
      if (_T_8781) begin
        bht_bank_rd_data_out_0_185 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_185 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_186 <= 2'h0;
    end else if (bht_bank_sel_0_11_10) begin
      if (_T_8790) begin
        bht_bank_rd_data_out_0_186 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_186 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_187 <= 2'h0;
    end else if (bht_bank_sel_0_11_11) begin
      if (_T_8799) begin
        bht_bank_rd_data_out_0_187 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_187 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_188 <= 2'h0;
    end else if (bht_bank_sel_0_11_12) begin
      if (_T_8808) begin
        bht_bank_rd_data_out_0_188 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_188 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_189 <= 2'h0;
    end else if (bht_bank_sel_0_11_13) begin
      if (_T_8817) begin
        bht_bank_rd_data_out_0_189 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_189 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_190 <= 2'h0;
    end else if (bht_bank_sel_0_11_14) begin
      if (_T_8826) begin
        bht_bank_rd_data_out_0_190 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_190 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_191 <= 2'h0;
    end else if (bht_bank_sel_0_11_15) begin
      if (_T_8835) begin
        bht_bank_rd_data_out_0_191 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_191 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_192 <= 2'h0;
    end else if (bht_bank_sel_0_12_0) begin
      if (_T_8844) begin
        bht_bank_rd_data_out_0_192 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_192 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_193 <= 2'h0;
    end else if (bht_bank_sel_0_12_1) begin
      if (_T_8853) begin
        bht_bank_rd_data_out_0_193 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_193 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_194 <= 2'h0;
    end else if (bht_bank_sel_0_12_2) begin
      if (_T_8862) begin
        bht_bank_rd_data_out_0_194 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_194 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_195 <= 2'h0;
    end else if (bht_bank_sel_0_12_3) begin
      if (_T_8871) begin
        bht_bank_rd_data_out_0_195 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_195 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_196 <= 2'h0;
    end else if (bht_bank_sel_0_12_4) begin
      if (_T_8880) begin
        bht_bank_rd_data_out_0_196 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_196 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_197 <= 2'h0;
    end else if (bht_bank_sel_0_12_5) begin
      if (_T_8889) begin
        bht_bank_rd_data_out_0_197 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_197 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_198 <= 2'h0;
    end else if (bht_bank_sel_0_12_6) begin
      if (_T_8898) begin
        bht_bank_rd_data_out_0_198 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_198 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_199 <= 2'h0;
    end else if (bht_bank_sel_0_12_7) begin
      if (_T_8907) begin
        bht_bank_rd_data_out_0_199 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_199 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_200 <= 2'h0;
    end else if (bht_bank_sel_0_12_8) begin
      if (_T_8916) begin
        bht_bank_rd_data_out_0_200 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_200 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_201 <= 2'h0;
    end else if (bht_bank_sel_0_12_9) begin
      if (_T_8925) begin
        bht_bank_rd_data_out_0_201 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_201 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_202 <= 2'h0;
    end else if (bht_bank_sel_0_12_10) begin
      if (_T_8934) begin
        bht_bank_rd_data_out_0_202 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_202 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_203 <= 2'h0;
    end else if (bht_bank_sel_0_12_11) begin
      if (_T_8943) begin
        bht_bank_rd_data_out_0_203 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_203 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_204 <= 2'h0;
    end else if (bht_bank_sel_0_12_12) begin
      if (_T_8952) begin
        bht_bank_rd_data_out_0_204 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_204 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_205 <= 2'h0;
    end else if (bht_bank_sel_0_12_13) begin
      if (_T_8961) begin
        bht_bank_rd_data_out_0_205 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_205 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_206 <= 2'h0;
    end else if (bht_bank_sel_0_12_14) begin
      if (_T_8970) begin
        bht_bank_rd_data_out_0_206 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_206 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_207 <= 2'h0;
    end else if (bht_bank_sel_0_12_15) begin
      if (_T_8979) begin
        bht_bank_rd_data_out_0_207 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_207 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_208 <= 2'h0;
    end else if (bht_bank_sel_0_13_0) begin
      if (_T_8988) begin
        bht_bank_rd_data_out_0_208 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_208 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_209 <= 2'h0;
    end else if (bht_bank_sel_0_13_1) begin
      if (_T_8997) begin
        bht_bank_rd_data_out_0_209 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_209 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_210 <= 2'h0;
    end else if (bht_bank_sel_0_13_2) begin
      if (_T_9006) begin
        bht_bank_rd_data_out_0_210 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_210 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_211 <= 2'h0;
    end else if (bht_bank_sel_0_13_3) begin
      if (_T_9015) begin
        bht_bank_rd_data_out_0_211 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_211 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_212 <= 2'h0;
    end else if (bht_bank_sel_0_13_4) begin
      if (_T_9024) begin
        bht_bank_rd_data_out_0_212 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_212 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_213 <= 2'h0;
    end else if (bht_bank_sel_0_13_5) begin
      if (_T_9033) begin
        bht_bank_rd_data_out_0_213 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_213 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_214 <= 2'h0;
    end else if (bht_bank_sel_0_13_6) begin
      if (_T_9042) begin
        bht_bank_rd_data_out_0_214 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_214 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_215 <= 2'h0;
    end else if (bht_bank_sel_0_13_7) begin
      if (_T_9051) begin
        bht_bank_rd_data_out_0_215 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_215 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_216 <= 2'h0;
    end else if (bht_bank_sel_0_13_8) begin
      if (_T_9060) begin
        bht_bank_rd_data_out_0_216 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_216 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_217 <= 2'h0;
    end else if (bht_bank_sel_0_13_9) begin
      if (_T_9069) begin
        bht_bank_rd_data_out_0_217 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_217 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_218 <= 2'h0;
    end else if (bht_bank_sel_0_13_10) begin
      if (_T_9078) begin
        bht_bank_rd_data_out_0_218 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_218 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_219 <= 2'h0;
    end else if (bht_bank_sel_0_13_11) begin
      if (_T_9087) begin
        bht_bank_rd_data_out_0_219 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_219 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_220 <= 2'h0;
    end else if (bht_bank_sel_0_13_12) begin
      if (_T_9096) begin
        bht_bank_rd_data_out_0_220 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_220 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_221 <= 2'h0;
    end else if (bht_bank_sel_0_13_13) begin
      if (_T_9105) begin
        bht_bank_rd_data_out_0_221 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_221 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_222 <= 2'h0;
    end else if (bht_bank_sel_0_13_14) begin
      if (_T_9114) begin
        bht_bank_rd_data_out_0_222 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_222 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_223 <= 2'h0;
    end else if (bht_bank_sel_0_13_15) begin
      if (_T_9123) begin
        bht_bank_rd_data_out_0_223 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_223 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_224 <= 2'h0;
    end else if (bht_bank_sel_0_14_0) begin
      if (_T_9132) begin
        bht_bank_rd_data_out_0_224 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_224 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_225 <= 2'h0;
    end else if (bht_bank_sel_0_14_1) begin
      if (_T_9141) begin
        bht_bank_rd_data_out_0_225 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_225 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_226 <= 2'h0;
    end else if (bht_bank_sel_0_14_2) begin
      if (_T_9150) begin
        bht_bank_rd_data_out_0_226 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_226 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_227 <= 2'h0;
    end else if (bht_bank_sel_0_14_3) begin
      if (_T_9159) begin
        bht_bank_rd_data_out_0_227 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_227 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_228 <= 2'h0;
    end else if (bht_bank_sel_0_14_4) begin
      if (_T_9168) begin
        bht_bank_rd_data_out_0_228 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_228 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_229 <= 2'h0;
    end else if (bht_bank_sel_0_14_5) begin
      if (_T_9177) begin
        bht_bank_rd_data_out_0_229 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_229 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_230 <= 2'h0;
    end else if (bht_bank_sel_0_14_6) begin
      if (_T_9186) begin
        bht_bank_rd_data_out_0_230 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_230 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_231 <= 2'h0;
    end else if (bht_bank_sel_0_14_7) begin
      if (_T_9195) begin
        bht_bank_rd_data_out_0_231 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_231 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_232 <= 2'h0;
    end else if (bht_bank_sel_0_14_8) begin
      if (_T_9204) begin
        bht_bank_rd_data_out_0_232 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_232 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_233 <= 2'h0;
    end else if (bht_bank_sel_0_14_9) begin
      if (_T_9213) begin
        bht_bank_rd_data_out_0_233 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_233 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_234 <= 2'h0;
    end else if (bht_bank_sel_0_14_10) begin
      if (_T_9222) begin
        bht_bank_rd_data_out_0_234 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_234 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_235 <= 2'h0;
    end else if (bht_bank_sel_0_14_11) begin
      if (_T_9231) begin
        bht_bank_rd_data_out_0_235 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_235 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_236 <= 2'h0;
    end else if (bht_bank_sel_0_14_12) begin
      if (_T_9240) begin
        bht_bank_rd_data_out_0_236 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_236 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_237 <= 2'h0;
    end else if (bht_bank_sel_0_14_13) begin
      if (_T_9249) begin
        bht_bank_rd_data_out_0_237 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_237 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_238 <= 2'h0;
    end else if (bht_bank_sel_0_14_14) begin
      if (_T_9258) begin
        bht_bank_rd_data_out_0_238 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_238 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_239 <= 2'h0;
    end else if (bht_bank_sel_0_14_15) begin
      if (_T_9267) begin
        bht_bank_rd_data_out_0_239 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_239 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_240 <= 2'h0;
    end else if (bht_bank_sel_0_15_0) begin
      if (_T_9276) begin
        bht_bank_rd_data_out_0_240 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_240 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_241 <= 2'h0;
    end else if (bht_bank_sel_0_15_1) begin
      if (_T_9285) begin
        bht_bank_rd_data_out_0_241 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_241 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_242 <= 2'h0;
    end else if (bht_bank_sel_0_15_2) begin
      if (_T_9294) begin
        bht_bank_rd_data_out_0_242 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_242 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_243 <= 2'h0;
    end else if (bht_bank_sel_0_15_3) begin
      if (_T_9303) begin
        bht_bank_rd_data_out_0_243 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_243 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_244 <= 2'h0;
    end else if (bht_bank_sel_0_15_4) begin
      if (_T_9312) begin
        bht_bank_rd_data_out_0_244 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_244 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_245 <= 2'h0;
    end else if (bht_bank_sel_0_15_5) begin
      if (_T_9321) begin
        bht_bank_rd_data_out_0_245 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_245 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_246 <= 2'h0;
    end else if (bht_bank_sel_0_15_6) begin
      if (_T_9330) begin
        bht_bank_rd_data_out_0_246 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_246 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_247 <= 2'h0;
    end else if (bht_bank_sel_0_15_7) begin
      if (_T_9339) begin
        bht_bank_rd_data_out_0_247 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_247 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_248 <= 2'h0;
    end else if (bht_bank_sel_0_15_8) begin
      if (_T_9348) begin
        bht_bank_rd_data_out_0_248 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_248 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_249 <= 2'h0;
    end else if (bht_bank_sel_0_15_9) begin
      if (_T_9357) begin
        bht_bank_rd_data_out_0_249 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_249 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_250 <= 2'h0;
    end else if (bht_bank_sel_0_15_10) begin
      if (_T_9366) begin
        bht_bank_rd_data_out_0_250 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_250 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_251 <= 2'h0;
    end else if (bht_bank_sel_0_15_11) begin
      if (_T_9375) begin
        bht_bank_rd_data_out_0_251 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_251 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_252 <= 2'h0;
    end else if (bht_bank_sel_0_15_12) begin
      if (_T_9384) begin
        bht_bank_rd_data_out_0_252 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_252 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_253 <= 2'h0;
    end else if (bht_bank_sel_0_15_13) begin
      if (_T_9393) begin
        bht_bank_rd_data_out_0_253 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_253 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_254 <= 2'h0;
    end else if (bht_bank_sel_0_15_14) begin
      if (_T_9402) begin
        bht_bank_rd_data_out_0_254 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_254 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      bht_bank_rd_data_out_0_255 <= 2'h0;
    end else if (bht_bank_sel_0_15_15) begin
      if (_T_9411) begin
        bht_bank_rd_data_out_0_255 <= io_dec_bp_dec_tlu_br0_r_pkt_bits_hist;
      end else begin
        bht_bank_rd_data_out_0_255 <= io_exu_bp_exu_mp_pkt_bits_hist;
      end
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      exu_mp_way_f <= 1'h0;
    end else if (_T_341) begin
      exu_mp_way_f <= io_exu_bp_exu_mp_pkt_bits_way;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      btb_lru_b0_f <= 256'h0;
    end else if (_T_208) begin
      btb_lru_b0_f <= btb_lru_b0_ns;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      exu_flush_final_d1 <= 1'h0;
    end else if (_T_345) begin
      exu_flush_final_d1 <= io_exu_flush_final;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      ifc_fetch_adder_prior <= 30'h0;
    end else if (_T_385) begin
      ifc_fetch_adder_prior <= io_ifc_fetch_addr_f[30:1];
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_0 <= 32'h0;
    end else if (rsenable_0) begin
      rets_out_0 <= rets_in_0;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_1 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_1 <= rets_in_1;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_2 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_2 <= rets_in_2;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_3 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_3 <= rets_in_3;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_4 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_4 <= rets_in_4;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_5 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_5 <= rets_in_5;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_6 <= 32'h0;
    end else if (rsenable_1) begin
      rets_out_6 <= rets_in_6;
    end
  end
  always @(posedge clock or posedge reset) begin
    if (reset) begin
      rets_out_7 <= 32'h0;
    end else if (rs_push) begin
      rets_out_7 <= rets_out_6;
    end
  end
endmodule
