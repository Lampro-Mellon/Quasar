module el2_dec_trigger(
  input         clock,
  input         reset,
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input         io_trigger_pkt_any_0_execute,
  input         io_trigger_pkt_any_0_m,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input         io_trigger_pkt_any_1_execute,
  input         io_trigger_pkt_any_1_m,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input         io_trigger_pkt_any_2_execute,
  input         io_trigger_pkt_any_2_m,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input         io_trigger_pkt_any_3_execute,
  input         io_trigger_pkt_any_3_m,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input  [30:0] io_dec_i0_pc_d,
  output [3:0]  io_dec_i0_trigger_match_d
);
  wire  _T = ~io_trigger_pkt_any_0_select; // @[el2_lsu_trigger.scala 15:63]
  wire  _T_1 = _T & io_trigger_pkt_any_0_execute; // @[el2_lsu_trigger.scala 15:93]
  wire [9:0] _T_11 = {_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [18:0] _T_20 = {_T_11,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [27:0] _T_29 = {_T_20,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_33 = {_T_29,_T_1,_T_1,_T_1,_T_1}; // @[Cat.scala 29:58]
  wire [31:0] _T_35 = {io_dec_i0_pc_d,io_trigger_pkt_any_0_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_0 = _T_33 & _T_35; // @[el2_lsu_trigger.scala 15:127]
  wire  _T_37 = ~io_trigger_pkt_any_1_select; // @[el2_lsu_trigger.scala 15:63]
  wire  _T_38 = _T_37 & io_trigger_pkt_any_1_execute; // @[el2_lsu_trigger.scala 15:93]
  wire [9:0] _T_48 = {_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [18:0] _T_57 = {_T_48,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [27:0] _T_66 = {_T_57,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [31:0] _T_70 = {_T_66,_T_38,_T_38,_T_38,_T_38}; // @[Cat.scala 29:58]
  wire [31:0] _T_72 = {io_dec_i0_pc_d,io_trigger_pkt_any_1_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_1 = _T_70 & _T_72; // @[el2_lsu_trigger.scala 15:127]
  wire  _T_74 = ~io_trigger_pkt_any_2_select; // @[el2_lsu_trigger.scala 15:63]
  wire  _T_75 = _T_74 & io_trigger_pkt_any_2_execute; // @[el2_lsu_trigger.scala 15:93]
  wire [9:0] _T_85 = {_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [18:0] _T_94 = {_T_85,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [27:0] _T_103 = {_T_94,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [31:0] _T_107 = {_T_103,_T_75,_T_75,_T_75,_T_75}; // @[Cat.scala 29:58]
  wire [31:0] _T_109 = {io_dec_i0_pc_d,io_trigger_pkt_any_2_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_2 = _T_107 & _T_109; // @[el2_lsu_trigger.scala 15:127]
  wire  _T_111 = ~io_trigger_pkt_any_3_select; // @[el2_lsu_trigger.scala 15:63]
  wire  _T_112 = _T_111 & io_trigger_pkt_any_3_execute; // @[el2_lsu_trigger.scala 15:93]
  wire [9:0] _T_122 = {_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [18:0] _T_131 = {_T_122,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [27:0] _T_140 = {_T_131,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [31:0] _T_144 = {_T_140,_T_112,_T_112,_T_112,_T_112}; // @[Cat.scala 29:58]
  wire [31:0] _T_146 = {io_dec_i0_pc_d,io_trigger_pkt_any_3_tdata2[0]}; // @[Cat.scala 29:58]
  wire [31:0] dec_i0_match_data_3 = _T_144 & _T_146; // @[el2_lsu_trigger.scala 15:127]
  wire  _T_148 = io_trigger_pkt_any_0_execute & io_trigger_pkt_any_0_m; // @[el2_lsu_trigger.scala 16:83]
  wire  _T_151 = &io_trigger_pkt_any_0_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_152 = ~_T_151; // @[el2_lib.scala 194:39]
  wire  _T_153 = io_trigger_pkt_any_0_match_ & _T_152; // @[el2_lib.scala 194:37]
  wire  _T_156 = io_trigger_pkt_any_0_tdata2[0] == dec_i0_match_data_0[0]; // @[el2_lib.scala 195:52]
  wire  _T_157 = _T_153 | _T_156; // @[el2_lib.scala 195:41]
  wire  _T_159 = &io_trigger_pkt_any_0_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_160 = _T_159 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_163 = io_trigger_pkt_any_0_tdata2[1] == dec_i0_match_data_0[1]; // @[el2_lib.scala 197:80]
  wire  _T_164 = _T_160 | _T_163; // @[el2_lib.scala 197:25]
  wire  _T_166 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_167 = _T_166 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_170 = io_trigger_pkt_any_0_tdata2[2] == dec_i0_match_data_0[2]; // @[el2_lib.scala 197:80]
  wire  _T_171 = _T_167 | _T_170; // @[el2_lib.scala 197:25]
  wire  _T_173 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_174 = _T_173 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_177 = io_trigger_pkt_any_0_tdata2[3] == dec_i0_match_data_0[3]; // @[el2_lib.scala 197:80]
  wire  _T_178 = _T_174 | _T_177; // @[el2_lib.scala 197:25]
  wire  _T_180 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_181 = _T_180 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_184 = io_trigger_pkt_any_0_tdata2[4] == dec_i0_match_data_0[4]; // @[el2_lib.scala 197:80]
  wire  _T_185 = _T_181 | _T_184; // @[el2_lib.scala 197:25]
  wire  _T_187 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_188 = _T_187 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_191 = io_trigger_pkt_any_0_tdata2[5] == dec_i0_match_data_0[5]; // @[el2_lib.scala 197:80]
  wire  _T_192 = _T_188 | _T_191; // @[el2_lib.scala 197:25]
  wire  _T_194 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_195 = _T_194 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_198 = io_trigger_pkt_any_0_tdata2[6] == dec_i0_match_data_0[6]; // @[el2_lib.scala 197:80]
  wire  _T_199 = _T_195 | _T_198; // @[el2_lib.scala 197:25]
  wire  _T_201 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_202 = _T_201 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_205 = io_trigger_pkt_any_0_tdata2[7] == dec_i0_match_data_0[7]; // @[el2_lib.scala 197:80]
  wire  _T_206 = _T_202 | _T_205; // @[el2_lib.scala 197:25]
  wire  _T_208 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_209 = _T_208 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_212 = io_trigger_pkt_any_0_tdata2[8] == dec_i0_match_data_0[8]; // @[el2_lib.scala 197:80]
  wire  _T_213 = _T_209 | _T_212; // @[el2_lib.scala 197:25]
  wire  _T_215 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_216 = _T_215 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_219 = io_trigger_pkt_any_0_tdata2[9] == dec_i0_match_data_0[9]; // @[el2_lib.scala 197:80]
  wire  _T_220 = _T_216 | _T_219; // @[el2_lib.scala 197:25]
  wire  _T_222 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_223 = _T_222 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_226 = io_trigger_pkt_any_0_tdata2[10] == dec_i0_match_data_0[10]; // @[el2_lib.scala 197:80]
  wire  _T_227 = _T_223 | _T_226; // @[el2_lib.scala 197:25]
  wire  _T_229 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_230 = _T_229 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_233 = io_trigger_pkt_any_0_tdata2[11] == dec_i0_match_data_0[11]; // @[el2_lib.scala 197:80]
  wire  _T_234 = _T_230 | _T_233; // @[el2_lib.scala 197:25]
  wire  _T_236 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_237 = _T_236 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_240 = io_trigger_pkt_any_0_tdata2[12] == dec_i0_match_data_0[12]; // @[el2_lib.scala 197:80]
  wire  _T_241 = _T_237 | _T_240; // @[el2_lib.scala 197:25]
  wire  _T_243 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_244 = _T_243 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_247 = io_trigger_pkt_any_0_tdata2[13] == dec_i0_match_data_0[13]; // @[el2_lib.scala 197:80]
  wire  _T_248 = _T_244 | _T_247; // @[el2_lib.scala 197:25]
  wire  _T_250 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_251 = _T_250 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_254 = io_trigger_pkt_any_0_tdata2[14] == dec_i0_match_data_0[14]; // @[el2_lib.scala 197:80]
  wire  _T_255 = _T_251 | _T_254; // @[el2_lib.scala 197:25]
  wire  _T_257 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_258 = _T_257 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_261 = io_trigger_pkt_any_0_tdata2[15] == dec_i0_match_data_0[15]; // @[el2_lib.scala 197:80]
  wire  _T_262 = _T_258 | _T_261; // @[el2_lib.scala 197:25]
  wire  _T_264 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_265 = _T_264 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_268 = io_trigger_pkt_any_0_tdata2[16] == dec_i0_match_data_0[16]; // @[el2_lib.scala 197:80]
  wire  _T_269 = _T_265 | _T_268; // @[el2_lib.scala 197:25]
  wire  _T_271 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_272 = _T_271 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_275 = io_trigger_pkt_any_0_tdata2[17] == dec_i0_match_data_0[17]; // @[el2_lib.scala 197:80]
  wire  _T_276 = _T_272 | _T_275; // @[el2_lib.scala 197:25]
  wire  _T_278 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_279 = _T_278 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_282 = io_trigger_pkt_any_0_tdata2[18] == dec_i0_match_data_0[18]; // @[el2_lib.scala 197:80]
  wire  _T_283 = _T_279 | _T_282; // @[el2_lib.scala 197:25]
  wire  _T_285 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_286 = _T_285 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_289 = io_trigger_pkt_any_0_tdata2[19] == dec_i0_match_data_0[19]; // @[el2_lib.scala 197:80]
  wire  _T_290 = _T_286 | _T_289; // @[el2_lib.scala 197:25]
  wire  _T_292 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_293 = _T_292 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_296 = io_trigger_pkt_any_0_tdata2[20] == dec_i0_match_data_0[20]; // @[el2_lib.scala 197:80]
  wire  _T_297 = _T_293 | _T_296; // @[el2_lib.scala 197:25]
  wire  _T_299 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_300 = _T_299 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_303 = io_trigger_pkt_any_0_tdata2[21] == dec_i0_match_data_0[21]; // @[el2_lib.scala 197:80]
  wire  _T_304 = _T_300 | _T_303; // @[el2_lib.scala 197:25]
  wire  _T_306 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_307 = _T_306 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_310 = io_trigger_pkt_any_0_tdata2[22] == dec_i0_match_data_0[22]; // @[el2_lib.scala 197:80]
  wire  _T_311 = _T_307 | _T_310; // @[el2_lib.scala 197:25]
  wire  _T_313 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_314 = _T_313 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_317 = io_trigger_pkt_any_0_tdata2[23] == dec_i0_match_data_0[23]; // @[el2_lib.scala 197:80]
  wire  _T_318 = _T_314 | _T_317; // @[el2_lib.scala 197:25]
  wire  _T_320 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_321 = _T_320 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_324 = io_trigger_pkt_any_0_tdata2[24] == dec_i0_match_data_0[24]; // @[el2_lib.scala 197:80]
  wire  _T_325 = _T_321 | _T_324; // @[el2_lib.scala 197:25]
  wire  _T_327 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_328 = _T_327 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_331 = io_trigger_pkt_any_0_tdata2[25] == dec_i0_match_data_0[25]; // @[el2_lib.scala 197:80]
  wire  _T_332 = _T_328 | _T_331; // @[el2_lib.scala 197:25]
  wire  _T_334 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_335 = _T_334 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_338 = io_trigger_pkt_any_0_tdata2[26] == dec_i0_match_data_0[26]; // @[el2_lib.scala 197:80]
  wire  _T_339 = _T_335 | _T_338; // @[el2_lib.scala 197:25]
  wire  _T_341 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_342 = _T_341 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_345 = io_trigger_pkt_any_0_tdata2[27] == dec_i0_match_data_0[27]; // @[el2_lib.scala 197:80]
  wire  _T_346 = _T_342 | _T_345; // @[el2_lib.scala 197:25]
  wire  _T_348 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_349 = _T_348 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_352 = io_trigger_pkt_any_0_tdata2[28] == dec_i0_match_data_0[28]; // @[el2_lib.scala 197:80]
  wire  _T_353 = _T_349 | _T_352; // @[el2_lib.scala 197:25]
  wire  _T_355 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_356 = _T_355 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_359 = io_trigger_pkt_any_0_tdata2[29] == dec_i0_match_data_0[29]; // @[el2_lib.scala 197:80]
  wire  _T_360 = _T_356 | _T_359; // @[el2_lib.scala 197:25]
  wire  _T_362 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_363 = _T_362 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_366 = io_trigger_pkt_any_0_tdata2[30] == dec_i0_match_data_0[30]; // @[el2_lib.scala 197:80]
  wire  _T_367 = _T_363 | _T_366; // @[el2_lib.scala 197:25]
  wire  _T_369 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_370 = _T_369 & _T_153; // @[el2_lib.scala 197:43]
  wire  _T_373 = io_trigger_pkt_any_0_tdata2[31] == dec_i0_match_data_0[31]; // @[el2_lib.scala 197:80]
  wire  _T_374 = _T_370 | _T_373; // @[el2_lib.scala 197:25]
  wire  _T_375 = _T_157 & _T_164; // @[el2_lib.scala 198:22]
  wire  _T_376 = _T_375 & _T_171; // @[el2_lib.scala 198:22]
  wire  _T_377 = _T_376 & _T_178; // @[el2_lib.scala 198:22]
  wire  _T_378 = _T_377 & _T_185; // @[el2_lib.scala 198:22]
  wire  _T_379 = _T_378 & _T_192; // @[el2_lib.scala 198:22]
  wire  _T_380 = _T_379 & _T_199; // @[el2_lib.scala 198:22]
  wire  _T_381 = _T_380 & _T_206; // @[el2_lib.scala 198:22]
  wire  _T_382 = _T_381 & _T_213; // @[el2_lib.scala 198:22]
  wire  _T_383 = _T_382 & _T_220; // @[el2_lib.scala 198:22]
  wire  _T_384 = _T_383 & _T_227; // @[el2_lib.scala 198:22]
  wire  _T_385 = _T_384 & _T_234; // @[el2_lib.scala 198:22]
  wire  _T_386 = _T_385 & _T_241; // @[el2_lib.scala 198:22]
  wire  _T_387 = _T_386 & _T_248; // @[el2_lib.scala 198:22]
  wire  _T_388 = _T_387 & _T_255; // @[el2_lib.scala 198:22]
  wire  _T_389 = _T_388 & _T_262; // @[el2_lib.scala 198:22]
  wire  _T_390 = _T_389 & _T_269; // @[el2_lib.scala 198:22]
  wire  _T_391 = _T_390 & _T_276; // @[el2_lib.scala 198:22]
  wire  _T_392 = _T_391 & _T_283; // @[el2_lib.scala 198:22]
  wire  _T_393 = _T_392 & _T_290; // @[el2_lib.scala 198:22]
  wire  _T_394 = _T_393 & _T_297; // @[el2_lib.scala 198:22]
  wire  _T_395 = _T_394 & _T_304; // @[el2_lib.scala 198:22]
  wire  _T_396 = _T_395 & _T_311; // @[el2_lib.scala 198:22]
  wire  _T_397 = _T_396 & _T_318; // @[el2_lib.scala 198:22]
  wire  _T_398 = _T_397 & _T_325; // @[el2_lib.scala 198:22]
  wire  _T_399 = _T_398 & _T_332; // @[el2_lib.scala 198:22]
  wire  _T_400 = _T_399 & _T_339; // @[el2_lib.scala 198:22]
  wire  _T_401 = _T_400 & _T_346; // @[el2_lib.scala 198:22]
  wire  _T_402 = _T_401 & _T_353; // @[el2_lib.scala 198:22]
  wire  _T_403 = _T_402 & _T_360; // @[el2_lib.scala 198:22]
  wire  _T_404 = _T_403 & _T_367; // @[el2_lib.scala 198:22]
  wire  _T_405 = _T_404 & _T_374; // @[el2_lib.scala 198:22]
  wire  _T_406 = _T_148 & _T_405; // @[el2_lsu_trigger.scala 16:109]
  wire  _T_407 = io_trigger_pkt_any_1_execute & io_trigger_pkt_any_1_m; // @[el2_lsu_trigger.scala 16:83]
  wire  _T_410 = &io_trigger_pkt_any_1_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_411 = ~_T_410; // @[el2_lib.scala 194:39]
  wire  _T_412 = io_trigger_pkt_any_1_match_ & _T_411; // @[el2_lib.scala 194:37]
  wire  _T_415 = io_trigger_pkt_any_1_tdata2[0] == dec_i0_match_data_1[0]; // @[el2_lib.scala 195:52]
  wire  _T_416 = _T_412 | _T_415; // @[el2_lib.scala 195:41]
  wire  _T_418 = &io_trigger_pkt_any_1_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_419 = _T_418 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_422 = io_trigger_pkt_any_1_tdata2[1] == dec_i0_match_data_1[1]; // @[el2_lib.scala 197:80]
  wire  _T_423 = _T_419 | _T_422; // @[el2_lib.scala 197:25]
  wire  _T_425 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_426 = _T_425 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_429 = io_trigger_pkt_any_1_tdata2[2] == dec_i0_match_data_1[2]; // @[el2_lib.scala 197:80]
  wire  _T_430 = _T_426 | _T_429; // @[el2_lib.scala 197:25]
  wire  _T_432 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_433 = _T_432 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_436 = io_trigger_pkt_any_1_tdata2[3] == dec_i0_match_data_1[3]; // @[el2_lib.scala 197:80]
  wire  _T_437 = _T_433 | _T_436; // @[el2_lib.scala 197:25]
  wire  _T_439 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_440 = _T_439 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_443 = io_trigger_pkt_any_1_tdata2[4] == dec_i0_match_data_1[4]; // @[el2_lib.scala 197:80]
  wire  _T_444 = _T_440 | _T_443; // @[el2_lib.scala 197:25]
  wire  _T_446 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_447 = _T_446 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_450 = io_trigger_pkt_any_1_tdata2[5] == dec_i0_match_data_1[5]; // @[el2_lib.scala 197:80]
  wire  _T_451 = _T_447 | _T_450; // @[el2_lib.scala 197:25]
  wire  _T_453 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_454 = _T_453 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_457 = io_trigger_pkt_any_1_tdata2[6] == dec_i0_match_data_1[6]; // @[el2_lib.scala 197:80]
  wire  _T_458 = _T_454 | _T_457; // @[el2_lib.scala 197:25]
  wire  _T_460 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_461 = _T_460 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_464 = io_trigger_pkt_any_1_tdata2[7] == dec_i0_match_data_1[7]; // @[el2_lib.scala 197:80]
  wire  _T_465 = _T_461 | _T_464; // @[el2_lib.scala 197:25]
  wire  _T_467 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_468 = _T_467 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_471 = io_trigger_pkt_any_1_tdata2[8] == dec_i0_match_data_1[8]; // @[el2_lib.scala 197:80]
  wire  _T_472 = _T_468 | _T_471; // @[el2_lib.scala 197:25]
  wire  _T_474 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_475 = _T_474 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_478 = io_trigger_pkt_any_1_tdata2[9] == dec_i0_match_data_1[9]; // @[el2_lib.scala 197:80]
  wire  _T_479 = _T_475 | _T_478; // @[el2_lib.scala 197:25]
  wire  _T_481 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_482 = _T_481 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_485 = io_trigger_pkt_any_1_tdata2[10] == dec_i0_match_data_1[10]; // @[el2_lib.scala 197:80]
  wire  _T_486 = _T_482 | _T_485; // @[el2_lib.scala 197:25]
  wire  _T_488 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_489 = _T_488 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_492 = io_trigger_pkt_any_1_tdata2[11] == dec_i0_match_data_1[11]; // @[el2_lib.scala 197:80]
  wire  _T_493 = _T_489 | _T_492; // @[el2_lib.scala 197:25]
  wire  _T_495 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_496 = _T_495 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_499 = io_trigger_pkt_any_1_tdata2[12] == dec_i0_match_data_1[12]; // @[el2_lib.scala 197:80]
  wire  _T_500 = _T_496 | _T_499; // @[el2_lib.scala 197:25]
  wire  _T_502 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_503 = _T_502 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_506 = io_trigger_pkt_any_1_tdata2[13] == dec_i0_match_data_1[13]; // @[el2_lib.scala 197:80]
  wire  _T_507 = _T_503 | _T_506; // @[el2_lib.scala 197:25]
  wire  _T_509 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_510 = _T_509 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_513 = io_trigger_pkt_any_1_tdata2[14] == dec_i0_match_data_1[14]; // @[el2_lib.scala 197:80]
  wire  _T_514 = _T_510 | _T_513; // @[el2_lib.scala 197:25]
  wire  _T_516 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_517 = _T_516 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_520 = io_trigger_pkt_any_1_tdata2[15] == dec_i0_match_data_1[15]; // @[el2_lib.scala 197:80]
  wire  _T_521 = _T_517 | _T_520; // @[el2_lib.scala 197:25]
  wire  _T_523 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_524 = _T_523 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_527 = io_trigger_pkt_any_1_tdata2[16] == dec_i0_match_data_1[16]; // @[el2_lib.scala 197:80]
  wire  _T_528 = _T_524 | _T_527; // @[el2_lib.scala 197:25]
  wire  _T_530 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_531 = _T_530 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_534 = io_trigger_pkt_any_1_tdata2[17] == dec_i0_match_data_1[17]; // @[el2_lib.scala 197:80]
  wire  _T_535 = _T_531 | _T_534; // @[el2_lib.scala 197:25]
  wire  _T_537 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_538 = _T_537 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_541 = io_trigger_pkt_any_1_tdata2[18] == dec_i0_match_data_1[18]; // @[el2_lib.scala 197:80]
  wire  _T_542 = _T_538 | _T_541; // @[el2_lib.scala 197:25]
  wire  _T_544 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_545 = _T_544 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_548 = io_trigger_pkt_any_1_tdata2[19] == dec_i0_match_data_1[19]; // @[el2_lib.scala 197:80]
  wire  _T_549 = _T_545 | _T_548; // @[el2_lib.scala 197:25]
  wire  _T_551 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_552 = _T_551 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_555 = io_trigger_pkt_any_1_tdata2[20] == dec_i0_match_data_1[20]; // @[el2_lib.scala 197:80]
  wire  _T_556 = _T_552 | _T_555; // @[el2_lib.scala 197:25]
  wire  _T_558 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_559 = _T_558 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_562 = io_trigger_pkt_any_1_tdata2[21] == dec_i0_match_data_1[21]; // @[el2_lib.scala 197:80]
  wire  _T_563 = _T_559 | _T_562; // @[el2_lib.scala 197:25]
  wire  _T_565 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_566 = _T_565 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_569 = io_trigger_pkt_any_1_tdata2[22] == dec_i0_match_data_1[22]; // @[el2_lib.scala 197:80]
  wire  _T_570 = _T_566 | _T_569; // @[el2_lib.scala 197:25]
  wire  _T_572 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_573 = _T_572 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_576 = io_trigger_pkt_any_1_tdata2[23] == dec_i0_match_data_1[23]; // @[el2_lib.scala 197:80]
  wire  _T_577 = _T_573 | _T_576; // @[el2_lib.scala 197:25]
  wire  _T_579 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_580 = _T_579 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_583 = io_trigger_pkt_any_1_tdata2[24] == dec_i0_match_data_1[24]; // @[el2_lib.scala 197:80]
  wire  _T_584 = _T_580 | _T_583; // @[el2_lib.scala 197:25]
  wire  _T_586 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_587 = _T_586 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_590 = io_trigger_pkt_any_1_tdata2[25] == dec_i0_match_data_1[25]; // @[el2_lib.scala 197:80]
  wire  _T_591 = _T_587 | _T_590; // @[el2_lib.scala 197:25]
  wire  _T_593 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_594 = _T_593 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_597 = io_trigger_pkt_any_1_tdata2[26] == dec_i0_match_data_1[26]; // @[el2_lib.scala 197:80]
  wire  _T_598 = _T_594 | _T_597; // @[el2_lib.scala 197:25]
  wire  _T_600 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_601 = _T_600 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_604 = io_trigger_pkt_any_1_tdata2[27] == dec_i0_match_data_1[27]; // @[el2_lib.scala 197:80]
  wire  _T_605 = _T_601 | _T_604; // @[el2_lib.scala 197:25]
  wire  _T_607 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_608 = _T_607 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_611 = io_trigger_pkt_any_1_tdata2[28] == dec_i0_match_data_1[28]; // @[el2_lib.scala 197:80]
  wire  _T_612 = _T_608 | _T_611; // @[el2_lib.scala 197:25]
  wire  _T_614 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_615 = _T_614 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_618 = io_trigger_pkt_any_1_tdata2[29] == dec_i0_match_data_1[29]; // @[el2_lib.scala 197:80]
  wire  _T_619 = _T_615 | _T_618; // @[el2_lib.scala 197:25]
  wire  _T_621 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_622 = _T_621 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_625 = io_trigger_pkt_any_1_tdata2[30] == dec_i0_match_data_1[30]; // @[el2_lib.scala 197:80]
  wire  _T_626 = _T_622 | _T_625; // @[el2_lib.scala 197:25]
  wire  _T_628 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_629 = _T_628 & _T_412; // @[el2_lib.scala 197:43]
  wire  _T_632 = io_trigger_pkt_any_1_tdata2[31] == dec_i0_match_data_1[31]; // @[el2_lib.scala 197:80]
  wire  _T_633 = _T_629 | _T_632; // @[el2_lib.scala 197:25]
  wire  _T_634 = _T_416 & _T_423; // @[el2_lib.scala 198:22]
  wire  _T_635 = _T_634 & _T_430; // @[el2_lib.scala 198:22]
  wire  _T_636 = _T_635 & _T_437; // @[el2_lib.scala 198:22]
  wire  _T_637 = _T_636 & _T_444; // @[el2_lib.scala 198:22]
  wire  _T_638 = _T_637 & _T_451; // @[el2_lib.scala 198:22]
  wire  _T_639 = _T_638 & _T_458; // @[el2_lib.scala 198:22]
  wire  _T_640 = _T_639 & _T_465; // @[el2_lib.scala 198:22]
  wire  _T_641 = _T_640 & _T_472; // @[el2_lib.scala 198:22]
  wire  _T_642 = _T_641 & _T_479; // @[el2_lib.scala 198:22]
  wire  _T_643 = _T_642 & _T_486; // @[el2_lib.scala 198:22]
  wire  _T_644 = _T_643 & _T_493; // @[el2_lib.scala 198:22]
  wire  _T_645 = _T_644 & _T_500; // @[el2_lib.scala 198:22]
  wire  _T_646 = _T_645 & _T_507; // @[el2_lib.scala 198:22]
  wire  _T_647 = _T_646 & _T_514; // @[el2_lib.scala 198:22]
  wire  _T_648 = _T_647 & _T_521; // @[el2_lib.scala 198:22]
  wire  _T_649 = _T_648 & _T_528; // @[el2_lib.scala 198:22]
  wire  _T_650 = _T_649 & _T_535; // @[el2_lib.scala 198:22]
  wire  _T_651 = _T_650 & _T_542; // @[el2_lib.scala 198:22]
  wire  _T_652 = _T_651 & _T_549; // @[el2_lib.scala 198:22]
  wire  _T_653 = _T_652 & _T_556; // @[el2_lib.scala 198:22]
  wire  _T_654 = _T_653 & _T_563; // @[el2_lib.scala 198:22]
  wire  _T_655 = _T_654 & _T_570; // @[el2_lib.scala 198:22]
  wire  _T_656 = _T_655 & _T_577; // @[el2_lib.scala 198:22]
  wire  _T_657 = _T_656 & _T_584; // @[el2_lib.scala 198:22]
  wire  _T_658 = _T_657 & _T_591; // @[el2_lib.scala 198:22]
  wire  _T_659 = _T_658 & _T_598; // @[el2_lib.scala 198:22]
  wire  _T_660 = _T_659 & _T_605; // @[el2_lib.scala 198:22]
  wire  _T_661 = _T_660 & _T_612; // @[el2_lib.scala 198:22]
  wire  _T_662 = _T_661 & _T_619; // @[el2_lib.scala 198:22]
  wire  _T_663 = _T_662 & _T_626; // @[el2_lib.scala 198:22]
  wire  _T_664 = _T_663 & _T_633; // @[el2_lib.scala 198:22]
  wire  _T_665 = _T_407 & _T_664; // @[el2_lsu_trigger.scala 16:109]
  wire  _T_666 = io_trigger_pkt_any_2_execute & io_trigger_pkt_any_2_m; // @[el2_lsu_trigger.scala 16:83]
  wire  _T_669 = &io_trigger_pkt_any_2_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_670 = ~_T_669; // @[el2_lib.scala 194:39]
  wire  _T_671 = io_trigger_pkt_any_2_match_ & _T_670; // @[el2_lib.scala 194:37]
  wire  _T_674 = io_trigger_pkt_any_2_tdata2[0] == dec_i0_match_data_2[0]; // @[el2_lib.scala 195:52]
  wire  _T_675 = _T_671 | _T_674; // @[el2_lib.scala 195:41]
  wire  _T_677 = &io_trigger_pkt_any_2_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_678 = _T_677 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_681 = io_trigger_pkt_any_2_tdata2[1] == dec_i0_match_data_2[1]; // @[el2_lib.scala 197:80]
  wire  _T_682 = _T_678 | _T_681; // @[el2_lib.scala 197:25]
  wire  _T_684 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_685 = _T_684 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_688 = io_trigger_pkt_any_2_tdata2[2] == dec_i0_match_data_2[2]; // @[el2_lib.scala 197:80]
  wire  _T_689 = _T_685 | _T_688; // @[el2_lib.scala 197:25]
  wire  _T_691 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_692 = _T_691 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_695 = io_trigger_pkt_any_2_tdata2[3] == dec_i0_match_data_2[3]; // @[el2_lib.scala 197:80]
  wire  _T_696 = _T_692 | _T_695; // @[el2_lib.scala 197:25]
  wire  _T_698 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_699 = _T_698 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_702 = io_trigger_pkt_any_2_tdata2[4] == dec_i0_match_data_2[4]; // @[el2_lib.scala 197:80]
  wire  _T_703 = _T_699 | _T_702; // @[el2_lib.scala 197:25]
  wire  _T_705 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_706 = _T_705 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_709 = io_trigger_pkt_any_2_tdata2[5] == dec_i0_match_data_2[5]; // @[el2_lib.scala 197:80]
  wire  _T_710 = _T_706 | _T_709; // @[el2_lib.scala 197:25]
  wire  _T_712 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_713 = _T_712 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_716 = io_trigger_pkt_any_2_tdata2[6] == dec_i0_match_data_2[6]; // @[el2_lib.scala 197:80]
  wire  _T_717 = _T_713 | _T_716; // @[el2_lib.scala 197:25]
  wire  _T_719 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_720 = _T_719 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_723 = io_trigger_pkt_any_2_tdata2[7] == dec_i0_match_data_2[7]; // @[el2_lib.scala 197:80]
  wire  _T_724 = _T_720 | _T_723; // @[el2_lib.scala 197:25]
  wire  _T_726 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_727 = _T_726 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_730 = io_trigger_pkt_any_2_tdata2[8] == dec_i0_match_data_2[8]; // @[el2_lib.scala 197:80]
  wire  _T_731 = _T_727 | _T_730; // @[el2_lib.scala 197:25]
  wire  _T_733 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_734 = _T_733 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_737 = io_trigger_pkt_any_2_tdata2[9] == dec_i0_match_data_2[9]; // @[el2_lib.scala 197:80]
  wire  _T_738 = _T_734 | _T_737; // @[el2_lib.scala 197:25]
  wire  _T_740 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_741 = _T_740 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_744 = io_trigger_pkt_any_2_tdata2[10] == dec_i0_match_data_2[10]; // @[el2_lib.scala 197:80]
  wire  _T_745 = _T_741 | _T_744; // @[el2_lib.scala 197:25]
  wire  _T_747 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_748 = _T_747 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_751 = io_trigger_pkt_any_2_tdata2[11] == dec_i0_match_data_2[11]; // @[el2_lib.scala 197:80]
  wire  _T_752 = _T_748 | _T_751; // @[el2_lib.scala 197:25]
  wire  _T_754 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_755 = _T_754 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_758 = io_trigger_pkt_any_2_tdata2[12] == dec_i0_match_data_2[12]; // @[el2_lib.scala 197:80]
  wire  _T_759 = _T_755 | _T_758; // @[el2_lib.scala 197:25]
  wire  _T_761 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_762 = _T_761 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_765 = io_trigger_pkt_any_2_tdata2[13] == dec_i0_match_data_2[13]; // @[el2_lib.scala 197:80]
  wire  _T_766 = _T_762 | _T_765; // @[el2_lib.scala 197:25]
  wire  _T_768 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_769 = _T_768 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_772 = io_trigger_pkt_any_2_tdata2[14] == dec_i0_match_data_2[14]; // @[el2_lib.scala 197:80]
  wire  _T_773 = _T_769 | _T_772; // @[el2_lib.scala 197:25]
  wire  _T_775 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_776 = _T_775 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_779 = io_trigger_pkt_any_2_tdata2[15] == dec_i0_match_data_2[15]; // @[el2_lib.scala 197:80]
  wire  _T_780 = _T_776 | _T_779; // @[el2_lib.scala 197:25]
  wire  _T_782 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_783 = _T_782 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_786 = io_trigger_pkt_any_2_tdata2[16] == dec_i0_match_data_2[16]; // @[el2_lib.scala 197:80]
  wire  _T_787 = _T_783 | _T_786; // @[el2_lib.scala 197:25]
  wire  _T_789 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_790 = _T_789 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_793 = io_trigger_pkt_any_2_tdata2[17] == dec_i0_match_data_2[17]; // @[el2_lib.scala 197:80]
  wire  _T_794 = _T_790 | _T_793; // @[el2_lib.scala 197:25]
  wire  _T_796 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_797 = _T_796 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_800 = io_trigger_pkt_any_2_tdata2[18] == dec_i0_match_data_2[18]; // @[el2_lib.scala 197:80]
  wire  _T_801 = _T_797 | _T_800; // @[el2_lib.scala 197:25]
  wire  _T_803 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_804 = _T_803 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_807 = io_trigger_pkt_any_2_tdata2[19] == dec_i0_match_data_2[19]; // @[el2_lib.scala 197:80]
  wire  _T_808 = _T_804 | _T_807; // @[el2_lib.scala 197:25]
  wire  _T_810 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_811 = _T_810 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_814 = io_trigger_pkt_any_2_tdata2[20] == dec_i0_match_data_2[20]; // @[el2_lib.scala 197:80]
  wire  _T_815 = _T_811 | _T_814; // @[el2_lib.scala 197:25]
  wire  _T_817 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_818 = _T_817 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_821 = io_trigger_pkt_any_2_tdata2[21] == dec_i0_match_data_2[21]; // @[el2_lib.scala 197:80]
  wire  _T_822 = _T_818 | _T_821; // @[el2_lib.scala 197:25]
  wire  _T_824 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_825 = _T_824 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_828 = io_trigger_pkt_any_2_tdata2[22] == dec_i0_match_data_2[22]; // @[el2_lib.scala 197:80]
  wire  _T_829 = _T_825 | _T_828; // @[el2_lib.scala 197:25]
  wire  _T_831 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_832 = _T_831 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_835 = io_trigger_pkt_any_2_tdata2[23] == dec_i0_match_data_2[23]; // @[el2_lib.scala 197:80]
  wire  _T_836 = _T_832 | _T_835; // @[el2_lib.scala 197:25]
  wire  _T_838 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_839 = _T_838 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_842 = io_trigger_pkt_any_2_tdata2[24] == dec_i0_match_data_2[24]; // @[el2_lib.scala 197:80]
  wire  _T_843 = _T_839 | _T_842; // @[el2_lib.scala 197:25]
  wire  _T_845 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_846 = _T_845 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_849 = io_trigger_pkt_any_2_tdata2[25] == dec_i0_match_data_2[25]; // @[el2_lib.scala 197:80]
  wire  _T_850 = _T_846 | _T_849; // @[el2_lib.scala 197:25]
  wire  _T_852 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_853 = _T_852 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_856 = io_trigger_pkt_any_2_tdata2[26] == dec_i0_match_data_2[26]; // @[el2_lib.scala 197:80]
  wire  _T_857 = _T_853 | _T_856; // @[el2_lib.scala 197:25]
  wire  _T_859 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_860 = _T_859 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_863 = io_trigger_pkt_any_2_tdata2[27] == dec_i0_match_data_2[27]; // @[el2_lib.scala 197:80]
  wire  _T_864 = _T_860 | _T_863; // @[el2_lib.scala 197:25]
  wire  _T_866 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_867 = _T_866 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_870 = io_trigger_pkt_any_2_tdata2[28] == dec_i0_match_data_2[28]; // @[el2_lib.scala 197:80]
  wire  _T_871 = _T_867 | _T_870; // @[el2_lib.scala 197:25]
  wire  _T_873 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_874 = _T_873 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_877 = io_trigger_pkt_any_2_tdata2[29] == dec_i0_match_data_2[29]; // @[el2_lib.scala 197:80]
  wire  _T_878 = _T_874 | _T_877; // @[el2_lib.scala 197:25]
  wire  _T_880 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_881 = _T_880 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_884 = io_trigger_pkt_any_2_tdata2[30] == dec_i0_match_data_2[30]; // @[el2_lib.scala 197:80]
  wire  _T_885 = _T_881 | _T_884; // @[el2_lib.scala 197:25]
  wire  _T_887 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_888 = _T_887 & _T_671; // @[el2_lib.scala 197:43]
  wire  _T_891 = io_trigger_pkt_any_2_tdata2[31] == dec_i0_match_data_2[31]; // @[el2_lib.scala 197:80]
  wire  _T_892 = _T_888 | _T_891; // @[el2_lib.scala 197:25]
  wire  _T_893 = _T_675 & _T_682; // @[el2_lib.scala 198:22]
  wire  _T_894 = _T_893 & _T_689; // @[el2_lib.scala 198:22]
  wire  _T_895 = _T_894 & _T_696; // @[el2_lib.scala 198:22]
  wire  _T_896 = _T_895 & _T_703; // @[el2_lib.scala 198:22]
  wire  _T_897 = _T_896 & _T_710; // @[el2_lib.scala 198:22]
  wire  _T_898 = _T_897 & _T_717; // @[el2_lib.scala 198:22]
  wire  _T_899 = _T_898 & _T_724; // @[el2_lib.scala 198:22]
  wire  _T_900 = _T_899 & _T_731; // @[el2_lib.scala 198:22]
  wire  _T_901 = _T_900 & _T_738; // @[el2_lib.scala 198:22]
  wire  _T_902 = _T_901 & _T_745; // @[el2_lib.scala 198:22]
  wire  _T_903 = _T_902 & _T_752; // @[el2_lib.scala 198:22]
  wire  _T_904 = _T_903 & _T_759; // @[el2_lib.scala 198:22]
  wire  _T_905 = _T_904 & _T_766; // @[el2_lib.scala 198:22]
  wire  _T_906 = _T_905 & _T_773; // @[el2_lib.scala 198:22]
  wire  _T_907 = _T_906 & _T_780; // @[el2_lib.scala 198:22]
  wire  _T_908 = _T_907 & _T_787; // @[el2_lib.scala 198:22]
  wire  _T_909 = _T_908 & _T_794; // @[el2_lib.scala 198:22]
  wire  _T_910 = _T_909 & _T_801; // @[el2_lib.scala 198:22]
  wire  _T_911 = _T_910 & _T_808; // @[el2_lib.scala 198:22]
  wire  _T_912 = _T_911 & _T_815; // @[el2_lib.scala 198:22]
  wire  _T_913 = _T_912 & _T_822; // @[el2_lib.scala 198:22]
  wire  _T_914 = _T_913 & _T_829; // @[el2_lib.scala 198:22]
  wire  _T_915 = _T_914 & _T_836; // @[el2_lib.scala 198:22]
  wire  _T_916 = _T_915 & _T_843; // @[el2_lib.scala 198:22]
  wire  _T_917 = _T_916 & _T_850; // @[el2_lib.scala 198:22]
  wire  _T_918 = _T_917 & _T_857; // @[el2_lib.scala 198:22]
  wire  _T_919 = _T_918 & _T_864; // @[el2_lib.scala 198:22]
  wire  _T_920 = _T_919 & _T_871; // @[el2_lib.scala 198:22]
  wire  _T_921 = _T_920 & _T_878; // @[el2_lib.scala 198:22]
  wire  _T_922 = _T_921 & _T_885; // @[el2_lib.scala 198:22]
  wire  _T_923 = _T_922 & _T_892; // @[el2_lib.scala 198:22]
  wire  _T_924 = _T_666 & _T_923; // @[el2_lsu_trigger.scala 16:109]
  wire  _T_925 = io_trigger_pkt_any_3_execute & io_trigger_pkt_any_3_m; // @[el2_lsu_trigger.scala 16:83]
  wire  _T_928 = &io_trigger_pkt_any_3_tdata2; // @[el2_lib.scala 194:45]
  wire  _T_929 = ~_T_928; // @[el2_lib.scala 194:39]
  wire  _T_930 = io_trigger_pkt_any_3_match_ & _T_929; // @[el2_lib.scala 194:37]
  wire  _T_933 = io_trigger_pkt_any_3_tdata2[0] == dec_i0_match_data_3[0]; // @[el2_lib.scala 195:52]
  wire  _T_934 = _T_930 | _T_933; // @[el2_lib.scala 195:41]
  wire  _T_936 = &io_trigger_pkt_any_3_tdata2[0]; // @[el2_lib.scala 197:38]
  wire  _T_937 = _T_936 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_940 = io_trigger_pkt_any_3_tdata2[1] == dec_i0_match_data_3[1]; // @[el2_lib.scala 197:80]
  wire  _T_941 = _T_937 | _T_940; // @[el2_lib.scala 197:25]
  wire  _T_943 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[el2_lib.scala 197:38]
  wire  _T_944 = _T_943 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_947 = io_trigger_pkt_any_3_tdata2[2] == dec_i0_match_data_3[2]; // @[el2_lib.scala 197:80]
  wire  _T_948 = _T_944 | _T_947; // @[el2_lib.scala 197:25]
  wire  _T_950 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[el2_lib.scala 197:38]
  wire  _T_951 = _T_950 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_954 = io_trigger_pkt_any_3_tdata2[3] == dec_i0_match_data_3[3]; // @[el2_lib.scala 197:80]
  wire  _T_955 = _T_951 | _T_954; // @[el2_lib.scala 197:25]
  wire  _T_957 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[el2_lib.scala 197:38]
  wire  _T_958 = _T_957 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_961 = io_trigger_pkt_any_3_tdata2[4] == dec_i0_match_data_3[4]; // @[el2_lib.scala 197:80]
  wire  _T_962 = _T_958 | _T_961; // @[el2_lib.scala 197:25]
  wire  _T_964 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[el2_lib.scala 197:38]
  wire  _T_965 = _T_964 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_968 = io_trigger_pkt_any_3_tdata2[5] == dec_i0_match_data_3[5]; // @[el2_lib.scala 197:80]
  wire  _T_969 = _T_965 | _T_968; // @[el2_lib.scala 197:25]
  wire  _T_971 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[el2_lib.scala 197:38]
  wire  _T_972 = _T_971 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_975 = io_trigger_pkt_any_3_tdata2[6] == dec_i0_match_data_3[6]; // @[el2_lib.scala 197:80]
  wire  _T_976 = _T_972 | _T_975; // @[el2_lib.scala 197:25]
  wire  _T_978 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[el2_lib.scala 197:38]
  wire  _T_979 = _T_978 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_982 = io_trigger_pkt_any_3_tdata2[7] == dec_i0_match_data_3[7]; // @[el2_lib.scala 197:80]
  wire  _T_983 = _T_979 | _T_982; // @[el2_lib.scala 197:25]
  wire  _T_985 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[el2_lib.scala 197:38]
  wire  _T_986 = _T_985 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_989 = io_trigger_pkt_any_3_tdata2[8] == dec_i0_match_data_3[8]; // @[el2_lib.scala 197:80]
  wire  _T_990 = _T_986 | _T_989; // @[el2_lib.scala 197:25]
  wire  _T_992 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[el2_lib.scala 197:38]
  wire  _T_993 = _T_992 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_996 = io_trigger_pkt_any_3_tdata2[9] == dec_i0_match_data_3[9]; // @[el2_lib.scala 197:80]
  wire  _T_997 = _T_993 | _T_996; // @[el2_lib.scala 197:25]
  wire  _T_999 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[el2_lib.scala 197:38]
  wire  _T_1000 = _T_999 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1003 = io_trigger_pkt_any_3_tdata2[10] == dec_i0_match_data_3[10]; // @[el2_lib.scala 197:80]
  wire  _T_1004 = _T_1000 | _T_1003; // @[el2_lib.scala 197:25]
  wire  _T_1006 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[el2_lib.scala 197:38]
  wire  _T_1007 = _T_1006 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1010 = io_trigger_pkt_any_3_tdata2[11] == dec_i0_match_data_3[11]; // @[el2_lib.scala 197:80]
  wire  _T_1011 = _T_1007 | _T_1010; // @[el2_lib.scala 197:25]
  wire  _T_1013 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[el2_lib.scala 197:38]
  wire  _T_1014 = _T_1013 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1017 = io_trigger_pkt_any_3_tdata2[12] == dec_i0_match_data_3[12]; // @[el2_lib.scala 197:80]
  wire  _T_1018 = _T_1014 | _T_1017; // @[el2_lib.scala 197:25]
  wire  _T_1020 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[el2_lib.scala 197:38]
  wire  _T_1021 = _T_1020 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1024 = io_trigger_pkt_any_3_tdata2[13] == dec_i0_match_data_3[13]; // @[el2_lib.scala 197:80]
  wire  _T_1025 = _T_1021 | _T_1024; // @[el2_lib.scala 197:25]
  wire  _T_1027 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[el2_lib.scala 197:38]
  wire  _T_1028 = _T_1027 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1031 = io_trigger_pkt_any_3_tdata2[14] == dec_i0_match_data_3[14]; // @[el2_lib.scala 197:80]
  wire  _T_1032 = _T_1028 | _T_1031; // @[el2_lib.scala 197:25]
  wire  _T_1034 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[el2_lib.scala 197:38]
  wire  _T_1035 = _T_1034 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1038 = io_trigger_pkt_any_3_tdata2[15] == dec_i0_match_data_3[15]; // @[el2_lib.scala 197:80]
  wire  _T_1039 = _T_1035 | _T_1038; // @[el2_lib.scala 197:25]
  wire  _T_1041 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[el2_lib.scala 197:38]
  wire  _T_1042 = _T_1041 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1045 = io_trigger_pkt_any_3_tdata2[16] == dec_i0_match_data_3[16]; // @[el2_lib.scala 197:80]
  wire  _T_1046 = _T_1042 | _T_1045; // @[el2_lib.scala 197:25]
  wire  _T_1048 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[el2_lib.scala 197:38]
  wire  _T_1049 = _T_1048 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1052 = io_trigger_pkt_any_3_tdata2[17] == dec_i0_match_data_3[17]; // @[el2_lib.scala 197:80]
  wire  _T_1053 = _T_1049 | _T_1052; // @[el2_lib.scala 197:25]
  wire  _T_1055 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[el2_lib.scala 197:38]
  wire  _T_1056 = _T_1055 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1059 = io_trigger_pkt_any_3_tdata2[18] == dec_i0_match_data_3[18]; // @[el2_lib.scala 197:80]
  wire  _T_1060 = _T_1056 | _T_1059; // @[el2_lib.scala 197:25]
  wire  _T_1062 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[el2_lib.scala 197:38]
  wire  _T_1063 = _T_1062 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1066 = io_trigger_pkt_any_3_tdata2[19] == dec_i0_match_data_3[19]; // @[el2_lib.scala 197:80]
  wire  _T_1067 = _T_1063 | _T_1066; // @[el2_lib.scala 197:25]
  wire  _T_1069 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[el2_lib.scala 197:38]
  wire  _T_1070 = _T_1069 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1073 = io_trigger_pkt_any_3_tdata2[20] == dec_i0_match_data_3[20]; // @[el2_lib.scala 197:80]
  wire  _T_1074 = _T_1070 | _T_1073; // @[el2_lib.scala 197:25]
  wire  _T_1076 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[el2_lib.scala 197:38]
  wire  _T_1077 = _T_1076 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1080 = io_trigger_pkt_any_3_tdata2[21] == dec_i0_match_data_3[21]; // @[el2_lib.scala 197:80]
  wire  _T_1081 = _T_1077 | _T_1080; // @[el2_lib.scala 197:25]
  wire  _T_1083 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[el2_lib.scala 197:38]
  wire  _T_1084 = _T_1083 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1087 = io_trigger_pkt_any_3_tdata2[22] == dec_i0_match_data_3[22]; // @[el2_lib.scala 197:80]
  wire  _T_1088 = _T_1084 | _T_1087; // @[el2_lib.scala 197:25]
  wire  _T_1090 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[el2_lib.scala 197:38]
  wire  _T_1091 = _T_1090 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1094 = io_trigger_pkt_any_3_tdata2[23] == dec_i0_match_data_3[23]; // @[el2_lib.scala 197:80]
  wire  _T_1095 = _T_1091 | _T_1094; // @[el2_lib.scala 197:25]
  wire  _T_1097 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[el2_lib.scala 197:38]
  wire  _T_1098 = _T_1097 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1101 = io_trigger_pkt_any_3_tdata2[24] == dec_i0_match_data_3[24]; // @[el2_lib.scala 197:80]
  wire  _T_1102 = _T_1098 | _T_1101; // @[el2_lib.scala 197:25]
  wire  _T_1104 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[el2_lib.scala 197:38]
  wire  _T_1105 = _T_1104 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1108 = io_trigger_pkt_any_3_tdata2[25] == dec_i0_match_data_3[25]; // @[el2_lib.scala 197:80]
  wire  _T_1109 = _T_1105 | _T_1108; // @[el2_lib.scala 197:25]
  wire  _T_1111 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[el2_lib.scala 197:38]
  wire  _T_1112 = _T_1111 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1115 = io_trigger_pkt_any_3_tdata2[26] == dec_i0_match_data_3[26]; // @[el2_lib.scala 197:80]
  wire  _T_1116 = _T_1112 | _T_1115; // @[el2_lib.scala 197:25]
  wire  _T_1118 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[el2_lib.scala 197:38]
  wire  _T_1119 = _T_1118 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1122 = io_trigger_pkt_any_3_tdata2[27] == dec_i0_match_data_3[27]; // @[el2_lib.scala 197:80]
  wire  _T_1123 = _T_1119 | _T_1122; // @[el2_lib.scala 197:25]
  wire  _T_1125 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[el2_lib.scala 197:38]
  wire  _T_1126 = _T_1125 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1129 = io_trigger_pkt_any_3_tdata2[28] == dec_i0_match_data_3[28]; // @[el2_lib.scala 197:80]
  wire  _T_1130 = _T_1126 | _T_1129; // @[el2_lib.scala 197:25]
  wire  _T_1132 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[el2_lib.scala 197:38]
  wire  _T_1133 = _T_1132 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1136 = io_trigger_pkt_any_3_tdata2[29] == dec_i0_match_data_3[29]; // @[el2_lib.scala 197:80]
  wire  _T_1137 = _T_1133 | _T_1136; // @[el2_lib.scala 197:25]
  wire  _T_1139 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[el2_lib.scala 197:38]
  wire  _T_1140 = _T_1139 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1143 = io_trigger_pkt_any_3_tdata2[30] == dec_i0_match_data_3[30]; // @[el2_lib.scala 197:80]
  wire  _T_1144 = _T_1140 | _T_1143; // @[el2_lib.scala 197:25]
  wire  _T_1146 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[el2_lib.scala 197:38]
  wire  _T_1147 = _T_1146 & _T_930; // @[el2_lib.scala 197:43]
  wire  _T_1150 = io_trigger_pkt_any_3_tdata2[31] == dec_i0_match_data_3[31]; // @[el2_lib.scala 197:80]
  wire  _T_1151 = _T_1147 | _T_1150; // @[el2_lib.scala 197:25]
  wire  _T_1152 = _T_934 & _T_941; // @[el2_lib.scala 198:22]
  wire  _T_1153 = _T_1152 & _T_948; // @[el2_lib.scala 198:22]
  wire  _T_1154 = _T_1153 & _T_955; // @[el2_lib.scala 198:22]
  wire  _T_1155 = _T_1154 & _T_962; // @[el2_lib.scala 198:22]
  wire  _T_1156 = _T_1155 & _T_969; // @[el2_lib.scala 198:22]
  wire  _T_1157 = _T_1156 & _T_976; // @[el2_lib.scala 198:22]
  wire  _T_1158 = _T_1157 & _T_983; // @[el2_lib.scala 198:22]
  wire  _T_1159 = _T_1158 & _T_990; // @[el2_lib.scala 198:22]
  wire  _T_1160 = _T_1159 & _T_997; // @[el2_lib.scala 198:22]
  wire  _T_1161 = _T_1160 & _T_1004; // @[el2_lib.scala 198:22]
  wire  _T_1162 = _T_1161 & _T_1011; // @[el2_lib.scala 198:22]
  wire  _T_1163 = _T_1162 & _T_1018; // @[el2_lib.scala 198:22]
  wire  _T_1164 = _T_1163 & _T_1025; // @[el2_lib.scala 198:22]
  wire  _T_1165 = _T_1164 & _T_1032; // @[el2_lib.scala 198:22]
  wire  _T_1166 = _T_1165 & _T_1039; // @[el2_lib.scala 198:22]
  wire  _T_1167 = _T_1166 & _T_1046; // @[el2_lib.scala 198:22]
  wire  _T_1168 = _T_1167 & _T_1053; // @[el2_lib.scala 198:22]
  wire  _T_1169 = _T_1168 & _T_1060; // @[el2_lib.scala 198:22]
  wire  _T_1170 = _T_1169 & _T_1067; // @[el2_lib.scala 198:22]
  wire  _T_1171 = _T_1170 & _T_1074; // @[el2_lib.scala 198:22]
  wire  _T_1172 = _T_1171 & _T_1081; // @[el2_lib.scala 198:22]
  wire  _T_1173 = _T_1172 & _T_1088; // @[el2_lib.scala 198:22]
  wire  _T_1174 = _T_1173 & _T_1095; // @[el2_lib.scala 198:22]
  wire  _T_1175 = _T_1174 & _T_1102; // @[el2_lib.scala 198:22]
  wire  _T_1176 = _T_1175 & _T_1109; // @[el2_lib.scala 198:22]
  wire  _T_1177 = _T_1176 & _T_1116; // @[el2_lib.scala 198:22]
  wire  _T_1178 = _T_1177 & _T_1123; // @[el2_lib.scala 198:22]
  wire  _T_1179 = _T_1178 & _T_1130; // @[el2_lib.scala 198:22]
  wire  _T_1180 = _T_1179 & _T_1137; // @[el2_lib.scala 198:22]
  wire  _T_1181 = _T_1180 & _T_1144; // @[el2_lib.scala 198:22]
  wire  _T_1182 = _T_1181 & _T_1151; // @[el2_lib.scala 198:22]
  wire  _T_1183 = _T_925 & _T_1182; // @[el2_lsu_trigger.scala 16:109]
  wire [2:0] _T_1185 = {_T_1183,_T_924,_T_665}; // @[Cat.scala 29:58]
  assign io_dec_i0_trigger_match_d = {_T_1185,_T_406}; // @[el2_lsu_trigger.scala 16:29]
endmodule
