module el2_lsu_trigger(
  input         clock,
  input         reset,
  input         io_trigger_pkt_any_0_select,
  input         io_trigger_pkt_any_0_match_,
  input         io_trigger_pkt_any_0_store,
  input         io_trigger_pkt_any_0_load,
  input         io_trigger_pkt_any_0_execute,
  input         io_trigger_pkt_any_0_m,
  input  [31:0] io_trigger_pkt_any_0_tdata2,
  input         io_trigger_pkt_any_1_select,
  input         io_trigger_pkt_any_1_match_,
  input         io_trigger_pkt_any_1_store,
  input         io_trigger_pkt_any_1_load,
  input         io_trigger_pkt_any_1_execute,
  input         io_trigger_pkt_any_1_m,
  input  [31:0] io_trigger_pkt_any_1_tdata2,
  input         io_trigger_pkt_any_2_select,
  input         io_trigger_pkt_any_2_match_,
  input         io_trigger_pkt_any_2_store,
  input         io_trigger_pkt_any_2_load,
  input         io_trigger_pkt_any_2_execute,
  input         io_trigger_pkt_any_2_m,
  input  [31:0] io_trigger_pkt_any_2_tdata2,
  input         io_trigger_pkt_any_3_select,
  input         io_trigger_pkt_any_3_match_,
  input         io_trigger_pkt_any_3_store,
  input         io_trigger_pkt_any_3_load,
  input         io_trigger_pkt_any_3_execute,
  input         io_trigger_pkt_any_3_m,
  input  [31:0] io_trigger_pkt_any_3_tdata2,
  input         io_lsu_pkt_m_fast_int,
  input         io_lsu_pkt_m_by,
  input         io_lsu_pkt_m_half,
  input         io_lsu_pkt_m_word,
  input         io_lsu_pkt_m_dword,
  input         io_lsu_pkt_m_load,
  input         io_lsu_pkt_m_store,
  input         io_lsu_pkt_m_unsign,
  input         io_lsu_pkt_m_dma,
  input         io_lsu_pkt_m_store_data_bypass_d,
  input         io_lsu_pkt_m_load_ldst_bypass_d,
  input         io_lsu_pkt_m_store_data_bypass_m,
  input         io_lsu_pkt_m_valid,
  input  [31:0] io_lsu_addr_m,
  input  [31:0] io_store_data_m,
  output [3:0]  io_lsu_trigger_match_m
);
  wire [15:0] _T_1 = io_lsu_pkt_m_word ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _T_3 = _T_1 & io_store_data_m[31:16]; // @[el2_lsu_trigger.scala 16:61]
  wire  _T_4 = io_lsu_pkt_m_half | io_lsu_pkt_m_word; // @[el2_lsu_trigger.scala 16:114]
  wire [7:0] _T_6 = _T_4 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_8 = _T_6 & io_store_data_m[15:8]; // @[el2_lsu_trigger.scala 16:136]
  wire [31:0] store_data_trigger_m = {_T_3,_T_8,io_store_data_m[7:0]}; // @[Cat.scala 29:58]
  wire  _T_12 = ~io_trigger_pkt_any_0_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_13 = io_trigger_pkt_any_0_select & io_trigger_pkt_any_0_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_15 = _T_12 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_16 = _T_13 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_0 = _T_15 | _T_16; // @[Mux.scala 27:72]
  wire  _T_19 = ~io_trigger_pkt_any_1_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_20 = io_trigger_pkt_any_1_select & io_trigger_pkt_any_1_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_22 = _T_19 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_23 = _T_20 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_1 = _T_22 | _T_23; // @[Mux.scala 27:72]
  wire  _T_26 = ~io_trigger_pkt_any_2_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_27 = io_trigger_pkt_any_2_select & io_trigger_pkt_any_2_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_29 = _T_26 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_30 = _T_27 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_2 = _T_29 | _T_30; // @[Mux.scala 27:72]
  wire  _T_33 = ~io_trigger_pkt_any_3_select; // @[el2_lsu_trigger.scala 17:53]
  wire  _T_34 = io_trigger_pkt_any_3_select & io_trigger_pkt_any_3_store; // @[el2_lsu_trigger.scala 17:136]
  wire [31:0] _T_36 = _T_33 ? io_lsu_addr_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_37 = _T_34 ? store_data_trigger_m : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] lsu_match_data_3 = _T_36 | _T_37; // @[Mux.scala 27:72]
  wire  _T_39 = ~io_lsu_pkt_m_dma; // @[el2_lsu_trigger.scala 18:71]
  wire  _T_40 = io_lsu_pkt_m_valid & _T_39; // @[el2_lsu_trigger.scala 18:69]
  wire  _T_41 = io_trigger_pkt_any_0_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 18:121]
  wire  _T_42 = io_trigger_pkt_any_0_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_44 = _T_42 & _T_12; // @[el2_lsu_trigger.scala 19:53]
  wire  _T_45 = _T_41 | _T_44; // @[el2_lsu_trigger.scala 18:142]
  wire  _T_46 = _T_40 & _T_45; // @[el2_lsu_trigger.scala 18:89]
  wire  _T_51 = &io_trigger_pkt_any_0_tdata2; // @[el2_lib.scala 240:73]
  wire  _T_52 = ~_T_51; // @[el2_lib.scala 240:47]
  wire  _T_53 = io_trigger_pkt_any_0_match_ & _T_52; // @[el2_lib.scala 240:44]
  wire  _T_56 = io_trigger_pkt_any_0_tdata2[0] == lsu_match_data_0[0]; // @[el2_lib.scala 241:52]
  wire  _T_57 = _T_53 | _T_56; // @[el2_lib.scala 241:41]
  wire  _T_59 = &io_trigger_pkt_any_0_tdata2[0]; // @[el2_lib.scala 243:37]
  wire  _T_60 = _T_59 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_63 = io_trigger_pkt_any_0_tdata2[1] == lsu_match_data_0[1]; // @[el2_lib.scala 243:79]
  wire  _T_64 = _T_60 | _T_63; // @[el2_lib.scala 243:24]
  wire  _T_66 = &io_trigger_pkt_any_0_tdata2[1:0]; // @[el2_lib.scala 243:37]
  wire  _T_67 = _T_66 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_70 = io_trigger_pkt_any_0_tdata2[2] == lsu_match_data_0[2]; // @[el2_lib.scala 243:79]
  wire  _T_71 = _T_67 | _T_70; // @[el2_lib.scala 243:24]
  wire  _T_73 = &io_trigger_pkt_any_0_tdata2[2:0]; // @[el2_lib.scala 243:37]
  wire  _T_74 = _T_73 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_77 = io_trigger_pkt_any_0_tdata2[3] == lsu_match_data_0[3]; // @[el2_lib.scala 243:79]
  wire  _T_78 = _T_74 | _T_77; // @[el2_lib.scala 243:24]
  wire  _T_80 = &io_trigger_pkt_any_0_tdata2[3:0]; // @[el2_lib.scala 243:37]
  wire  _T_81 = _T_80 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_84 = io_trigger_pkt_any_0_tdata2[4] == lsu_match_data_0[4]; // @[el2_lib.scala 243:79]
  wire  _T_85 = _T_81 | _T_84; // @[el2_lib.scala 243:24]
  wire  _T_87 = &io_trigger_pkt_any_0_tdata2[4:0]; // @[el2_lib.scala 243:37]
  wire  _T_88 = _T_87 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_91 = io_trigger_pkt_any_0_tdata2[5] == lsu_match_data_0[5]; // @[el2_lib.scala 243:79]
  wire  _T_92 = _T_88 | _T_91; // @[el2_lib.scala 243:24]
  wire  _T_94 = &io_trigger_pkt_any_0_tdata2[5:0]; // @[el2_lib.scala 243:37]
  wire  _T_95 = _T_94 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_98 = io_trigger_pkt_any_0_tdata2[6] == lsu_match_data_0[6]; // @[el2_lib.scala 243:79]
  wire  _T_99 = _T_95 | _T_98; // @[el2_lib.scala 243:24]
  wire  _T_101 = &io_trigger_pkt_any_0_tdata2[6:0]; // @[el2_lib.scala 243:37]
  wire  _T_102 = _T_101 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_105 = io_trigger_pkt_any_0_tdata2[7] == lsu_match_data_0[7]; // @[el2_lib.scala 243:79]
  wire  _T_106 = _T_102 | _T_105; // @[el2_lib.scala 243:24]
  wire  _T_108 = &io_trigger_pkt_any_0_tdata2[7:0]; // @[el2_lib.scala 243:37]
  wire  _T_109 = _T_108 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_112 = io_trigger_pkt_any_0_tdata2[8] == lsu_match_data_0[8]; // @[el2_lib.scala 243:79]
  wire  _T_113 = _T_109 | _T_112; // @[el2_lib.scala 243:24]
  wire  _T_115 = &io_trigger_pkt_any_0_tdata2[8:0]; // @[el2_lib.scala 243:37]
  wire  _T_116 = _T_115 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_119 = io_trigger_pkt_any_0_tdata2[9] == lsu_match_data_0[9]; // @[el2_lib.scala 243:79]
  wire  _T_120 = _T_116 | _T_119; // @[el2_lib.scala 243:24]
  wire  _T_122 = &io_trigger_pkt_any_0_tdata2[9:0]; // @[el2_lib.scala 243:37]
  wire  _T_123 = _T_122 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_126 = io_trigger_pkt_any_0_tdata2[10] == lsu_match_data_0[10]; // @[el2_lib.scala 243:79]
  wire  _T_127 = _T_123 | _T_126; // @[el2_lib.scala 243:24]
  wire  _T_129 = &io_trigger_pkt_any_0_tdata2[10:0]; // @[el2_lib.scala 243:37]
  wire  _T_130 = _T_129 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_133 = io_trigger_pkt_any_0_tdata2[11] == lsu_match_data_0[11]; // @[el2_lib.scala 243:79]
  wire  _T_134 = _T_130 | _T_133; // @[el2_lib.scala 243:24]
  wire  _T_136 = &io_trigger_pkt_any_0_tdata2[11:0]; // @[el2_lib.scala 243:37]
  wire  _T_137 = _T_136 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_140 = io_trigger_pkt_any_0_tdata2[12] == lsu_match_data_0[12]; // @[el2_lib.scala 243:79]
  wire  _T_141 = _T_137 | _T_140; // @[el2_lib.scala 243:24]
  wire  _T_143 = &io_trigger_pkt_any_0_tdata2[12:0]; // @[el2_lib.scala 243:37]
  wire  _T_144 = _T_143 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_147 = io_trigger_pkt_any_0_tdata2[13] == lsu_match_data_0[13]; // @[el2_lib.scala 243:79]
  wire  _T_148 = _T_144 | _T_147; // @[el2_lib.scala 243:24]
  wire  _T_150 = &io_trigger_pkt_any_0_tdata2[13:0]; // @[el2_lib.scala 243:37]
  wire  _T_151 = _T_150 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_154 = io_trigger_pkt_any_0_tdata2[14] == lsu_match_data_0[14]; // @[el2_lib.scala 243:79]
  wire  _T_155 = _T_151 | _T_154; // @[el2_lib.scala 243:24]
  wire  _T_157 = &io_trigger_pkt_any_0_tdata2[14:0]; // @[el2_lib.scala 243:37]
  wire  _T_158 = _T_157 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_161 = io_trigger_pkt_any_0_tdata2[15] == lsu_match_data_0[15]; // @[el2_lib.scala 243:79]
  wire  _T_162 = _T_158 | _T_161; // @[el2_lib.scala 243:24]
  wire  _T_164 = &io_trigger_pkt_any_0_tdata2[15:0]; // @[el2_lib.scala 243:37]
  wire  _T_165 = _T_164 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_168 = io_trigger_pkt_any_0_tdata2[16] == lsu_match_data_0[16]; // @[el2_lib.scala 243:79]
  wire  _T_169 = _T_165 | _T_168; // @[el2_lib.scala 243:24]
  wire  _T_171 = &io_trigger_pkt_any_0_tdata2[16:0]; // @[el2_lib.scala 243:37]
  wire  _T_172 = _T_171 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_175 = io_trigger_pkt_any_0_tdata2[17] == lsu_match_data_0[17]; // @[el2_lib.scala 243:79]
  wire  _T_176 = _T_172 | _T_175; // @[el2_lib.scala 243:24]
  wire  _T_178 = &io_trigger_pkt_any_0_tdata2[17:0]; // @[el2_lib.scala 243:37]
  wire  _T_179 = _T_178 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_182 = io_trigger_pkt_any_0_tdata2[18] == lsu_match_data_0[18]; // @[el2_lib.scala 243:79]
  wire  _T_183 = _T_179 | _T_182; // @[el2_lib.scala 243:24]
  wire  _T_185 = &io_trigger_pkt_any_0_tdata2[18:0]; // @[el2_lib.scala 243:37]
  wire  _T_186 = _T_185 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_189 = io_trigger_pkt_any_0_tdata2[19] == lsu_match_data_0[19]; // @[el2_lib.scala 243:79]
  wire  _T_190 = _T_186 | _T_189; // @[el2_lib.scala 243:24]
  wire  _T_192 = &io_trigger_pkt_any_0_tdata2[19:0]; // @[el2_lib.scala 243:37]
  wire  _T_193 = _T_192 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_196 = io_trigger_pkt_any_0_tdata2[20] == lsu_match_data_0[20]; // @[el2_lib.scala 243:79]
  wire  _T_197 = _T_193 | _T_196; // @[el2_lib.scala 243:24]
  wire  _T_199 = &io_trigger_pkt_any_0_tdata2[20:0]; // @[el2_lib.scala 243:37]
  wire  _T_200 = _T_199 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_203 = io_trigger_pkt_any_0_tdata2[21] == lsu_match_data_0[21]; // @[el2_lib.scala 243:79]
  wire  _T_204 = _T_200 | _T_203; // @[el2_lib.scala 243:24]
  wire  _T_206 = &io_trigger_pkt_any_0_tdata2[21:0]; // @[el2_lib.scala 243:37]
  wire  _T_207 = _T_206 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_210 = io_trigger_pkt_any_0_tdata2[22] == lsu_match_data_0[22]; // @[el2_lib.scala 243:79]
  wire  _T_211 = _T_207 | _T_210; // @[el2_lib.scala 243:24]
  wire  _T_213 = &io_trigger_pkt_any_0_tdata2[22:0]; // @[el2_lib.scala 243:37]
  wire  _T_214 = _T_213 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_217 = io_trigger_pkt_any_0_tdata2[23] == lsu_match_data_0[23]; // @[el2_lib.scala 243:79]
  wire  _T_218 = _T_214 | _T_217; // @[el2_lib.scala 243:24]
  wire  _T_220 = &io_trigger_pkt_any_0_tdata2[23:0]; // @[el2_lib.scala 243:37]
  wire  _T_221 = _T_220 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_224 = io_trigger_pkt_any_0_tdata2[24] == lsu_match_data_0[24]; // @[el2_lib.scala 243:79]
  wire  _T_225 = _T_221 | _T_224; // @[el2_lib.scala 243:24]
  wire  _T_227 = &io_trigger_pkt_any_0_tdata2[24:0]; // @[el2_lib.scala 243:37]
  wire  _T_228 = _T_227 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_231 = io_trigger_pkt_any_0_tdata2[25] == lsu_match_data_0[25]; // @[el2_lib.scala 243:79]
  wire  _T_232 = _T_228 | _T_231; // @[el2_lib.scala 243:24]
  wire  _T_234 = &io_trigger_pkt_any_0_tdata2[25:0]; // @[el2_lib.scala 243:37]
  wire  _T_235 = _T_234 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_238 = io_trigger_pkt_any_0_tdata2[26] == lsu_match_data_0[26]; // @[el2_lib.scala 243:79]
  wire  _T_239 = _T_235 | _T_238; // @[el2_lib.scala 243:24]
  wire  _T_241 = &io_trigger_pkt_any_0_tdata2[26:0]; // @[el2_lib.scala 243:37]
  wire  _T_242 = _T_241 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_245 = io_trigger_pkt_any_0_tdata2[27] == lsu_match_data_0[27]; // @[el2_lib.scala 243:79]
  wire  _T_246 = _T_242 | _T_245; // @[el2_lib.scala 243:24]
  wire  _T_248 = &io_trigger_pkt_any_0_tdata2[27:0]; // @[el2_lib.scala 243:37]
  wire  _T_249 = _T_248 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_252 = io_trigger_pkt_any_0_tdata2[28] == lsu_match_data_0[28]; // @[el2_lib.scala 243:79]
  wire  _T_253 = _T_249 | _T_252; // @[el2_lib.scala 243:24]
  wire  _T_255 = &io_trigger_pkt_any_0_tdata2[28:0]; // @[el2_lib.scala 243:37]
  wire  _T_256 = _T_255 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_259 = io_trigger_pkt_any_0_tdata2[29] == lsu_match_data_0[29]; // @[el2_lib.scala 243:79]
  wire  _T_260 = _T_256 | _T_259; // @[el2_lib.scala 243:24]
  wire  _T_262 = &io_trigger_pkt_any_0_tdata2[29:0]; // @[el2_lib.scala 243:37]
  wire  _T_263 = _T_262 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_266 = io_trigger_pkt_any_0_tdata2[30] == lsu_match_data_0[30]; // @[el2_lib.scala 243:79]
  wire  _T_267 = _T_263 | _T_266; // @[el2_lib.scala 243:24]
  wire  _T_269 = &io_trigger_pkt_any_0_tdata2[30:0]; // @[el2_lib.scala 243:37]
  wire  _T_270 = _T_269 & _T_53; // @[el2_lib.scala 243:42]
  wire  _T_273 = io_trigger_pkt_any_0_tdata2[31] == lsu_match_data_0[31]; // @[el2_lib.scala 243:79]
  wire  _T_274 = _T_270 | _T_273; // @[el2_lib.scala 243:24]
  wire [7:0] _T_281 = {_T_106,_T_99,_T_92,_T_85,_T_78,_T_71,_T_64,_T_57}; // @[el2_lib.scala 244:14]
  wire [15:0] _T_289 = {_T_162,_T_155,_T_148,_T_141,_T_134,_T_127,_T_120,_T_113,_T_281}; // @[el2_lib.scala 244:14]
  wire [7:0] _T_296 = {_T_218,_T_211,_T_204,_T_197,_T_190,_T_183,_T_176,_T_169}; // @[el2_lib.scala 244:14]
  wire [31:0] _T_305 = {_T_274,_T_267,_T_260,_T_253,_T_246,_T_239,_T_232,_T_225,_T_296,_T_289}; // @[el2_lib.scala 244:14]
  wire  _T_306 = &_T_305; // @[el2_lib.scala 244:21]
  wire  _T_307 = _T_46 & _T_306; // @[el2_lsu_trigger.scala 19:87]
  wire  _T_310 = io_trigger_pkt_any_1_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 18:121]
  wire  _T_311 = io_trigger_pkt_any_1_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_313 = _T_311 & _T_19; // @[el2_lsu_trigger.scala 19:53]
  wire  _T_314 = _T_310 | _T_313; // @[el2_lsu_trigger.scala 18:142]
  wire  _T_315 = _T_40 & _T_314; // @[el2_lsu_trigger.scala 18:89]
  wire  _T_320 = &io_trigger_pkt_any_1_tdata2; // @[el2_lib.scala 240:73]
  wire  _T_321 = ~_T_320; // @[el2_lib.scala 240:47]
  wire  _T_322 = io_trigger_pkt_any_1_match_ & _T_321; // @[el2_lib.scala 240:44]
  wire  _T_325 = io_trigger_pkt_any_1_tdata2[0] == lsu_match_data_1[0]; // @[el2_lib.scala 241:52]
  wire  _T_326 = _T_322 | _T_325; // @[el2_lib.scala 241:41]
  wire  _T_328 = &io_trigger_pkt_any_1_tdata2[0]; // @[el2_lib.scala 243:37]
  wire  _T_329 = _T_328 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_332 = io_trigger_pkt_any_1_tdata2[1] == lsu_match_data_1[1]; // @[el2_lib.scala 243:79]
  wire  _T_333 = _T_329 | _T_332; // @[el2_lib.scala 243:24]
  wire  _T_335 = &io_trigger_pkt_any_1_tdata2[1:0]; // @[el2_lib.scala 243:37]
  wire  _T_336 = _T_335 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_339 = io_trigger_pkt_any_1_tdata2[2] == lsu_match_data_1[2]; // @[el2_lib.scala 243:79]
  wire  _T_340 = _T_336 | _T_339; // @[el2_lib.scala 243:24]
  wire  _T_342 = &io_trigger_pkt_any_1_tdata2[2:0]; // @[el2_lib.scala 243:37]
  wire  _T_343 = _T_342 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_346 = io_trigger_pkt_any_1_tdata2[3] == lsu_match_data_1[3]; // @[el2_lib.scala 243:79]
  wire  _T_347 = _T_343 | _T_346; // @[el2_lib.scala 243:24]
  wire  _T_349 = &io_trigger_pkt_any_1_tdata2[3:0]; // @[el2_lib.scala 243:37]
  wire  _T_350 = _T_349 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_353 = io_trigger_pkt_any_1_tdata2[4] == lsu_match_data_1[4]; // @[el2_lib.scala 243:79]
  wire  _T_354 = _T_350 | _T_353; // @[el2_lib.scala 243:24]
  wire  _T_356 = &io_trigger_pkt_any_1_tdata2[4:0]; // @[el2_lib.scala 243:37]
  wire  _T_357 = _T_356 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_360 = io_trigger_pkt_any_1_tdata2[5] == lsu_match_data_1[5]; // @[el2_lib.scala 243:79]
  wire  _T_361 = _T_357 | _T_360; // @[el2_lib.scala 243:24]
  wire  _T_363 = &io_trigger_pkt_any_1_tdata2[5:0]; // @[el2_lib.scala 243:37]
  wire  _T_364 = _T_363 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_367 = io_trigger_pkt_any_1_tdata2[6] == lsu_match_data_1[6]; // @[el2_lib.scala 243:79]
  wire  _T_368 = _T_364 | _T_367; // @[el2_lib.scala 243:24]
  wire  _T_370 = &io_trigger_pkt_any_1_tdata2[6:0]; // @[el2_lib.scala 243:37]
  wire  _T_371 = _T_370 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_374 = io_trigger_pkt_any_1_tdata2[7] == lsu_match_data_1[7]; // @[el2_lib.scala 243:79]
  wire  _T_375 = _T_371 | _T_374; // @[el2_lib.scala 243:24]
  wire  _T_377 = &io_trigger_pkt_any_1_tdata2[7:0]; // @[el2_lib.scala 243:37]
  wire  _T_378 = _T_377 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_381 = io_trigger_pkt_any_1_tdata2[8] == lsu_match_data_1[8]; // @[el2_lib.scala 243:79]
  wire  _T_382 = _T_378 | _T_381; // @[el2_lib.scala 243:24]
  wire  _T_384 = &io_trigger_pkt_any_1_tdata2[8:0]; // @[el2_lib.scala 243:37]
  wire  _T_385 = _T_384 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_388 = io_trigger_pkt_any_1_tdata2[9] == lsu_match_data_1[9]; // @[el2_lib.scala 243:79]
  wire  _T_389 = _T_385 | _T_388; // @[el2_lib.scala 243:24]
  wire  _T_391 = &io_trigger_pkt_any_1_tdata2[9:0]; // @[el2_lib.scala 243:37]
  wire  _T_392 = _T_391 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_395 = io_trigger_pkt_any_1_tdata2[10] == lsu_match_data_1[10]; // @[el2_lib.scala 243:79]
  wire  _T_396 = _T_392 | _T_395; // @[el2_lib.scala 243:24]
  wire  _T_398 = &io_trigger_pkt_any_1_tdata2[10:0]; // @[el2_lib.scala 243:37]
  wire  _T_399 = _T_398 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_402 = io_trigger_pkt_any_1_tdata2[11] == lsu_match_data_1[11]; // @[el2_lib.scala 243:79]
  wire  _T_403 = _T_399 | _T_402; // @[el2_lib.scala 243:24]
  wire  _T_405 = &io_trigger_pkt_any_1_tdata2[11:0]; // @[el2_lib.scala 243:37]
  wire  _T_406 = _T_405 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_409 = io_trigger_pkt_any_1_tdata2[12] == lsu_match_data_1[12]; // @[el2_lib.scala 243:79]
  wire  _T_410 = _T_406 | _T_409; // @[el2_lib.scala 243:24]
  wire  _T_412 = &io_trigger_pkt_any_1_tdata2[12:0]; // @[el2_lib.scala 243:37]
  wire  _T_413 = _T_412 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_416 = io_trigger_pkt_any_1_tdata2[13] == lsu_match_data_1[13]; // @[el2_lib.scala 243:79]
  wire  _T_417 = _T_413 | _T_416; // @[el2_lib.scala 243:24]
  wire  _T_419 = &io_trigger_pkt_any_1_tdata2[13:0]; // @[el2_lib.scala 243:37]
  wire  _T_420 = _T_419 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_423 = io_trigger_pkt_any_1_tdata2[14] == lsu_match_data_1[14]; // @[el2_lib.scala 243:79]
  wire  _T_424 = _T_420 | _T_423; // @[el2_lib.scala 243:24]
  wire  _T_426 = &io_trigger_pkt_any_1_tdata2[14:0]; // @[el2_lib.scala 243:37]
  wire  _T_427 = _T_426 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_430 = io_trigger_pkt_any_1_tdata2[15] == lsu_match_data_1[15]; // @[el2_lib.scala 243:79]
  wire  _T_431 = _T_427 | _T_430; // @[el2_lib.scala 243:24]
  wire  _T_433 = &io_trigger_pkt_any_1_tdata2[15:0]; // @[el2_lib.scala 243:37]
  wire  _T_434 = _T_433 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_437 = io_trigger_pkt_any_1_tdata2[16] == lsu_match_data_1[16]; // @[el2_lib.scala 243:79]
  wire  _T_438 = _T_434 | _T_437; // @[el2_lib.scala 243:24]
  wire  _T_440 = &io_trigger_pkt_any_1_tdata2[16:0]; // @[el2_lib.scala 243:37]
  wire  _T_441 = _T_440 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_444 = io_trigger_pkt_any_1_tdata2[17] == lsu_match_data_1[17]; // @[el2_lib.scala 243:79]
  wire  _T_445 = _T_441 | _T_444; // @[el2_lib.scala 243:24]
  wire  _T_447 = &io_trigger_pkt_any_1_tdata2[17:0]; // @[el2_lib.scala 243:37]
  wire  _T_448 = _T_447 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_451 = io_trigger_pkt_any_1_tdata2[18] == lsu_match_data_1[18]; // @[el2_lib.scala 243:79]
  wire  _T_452 = _T_448 | _T_451; // @[el2_lib.scala 243:24]
  wire  _T_454 = &io_trigger_pkt_any_1_tdata2[18:0]; // @[el2_lib.scala 243:37]
  wire  _T_455 = _T_454 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_458 = io_trigger_pkt_any_1_tdata2[19] == lsu_match_data_1[19]; // @[el2_lib.scala 243:79]
  wire  _T_459 = _T_455 | _T_458; // @[el2_lib.scala 243:24]
  wire  _T_461 = &io_trigger_pkt_any_1_tdata2[19:0]; // @[el2_lib.scala 243:37]
  wire  _T_462 = _T_461 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_465 = io_trigger_pkt_any_1_tdata2[20] == lsu_match_data_1[20]; // @[el2_lib.scala 243:79]
  wire  _T_466 = _T_462 | _T_465; // @[el2_lib.scala 243:24]
  wire  _T_468 = &io_trigger_pkt_any_1_tdata2[20:0]; // @[el2_lib.scala 243:37]
  wire  _T_469 = _T_468 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_472 = io_trigger_pkt_any_1_tdata2[21] == lsu_match_data_1[21]; // @[el2_lib.scala 243:79]
  wire  _T_473 = _T_469 | _T_472; // @[el2_lib.scala 243:24]
  wire  _T_475 = &io_trigger_pkt_any_1_tdata2[21:0]; // @[el2_lib.scala 243:37]
  wire  _T_476 = _T_475 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_479 = io_trigger_pkt_any_1_tdata2[22] == lsu_match_data_1[22]; // @[el2_lib.scala 243:79]
  wire  _T_480 = _T_476 | _T_479; // @[el2_lib.scala 243:24]
  wire  _T_482 = &io_trigger_pkt_any_1_tdata2[22:0]; // @[el2_lib.scala 243:37]
  wire  _T_483 = _T_482 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_486 = io_trigger_pkt_any_1_tdata2[23] == lsu_match_data_1[23]; // @[el2_lib.scala 243:79]
  wire  _T_487 = _T_483 | _T_486; // @[el2_lib.scala 243:24]
  wire  _T_489 = &io_trigger_pkt_any_1_tdata2[23:0]; // @[el2_lib.scala 243:37]
  wire  _T_490 = _T_489 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_493 = io_trigger_pkt_any_1_tdata2[24] == lsu_match_data_1[24]; // @[el2_lib.scala 243:79]
  wire  _T_494 = _T_490 | _T_493; // @[el2_lib.scala 243:24]
  wire  _T_496 = &io_trigger_pkt_any_1_tdata2[24:0]; // @[el2_lib.scala 243:37]
  wire  _T_497 = _T_496 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_500 = io_trigger_pkt_any_1_tdata2[25] == lsu_match_data_1[25]; // @[el2_lib.scala 243:79]
  wire  _T_501 = _T_497 | _T_500; // @[el2_lib.scala 243:24]
  wire  _T_503 = &io_trigger_pkt_any_1_tdata2[25:0]; // @[el2_lib.scala 243:37]
  wire  _T_504 = _T_503 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_507 = io_trigger_pkt_any_1_tdata2[26] == lsu_match_data_1[26]; // @[el2_lib.scala 243:79]
  wire  _T_508 = _T_504 | _T_507; // @[el2_lib.scala 243:24]
  wire  _T_510 = &io_trigger_pkt_any_1_tdata2[26:0]; // @[el2_lib.scala 243:37]
  wire  _T_511 = _T_510 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_514 = io_trigger_pkt_any_1_tdata2[27] == lsu_match_data_1[27]; // @[el2_lib.scala 243:79]
  wire  _T_515 = _T_511 | _T_514; // @[el2_lib.scala 243:24]
  wire  _T_517 = &io_trigger_pkt_any_1_tdata2[27:0]; // @[el2_lib.scala 243:37]
  wire  _T_518 = _T_517 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_521 = io_trigger_pkt_any_1_tdata2[28] == lsu_match_data_1[28]; // @[el2_lib.scala 243:79]
  wire  _T_522 = _T_518 | _T_521; // @[el2_lib.scala 243:24]
  wire  _T_524 = &io_trigger_pkt_any_1_tdata2[28:0]; // @[el2_lib.scala 243:37]
  wire  _T_525 = _T_524 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_528 = io_trigger_pkt_any_1_tdata2[29] == lsu_match_data_1[29]; // @[el2_lib.scala 243:79]
  wire  _T_529 = _T_525 | _T_528; // @[el2_lib.scala 243:24]
  wire  _T_531 = &io_trigger_pkt_any_1_tdata2[29:0]; // @[el2_lib.scala 243:37]
  wire  _T_532 = _T_531 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_535 = io_trigger_pkt_any_1_tdata2[30] == lsu_match_data_1[30]; // @[el2_lib.scala 243:79]
  wire  _T_536 = _T_532 | _T_535; // @[el2_lib.scala 243:24]
  wire  _T_538 = &io_trigger_pkt_any_1_tdata2[30:0]; // @[el2_lib.scala 243:37]
  wire  _T_539 = _T_538 & _T_322; // @[el2_lib.scala 243:42]
  wire  _T_542 = io_trigger_pkt_any_1_tdata2[31] == lsu_match_data_1[31]; // @[el2_lib.scala 243:79]
  wire  _T_543 = _T_539 | _T_542; // @[el2_lib.scala 243:24]
  wire [7:0] _T_550 = {_T_375,_T_368,_T_361,_T_354,_T_347,_T_340,_T_333,_T_326}; // @[el2_lib.scala 244:14]
  wire [15:0] _T_558 = {_T_431,_T_424,_T_417,_T_410,_T_403,_T_396,_T_389,_T_382,_T_550}; // @[el2_lib.scala 244:14]
  wire [7:0] _T_565 = {_T_487,_T_480,_T_473,_T_466,_T_459,_T_452,_T_445,_T_438}; // @[el2_lib.scala 244:14]
  wire [31:0] _T_574 = {_T_543,_T_536,_T_529,_T_522,_T_515,_T_508,_T_501,_T_494,_T_565,_T_558}; // @[el2_lib.scala 244:14]
  wire  _T_575 = &_T_574; // @[el2_lib.scala 244:21]
  wire  _T_576 = _T_315 & _T_575; // @[el2_lsu_trigger.scala 19:87]
  wire  _T_579 = io_trigger_pkt_any_2_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 18:121]
  wire  _T_580 = io_trigger_pkt_any_2_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_582 = _T_580 & _T_26; // @[el2_lsu_trigger.scala 19:53]
  wire  _T_583 = _T_579 | _T_582; // @[el2_lsu_trigger.scala 18:142]
  wire  _T_584 = _T_40 & _T_583; // @[el2_lsu_trigger.scala 18:89]
  wire  _T_589 = &io_trigger_pkt_any_2_tdata2; // @[el2_lib.scala 240:73]
  wire  _T_590 = ~_T_589; // @[el2_lib.scala 240:47]
  wire  _T_591 = io_trigger_pkt_any_2_match_ & _T_590; // @[el2_lib.scala 240:44]
  wire  _T_594 = io_trigger_pkt_any_2_tdata2[0] == lsu_match_data_2[0]; // @[el2_lib.scala 241:52]
  wire  _T_595 = _T_591 | _T_594; // @[el2_lib.scala 241:41]
  wire  _T_597 = &io_trigger_pkt_any_2_tdata2[0]; // @[el2_lib.scala 243:37]
  wire  _T_598 = _T_597 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_601 = io_trigger_pkt_any_2_tdata2[1] == lsu_match_data_2[1]; // @[el2_lib.scala 243:79]
  wire  _T_602 = _T_598 | _T_601; // @[el2_lib.scala 243:24]
  wire  _T_604 = &io_trigger_pkt_any_2_tdata2[1:0]; // @[el2_lib.scala 243:37]
  wire  _T_605 = _T_604 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_608 = io_trigger_pkt_any_2_tdata2[2] == lsu_match_data_2[2]; // @[el2_lib.scala 243:79]
  wire  _T_609 = _T_605 | _T_608; // @[el2_lib.scala 243:24]
  wire  _T_611 = &io_trigger_pkt_any_2_tdata2[2:0]; // @[el2_lib.scala 243:37]
  wire  _T_612 = _T_611 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_615 = io_trigger_pkt_any_2_tdata2[3] == lsu_match_data_2[3]; // @[el2_lib.scala 243:79]
  wire  _T_616 = _T_612 | _T_615; // @[el2_lib.scala 243:24]
  wire  _T_618 = &io_trigger_pkt_any_2_tdata2[3:0]; // @[el2_lib.scala 243:37]
  wire  _T_619 = _T_618 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_622 = io_trigger_pkt_any_2_tdata2[4] == lsu_match_data_2[4]; // @[el2_lib.scala 243:79]
  wire  _T_623 = _T_619 | _T_622; // @[el2_lib.scala 243:24]
  wire  _T_625 = &io_trigger_pkt_any_2_tdata2[4:0]; // @[el2_lib.scala 243:37]
  wire  _T_626 = _T_625 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_629 = io_trigger_pkt_any_2_tdata2[5] == lsu_match_data_2[5]; // @[el2_lib.scala 243:79]
  wire  _T_630 = _T_626 | _T_629; // @[el2_lib.scala 243:24]
  wire  _T_632 = &io_trigger_pkt_any_2_tdata2[5:0]; // @[el2_lib.scala 243:37]
  wire  _T_633 = _T_632 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_636 = io_trigger_pkt_any_2_tdata2[6] == lsu_match_data_2[6]; // @[el2_lib.scala 243:79]
  wire  _T_637 = _T_633 | _T_636; // @[el2_lib.scala 243:24]
  wire  _T_639 = &io_trigger_pkt_any_2_tdata2[6:0]; // @[el2_lib.scala 243:37]
  wire  _T_640 = _T_639 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_643 = io_trigger_pkt_any_2_tdata2[7] == lsu_match_data_2[7]; // @[el2_lib.scala 243:79]
  wire  _T_644 = _T_640 | _T_643; // @[el2_lib.scala 243:24]
  wire  _T_646 = &io_trigger_pkt_any_2_tdata2[7:0]; // @[el2_lib.scala 243:37]
  wire  _T_647 = _T_646 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_650 = io_trigger_pkt_any_2_tdata2[8] == lsu_match_data_2[8]; // @[el2_lib.scala 243:79]
  wire  _T_651 = _T_647 | _T_650; // @[el2_lib.scala 243:24]
  wire  _T_653 = &io_trigger_pkt_any_2_tdata2[8:0]; // @[el2_lib.scala 243:37]
  wire  _T_654 = _T_653 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_657 = io_trigger_pkt_any_2_tdata2[9] == lsu_match_data_2[9]; // @[el2_lib.scala 243:79]
  wire  _T_658 = _T_654 | _T_657; // @[el2_lib.scala 243:24]
  wire  _T_660 = &io_trigger_pkt_any_2_tdata2[9:0]; // @[el2_lib.scala 243:37]
  wire  _T_661 = _T_660 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_664 = io_trigger_pkt_any_2_tdata2[10] == lsu_match_data_2[10]; // @[el2_lib.scala 243:79]
  wire  _T_665 = _T_661 | _T_664; // @[el2_lib.scala 243:24]
  wire  _T_667 = &io_trigger_pkt_any_2_tdata2[10:0]; // @[el2_lib.scala 243:37]
  wire  _T_668 = _T_667 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_671 = io_trigger_pkt_any_2_tdata2[11] == lsu_match_data_2[11]; // @[el2_lib.scala 243:79]
  wire  _T_672 = _T_668 | _T_671; // @[el2_lib.scala 243:24]
  wire  _T_674 = &io_trigger_pkt_any_2_tdata2[11:0]; // @[el2_lib.scala 243:37]
  wire  _T_675 = _T_674 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_678 = io_trigger_pkt_any_2_tdata2[12] == lsu_match_data_2[12]; // @[el2_lib.scala 243:79]
  wire  _T_679 = _T_675 | _T_678; // @[el2_lib.scala 243:24]
  wire  _T_681 = &io_trigger_pkt_any_2_tdata2[12:0]; // @[el2_lib.scala 243:37]
  wire  _T_682 = _T_681 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_685 = io_trigger_pkt_any_2_tdata2[13] == lsu_match_data_2[13]; // @[el2_lib.scala 243:79]
  wire  _T_686 = _T_682 | _T_685; // @[el2_lib.scala 243:24]
  wire  _T_688 = &io_trigger_pkt_any_2_tdata2[13:0]; // @[el2_lib.scala 243:37]
  wire  _T_689 = _T_688 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_692 = io_trigger_pkt_any_2_tdata2[14] == lsu_match_data_2[14]; // @[el2_lib.scala 243:79]
  wire  _T_693 = _T_689 | _T_692; // @[el2_lib.scala 243:24]
  wire  _T_695 = &io_trigger_pkt_any_2_tdata2[14:0]; // @[el2_lib.scala 243:37]
  wire  _T_696 = _T_695 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_699 = io_trigger_pkt_any_2_tdata2[15] == lsu_match_data_2[15]; // @[el2_lib.scala 243:79]
  wire  _T_700 = _T_696 | _T_699; // @[el2_lib.scala 243:24]
  wire  _T_702 = &io_trigger_pkt_any_2_tdata2[15:0]; // @[el2_lib.scala 243:37]
  wire  _T_703 = _T_702 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_706 = io_trigger_pkt_any_2_tdata2[16] == lsu_match_data_2[16]; // @[el2_lib.scala 243:79]
  wire  _T_707 = _T_703 | _T_706; // @[el2_lib.scala 243:24]
  wire  _T_709 = &io_trigger_pkt_any_2_tdata2[16:0]; // @[el2_lib.scala 243:37]
  wire  _T_710 = _T_709 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_713 = io_trigger_pkt_any_2_tdata2[17] == lsu_match_data_2[17]; // @[el2_lib.scala 243:79]
  wire  _T_714 = _T_710 | _T_713; // @[el2_lib.scala 243:24]
  wire  _T_716 = &io_trigger_pkt_any_2_tdata2[17:0]; // @[el2_lib.scala 243:37]
  wire  _T_717 = _T_716 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_720 = io_trigger_pkt_any_2_tdata2[18] == lsu_match_data_2[18]; // @[el2_lib.scala 243:79]
  wire  _T_721 = _T_717 | _T_720; // @[el2_lib.scala 243:24]
  wire  _T_723 = &io_trigger_pkt_any_2_tdata2[18:0]; // @[el2_lib.scala 243:37]
  wire  _T_724 = _T_723 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_727 = io_trigger_pkt_any_2_tdata2[19] == lsu_match_data_2[19]; // @[el2_lib.scala 243:79]
  wire  _T_728 = _T_724 | _T_727; // @[el2_lib.scala 243:24]
  wire  _T_730 = &io_trigger_pkt_any_2_tdata2[19:0]; // @[el2_lib.scala 243:37]
  wire  _T_731 = _T_730 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_734 = io_trigger_pkt_any_2_tdata2[20] == lsu_match_data_2[20]; // @[el2_lib.scala 243:79]
  wire  _T_735 = _T_731 | _T_734; // @[el2_lib.scala 243:24]
  wire  _T_737 = &io_trigger_pkt_any_2_tdata2[20:0]; // @[el2_lib.scala 243:37]
  wire  _T_738 = _T_737 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_741 = io_trigger_pkt_any_2_tdata2[21] == lsu_match_data_2[21]; // @[el2_lib.scala 243:79]
  wire  _T_742 = _T_738 | _T_741; // @[el2_lib.scala 243:24]
  wire  _T_744 = &io_trigger_pkt_any_2_tdata2[21:0]; // @[el2_lib.scala 243:37]
  wire  _T_745 = _T_744 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_748 = io_trigger_pkt_any_2_tdata2[22] == lsu_match_data_2[22]; // @[el2_lib.scala 243:79]
  wire  _T_749 = _T_745 | _T_748; // @[el2_lib.scala 243:24]
  wire  _T_751 = &io_trigger_pkt_any_2_tdata2[22:0]; // @[el2_lib.scala 243:37]
  wire  _T_752 = _T_751 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_755 = io_trigger_pkt_any_2_tdata2[23] == lsu_match_data_2[23]; // @[el2_lib.scala 243:79]
  wire  _T_756 = _T_752 | _T_755; // @[el2_lib.scala 243:24]
  wire  _T_758 = &io_trigger_pkt_any_2_tdata2[23:0]; // @[el2_lib.scala 243:37]
  wire  _T_759 = _T_758 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_762 = io_trigger_pkt_any_2_tdata2[24] == lsu_match_data_2[24]; // @[el2_lib.scala 243:79]
  wire  _T_763 = _T_759 | _T_762; // @[el2_lib.scala 243:24]
  wire  _T_765 = &io_trigger_pkt_any_2_tdata2[24:0]; // @[el2_lib.scala 243:37]
  wire  _T_766 = _T_765 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_769 = io_trigger_pkt_any_2_tdata2[25] == lsu_match_data_2[25]; // @[el2_lib.scala 243:79]
  wire  _T_770 = _T_766 | _T_769; // @[el2_lib.scala 243:24]
  wire  _T_772 = &io_trigger_pkt_any_2_tdata2[25:0]; // @[el2_lib.scala 243:37]
  wire  _T_773 = _T_772 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_776 = io_trigger_pkt_any_2_tdata2[26] == lsu_match_data_2[26]; // @[el2_lib.scala 243:79]
  wire  _T_777 = _T_773 | _T_776; // @[el2_lib.scala 243:24]
  wire  _T_779 = &io_trigger_pkt_any_2_tdata2[26:0]; // @[el2_lib.scala 243:37]
  wire  _T_780 = _T_779 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_783 = io_trigger_pkt_any_2_tdata2[27] == lsu_match_data_2[27]; // @[el2_lib.scala 243:79]
  wire  _T_784 = _T_780 | _T_783; // @[el2_lib.scala 243:24]
  wire  _T_786 = &io_trigger_pkt_any_2_tdata2[27:0]; // @[el2_lib.scala 243:37]
  wire  _T_787 = _T_786 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_790 = io_trigger_pkt_any_2_tdata2[28] == lsu_match_data_2[28]; // @[el2_lib.scala 243:79]
  wire  _T_791 = _T_787 | _T_790; // @[el2_lib.scala 243:24]
  wire  _T_793 = &io_trigger_pkt_any_2_tdata2[28:0]; // @[el2_lib.scala 243:37]
  wire  _T_794 = _T_793 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_797 = io_trigger_pkt_any_2_tdata2[29] == lsu_match_data_2[29]; // @[el2_lib.scala 243:79]
  wire  _T_798 = _T_794 | _T_797; // @[el2_lib.scala 243:24]
  wire  _T_800 = &io_trigger_pkt_any_2_tdata2[29:0]; // @[el2_lib.scala 243:37]
  wire  _T_801 = _T_800 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_804 = io_trigger_pkt_any_2_tdata2[30] == lsu_match_data_2[30]; // @[el2_lib.scala 243:79]
  wire  _T_805 = _T_801 | _T_804; // @[el2_lib.scala 243:24]
  wire  _T_807 = &io_trigger_pkt_any_2_tdata2[30:0]; // @[el2_lib.scala 243:37]
  wire  _T_808 = _T_807 & _T_591; // @[el2_lib.scala 243:42]
  wire  _T_811 = io_trigger_pkt_any_2_tdata2[31] == lsu_match_data_2[31]; // @[el2_lib.scala 243:79]
  wire  _T_812 = _T_808 | _T_811; // @[el2_lib.scala 243:24]
  wire [7:0] _T_819 = {_T_644,_T_637,_T_630,_T_623,_T_616,_T_609,_T_602,_T_595}; // @[el2_lib.scala 244:14]
  wire [15:0] _T_827 = {_T_700,_T_693,_T_686,_T_679,_T_672,_T_665,_T_658,_T_651,_T_819}; // @[el2_lib.scala 244:14]
  wire [7:0] _T_834 = {_T_756,_T_749,_T_742,_T_735,_T_728,_T_721,_T_714,_T_707}; // @[el2_lib.scala 244:14]
  wire [31:0] _T_843 = {_T_812,_T_805,_T_798,_T_791,_T_784,_T_777,_T_770,_T_763,_T_834,_T_827}; // @[el2_lib.scala 244:14]
  wire  _T_844 = &_T_843; // @[el2_lib.scala 244:21]
  wire  _T_845 = _T_584 & _T_844; // @[el2_lsu_trigger.scala 19:87]
  wire  _T_848 = io_trigger_pkt_any_3_store & io_lsu_pkt_m_store; // @[el2_lsu_trigger.scala 18:121]
  wire  _T_849 = io_trigger_pkt_any_3_load & io_lsu_pkt_m_load; // @[el2_lsu_trigger.scala 19:33]
  wire  _T_851 = _T_849 & _T_33; // @[el2_lsu_trigger.scala 19:53]
  wire  _T_852 = _T_848 | _T_851; // @[el2_lsu_trigger.scala 18:142]
  wire  _T_853 = _T_40 & _T_852; // @[el2_lsu_trigger.scala 18:89]
  wire  _T_858 = &io_trigger_pkt_any_3_tdata2; // @[el2_lib.scala 240:73]
  wire  _T_859 = ~_T_858; // @[el2_lib.scala 240:47]
  wire  _T_860 = io_trigger_pkt_any_3_match_ & _T_859; // @[el2_lib.scala 240:44]
  wire  _T_863 = io_trigger_pkt_any_3_tdata2[0] == lsu_match_data_3[0]; // @[el2_lib.scala 241:52]
  wire  _T_864 = _T_860 | _T_863; // @[el2_lib.scala 241:41]
  wire  _T_866 = &io_trigger_pkt_any_3_tdata2[0]; // @[el2_lib.scala 243:37]
  wire  _T_867 = _T_866 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_870 = io_trigger_pkt_any_3_tdata2[1] == lsu_match_data_3[1]; // @[el2_lib.scala 243:79]
  wire  _T_871 = _T_867 | _T_870; // @[el2_lib.scala 243:24]
  wire  _T_873 = &io_trigger_pkt_any_3_tdata2[1:0]; // @[el2_lib.scala 243:37]
  wire  _T_874 = _T_873 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_877 = io_trigger_pkt_any_3_tdata2[2] == lsu_match_data_3[2]; // @[el2_lib.scala 243:79]
  wire  _T_878 = _T_874 | _T_877; // @[el2_lib.scala 243:24]
  wire  _T_880 = &io_trigger_pkt_any_3_tdata2[2:0]; // @[el2_lib.scala 243:37]
  wire  _T_881 = _T_880 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_884 = io_trigger_pkt_any_3_tdata2[3] == lsu_match_data_3[3]; // @[el2_lib.scala 243:79]
  wire  _T_885 = _T_881 | _T_884; // @[el2_lib.scala 243:24]
  wire  _T_887 = &io_trigger_pkt_any_3_tdata2[3:0]; // @[el2_lib.scala 243:37]
  wire  _T_888 = _T_887 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_891 = io_trigger_pkt_any_3_tdata2[4] == lsu_match_data_3[4]; // @[el2_lib.scala 243:79]
  wire  _T_892 = _T_888 | _T_891; // @[el2_lib.scala 243:24]
  wire  _T_894 = &io_trigger_pkt_any_3_tdata2[4:0]; // @[el2_lib.scala 243:37]
  wire  _T_895 = _T_894 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_898 = io_trigger_pkt_any_3_tdata2[5] == lsu_match_data_3[5]; // @[el2_lib.scala 243:79]
  wire  _T_899 = _T_895 | _T_898; // @[el2_lib.scala 243:24]
  wire  _T_901 = &io_trigger_pkt_any_3_tdata2[5:0]; // @[el2_lib.scala 243:37]
  wire  _T_902 = _T_901 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_905 = io_trigger_pkt_any_3_tdata2[6] == lsu_match_data_3[6]; // @[el2_lib.scala 243:79]
  wire  _T_906 = _T_902 | _T_905; // @[el2_lib.scala 243:24]
  wire  _T_908 = &io_trigger_pkt_any_3_tdata2[6:0]; // @[el2_lib.scala 243:37]
  wire  _T_909 = _T_908 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_912 = io_trigger_pkt_any_3_tdata2[7] == lsu_match_data_3[7]; // @[el2_lib.scala 243:79]
  wire  _T_913 = _T_909 | _T_912; // @[el2_lib.scala 243:24]
  wire  _T_915 = &io_trigger_pkt_any_3_tdata2[7:0]; // @[el2_lib.scala 243:37]
  wire  _T_916 = _T_915 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_919 = io_trigger_pkt_any_3_tdata2[8] == lsu_match_data_3[8]; // @[el2_lib.scala 243:79]
  wire  _T_920 = _T_916 | _T_919; // @[el2_lib.scala 243:24]
  wire  _T_922 = &io_trigger_pkt_any_3_tdata2[8:0]; // @[el2_lib.scala 243:37]
  wire  _T_923 = _T_922 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_926 = io_trigger_pkt_any_3_tdata2[9] == lsu_match_data_3[9]; // @[el2_lib.scala 243:79]
  wire  _T_927 = _T_923 | _T_926; // @[el2_lib.scala 243:24]
  wire  _T_929 = &io_trigger_pkt_any_3_tdata2[9:0]; // @[el2_lib.scala 243:37]
  wire  _T_930 = _T_929 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_933 = io_trigger_pkt_any_3_tdata2[10] == lsu_match_data_3[10]; // @[el2_lib.scala 243:79]
  wire  _T_934 = _T_930 | _T_933; // @[el2_lib.scala 243:24]
  wire  _T_936 = &io_trigger_pkt_any_3_tdata2[10:0]; // @[el2_lib.scala 243:37]
  wire  _T_937 = _T_936 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_940 = io_trigger_pkt_any_3_tdata2[11] == lsu_match_data_3[11]; // @[el2_lib.scala 243:79]
  wire  _T_941 = _T_937 | _T_940; // @[el2_lib.scala 243:24]
  wire  _T_943 = &io_trigger_pkt_any_3_tdata2[11:0]; // @[el2_lib.scala 243:37]
  wire  _T_944 = _T_943 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_947 = io_trigger_pkt_any_3_tdata2[12] == lsu_match_data_3[12]; // @[el2_lib.scala 243:79]
  wire  _T_948 = _T_944 | _T_947; // @[el2_lib.scala 243:24]
  wire  _T_950 = &io_trigger_pkt_any_3_tdata2[12:0]; // @[el2_lib.scala 243:37]
  wire  _T_951 = _T_950 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_954 = io_trigger_pkt_any_3_tdata2[13] == lsu_match_data_3[13]; // @[el2_lib.scala 243:79]
  wire  _T_955 = _T_951 | _T_954; // @[el2_lib.scala 243:24]
  wire  _T_957 = &io_trigger_pkt_any_3_tdata2[13:0]; // @[el2_lib.scala 243:37]
  wire  _T_958 = _T_957 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_961 = io_trigger_pkt_any_3_tdata2[14] == lsu_match_data_3[14]; // @[el2_lib.scala 243:79]
  wire  _T_962 = _T_958 | _T_961; // @[el2_lib.scala 243:24]
  wire  _T_964 = &io_trigger_pkt_any_3_tdata2[14:0]; // @[el2_lib.scala 243:37]
  wire  _T_965 = _T_964 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_968 = io_trigger_pkt_any_3_tdata2[15] == lsu_match_data_3[15]; // @[el2_lib.scala 243:79]
  wire  _T_969 = _T_965 | _T_968; // @[el2_lib.scala 243:24]
  wire  _T_971 = &io_trigger_pkt_any_3_tdata2[15:0]; // @[el2_lib.scala 243:37]
  wire  _T_972 = _T_971 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_975 = io_trigger_pkt_any_3_tdata2[16] == lsu_match_data_3[16]; // @[el2_lib.scala 243:79]
  wire  _T_976 = _T_972 | _T_975; // @[el2_lib.scala 243:24]
  wire  _T_978 = &io_trigger_pkt_any_3_tdata2[16:0]; // @[el2_lib.scala 243:37]
  wire  _T_979 = _T_978 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_982 = io_trigger_pkt_any_3_tdata2[17] == lsu_match_data_3[17]; // @[el2_lib.scala 243:79]
  wire  _T_983 = _T_979 | _T_982; // @[el2_lib.scala 243:24]
  wire  _T_985 = &io_trigger_pkt_any_3_tdata2[17:0]; // @[el2_lib.scala 243:37]
  wire  _T_986 = _T_985 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_989 = io_trigger_pkt_any_3_tdata2[18] == lsu_match_data_3[18]; // @[el2_lib.scala 243:79]
  wire  _T_990 = _T_986 | _T_989; // @[el2_lib.scala 243:24]
  wire  _T_992 = &io_trigger_pkt_any_3_tdata2[18:0]; // @[el2_lib.scala 243:37]
  wire  _T_993 = _T_992 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_996 = io_trigger_pkt_any_3_tdata2[19] == lsu_match_data_3[19]; // @[el2_lib.scala 243:79]
  wire  _T_997 = _T_993 | _T_996; // @[el2_lib.scala 243:24]
  wire  _T_999 = &io_trigger_pkt_any_3_tdata2[19:0]; // @[el2_lib.scala 243:37]
  wire  _T_1000 = _T_999 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1003 = io_trigger_pkt_any_3_tdata2[20] == lsu_match_data_3[20]; // @[el2_lib.scala 243:79]
  wire  _T_1004 = _T_1000 | _T_1003; // @[el2_lib.scala 243:24]
  wire  _T_1006 = &io_trigger_pkt_any_3_tdata2[20:0]; // @[el2_lib.scala 243:37]
  wire  _T_1007 = _T_1006 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1010 = io_trigger_pkt_any_3_tdata2[21] == lsu_match_data_3[21]; // @[el2_lib.scala 243:79]
  wire  _T_1011 = _T_1007 | _T_1010; // @[el2_lib.scala 243:24]
  wire  _T_1013 = &io_trigger_pkt_any_3_tdata2[21:0]; // @[el2_lib.scala 243:37]
  wire  _T_1014 = _T_1013 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1017 = io_trigger_pkt_any_3_tdata2[22] == lsu_match_data_3[22]; // @[el2_lib.scala 243:79]
  wire  _T_1018 = _T_1014 | _T_1017; // @[el2_lib.scala 243:24]
  wire  _T_1020 = &io_trigger_pkt_any_3_tdata2[22:0]; // @[el2_lib.scala 243:37]
  wire  _T_1021 = _T_1020 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1024 = io_trigger_pkt_any_3_tdata2[23] == lsu_match_data_3[23]; // @[el2_lib.scala 243:79]
  wire  _T_1025 = _T_1021 | _T_1024; // @[el2_lib.scala 243:24]
  wire  _T_1027 = &io_trigger_pkt_any_3_tdata2[23:0]; // @[el2_lib.scala 243:37]
  wire  _T_1028 = _T_1027 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1031 = io_trigger_pkt_any_3_tdata2[24] == lsu_match_data_3[24]; // @[el2_lib.scala 243:79]
  wire  _T_1032 = _T_1028 | _T_1031; // @[el2_lib.scala 243:24]
  wire  _T_1034 = &io_trigger_pkt_any_3_tdata2[24:0]; // @[el2_lib.scala 243:37]
  wire  _T_1035 = _T_1034 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1038 = io_trigger_pkt_any_3_tdata2[25] == lsu_match_data_3[25]; // @[el2_lib.scala 243:79]
  wire  _T_1039 = _T_1035 | _T_1038; // @[el2_lib.scala 243:24]
  wire  _T_1041 = &io_trigger_pkt_any_3_tdata2[25:0]; // @[el2_lib.scala 243:37]
  wire  _T_1042 = _T_1041 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1045 = io_trigger_pkt_any_3_tdata2[26] == lsu_match_data_3[26]; // @[el2_lib.scala 243:79]
  wire  _T_1046 = _T_1042 | _T_1045; // @[el2_lib.scala 243:24]
  wire  _T_1048 = &io_trigger_pkt_any_3_tdata2[26:0]; // @[el2_lib.scala 243:37]
  wire  _T_1049 = _T_1048 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1052 = io_trigger_pkt_any_3_tdata2[27] == lsu_match_data_3[27]; // @[el2_lib.scala 243:79]
  wire  _T_1053 = _T_1049 | _T_1052; // @[el2_lib.scala 243:24]
  wire  _T_1055 = &io_trigger_pkt_any_3_tdata2[27:0]; // @[el2_lib.scala 243:37]
  wire  _T_1056 = _T_1055 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1059 = io_trigger_pkt_any_3_tdata2[28] == lsu_match_data_3[28]; // @[el2_lib.scala 243:79]
  wire  _T_1060 = _T_1056 | _T_1059; // @[el2_lib.scala 243:24]
  wire  _T_1062 = &io_trigger_pkt_any_3_tdata2[28:0]; // @[el2_lib.scala 243:37]
  wire  _T_1063 = _T_1062 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1066 = io_trigger_pkt_any_3_tdata2[29] == lsu_match_data_3[29]; // @[el2_lib.scala 243:79]
  wire  _T_1067 = _T_1063 | _T_1066; // @[el2_lib.scala 243:24]
  wire  _T_1069 = &io_trigger_pkt_any_3_tdata2[29:0]; // @[el2_lib.scala 243:37]
  wire  _T_1070 = _T_1069 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1073 = io_trigger_pkt_any_3_tdata2[30] == lsu_match_data_3[30]; // @[el2_lib.scala 243:79]
  wire  _T_1074 = _T_1070 | _T_1073; // @[el2_lib.scala 243:24]
  wire  _T_1076 = &io_trigger_pkt_any_3_tdata2[30:0]; // @[el2_lib.scala 243:37]
  wire  _T_1077 = _T_1076 & _T_860; // @[el2_lib.scala 243:42]
  wire  _T_1080 = io_trigger_pkt_any_3_tdata2[31] == lsu_match_data_3[31]; // @[el2_lib.scala 243:79]
  wire  _T_1081 = _T_1077 | _T_1080; // @[el2_lib.scala 243:24]
  wire [7:0] _T_1088 = {_T_913,_T_906,_T_899,_T_892,_T_885,_T_878,_T_871,_T_864}; // @[el2_lib.scala 244:14]
  wire [15:0] _T_1096 = {_T_969,_T_962,_T_955,_T_948,_T_941,_T_934,_T_927,_T_920,_T_1088}; // @[el2_lib.scala 244:14]
  wire [7:0] _T_1103 = {_T_1025,_T_1018,_T_1011,_T_1004,_T_997,_T_990,_T_983,_T_976}; // @[el2_lib.scala 244:14]
  wire [31:0] _T_1112 = {_T_1081,_T_1074,_T_1067,_T_1060,_T_1053,_T_1046,_T_1039,_T_1032,_T_1103,_T_1096}; // @[el2_lib.scala 244:14]
  wire  _T_1113 = &_T_1112; // @[el2_lib.scala 244:21]
  wire  _T_1114 = _T_853 & _T_1113; // @[el2_lsu_trigger.scala 19:87]
  wire [2:0] _T_1116 = {_T_1114,_T_845,_T_576}; // @[Cat.scala 29:58]
  assign io_lsu_trigger_match_m = {_T_1116,_T_307}; // @[el2_lsu_trigger.scala 18:26]
endmodule
