module RVCExpander(
  input         clock,
  input         reset,
  input  [31:0] io_in,
  output [31:0] io_out_bits,
  output [4:0]  io_out_rd,
  output [4:0]  io_out_rs1,
  output [4:0]  io_out_rs2,
  output [4:0]  io_out_rs3,
  output        io_rvc
);
  wire  _T_3 = |io_in[12:5]; // @[el2_ifu_compress.scala 49:29]
  wire [6:0] _T_4 = _T_3 ? 7'h13 : 7'h1f; // @[el2_ifu_compress.scala 49:20]
  wire [4:0] _T_14 = {2'h1,io_in[4:2]}; // @[Cat.scala 29:58]
  wire [29:0] _T_18 = {io_in[10:7],io_in[12:11],io_in[5],io_in[6],2'h0,5'h2,3'h0,2'h1,io_in[4:2],_T_4}; // @[Cat.scala 29:58]
  wire [7:0] _T_28 = {io_in[6:5],io_in[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [4:0] _T_30 = {2'h1,io_in[9:7]}; // @[Cat.scala 29:58]
  wire [27:0] _T_36 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h7}; // @[Cat.scala 29:58]
  wire [6:0] _T_50 = {io_in[5],io_in[12:10],io_in[6],2'h0}; // @[Cat.scala 29:58]
  wire [26:0] _T_58 = {io_in[5],io_in[12:10],io_in[6],2'h0,2'h1,io_in[9:7],3'h2,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [27:0] _T_78 = {io_in[6:5],io_in[12:10],3'h0,2'h1,io_in[9:7],3'h3,2'h1,io_in[4:2],7'h3}; // @[Cat.scala 29:58]
  wire [26:0] _T_109 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h3f}; // @[Cat.scala 29:58]
  wire [27:0] _T_136 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [26:0] _T_167 = {_T_50[6:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h2,_T_50[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [27:0] _T_194 = {_T_28[7:5],2'h1,io_in[4:2],2'h1,io_in[9:7],3'h3,_T_28[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [6:0] _T_205 = io_in[12] ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12]
  wire [11:0] _T_207 = {_T_205,io_in[6:2]}; // @[Cat.scala 29:58]
  wire [31:0] _T_213 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_221 = |io_in[11:7]; // @[el2_ifu_compress.scala 73:24]
  wire [6:0] _T_222 = _T_221 ? 7'h1b : 7'h1f; // @[el2_ifu_compress.scala 73:20]
  wire [31:0] _T_233 = {_T_205,io_in[6:2],io_in[11:7],3'h0,io_in[11:7],_T_222}; // @[Cat.scala 29:58]
  wire [31:0] _T_249 = {_T_205,io_in[6:2],5'h0,3'h0,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  wire  _T_260 = |_T_207; // @[el2_ifu_compress.scala 86:29]
  wire [6:0] _T_261 = _T_260 ? 7'h37 : 7'h3f; // @[el2_ifu_compress.scala 86:20]
  wire [14:0] _T_264 = io_in[12] ? 15'h7fff : 15'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_267 = {_T_264,io_in[6:2],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_271 = {_T_267[31:12],io_in[11:7],_T_261}; // @[Cat.scala 29:58]
  wire  _T_279 = io_in[11:7] == 5'h0; // @[el2_ifu_compress.scala 88:14]
  wire  _T_281 = io_in[11:7] == 5'h2; // @[el2_ifu_compress.scala 88:27]
  wire  _T_282 = _T_279 | _T_281; // @[el2_ifu_compress.scala 88:21]
  wire [6:0] _T_289 = _T_260 ? 7'h13 : 7'h1f; // @[el2_ifu_compress.scala 82:20]
  wire [2:0] _T_292 = io_in[12] ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_307 = {_T_292,io_in[4:3],io_in[5],io_in[2],io_in[6],4'h0,io_in[11:7],3'h0,io_in[11:7],_T_289}; // @[Cat.scala 29:58]
  wire [31:0] _T_314_bits = _T_282 ? _T_307 : _T_271; // @[el2_ifu_compress.scala 88:10]
  wire [4:0] _T_314_rd = _T_282 ? io_in[11:7] : io_in[11:7]; // @[el2_ifu_compress.scala 88:10]
  wire [4:0] _T_314_rs2 = _T_282 ? _T_14 : _T_14; // @[el2_ifu_compress.scala 88:10]
  wire [4:0] _T_314_rs3 = _T_282 ? io_in[31:27] : io_in[31:27]; // @[el2_ifu_compress.scala 88:10]
  wire [25:0] _T_325 = {io_in[12],io_in[6:2],2'h1,io_in[9:7],3'h5,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_172 = {{5'd0}, _T_325}; // @[el2_ifu_compress.scala 95:23]
  wire [30:0] _T_337 = _GEN_172 | 31'h40000000; // @[el2_ifu_compress.scala 95:23]
  wire [31:0] _T_350 = {_T_205,io_in[6:2],2'h1,io_in[9:7],3'h7,2'h1,io_in[9:7],7'h13}; // @[Cat.scala 29:58]
  wire [2:0] _T_354 = {io_in[12],io_in[6:5]}; // @[Cat.scala 29:58]
  wire  _T_356 = io_in[6:5] == 2'h0; // @[el2_ifu_compress.scala 99:30]
  wire [30:0] _T_357 = _T_356 ? 31'h40000000 : 31'h0; // @[el2_ifu_compress.scala 99:22]
  wire [6:0] _T_359 = io_in[12] ? 7'h3b : 7'h33; // @[el2_ifu_compress.scala 100:22]
  wire [2:0] _GEN_1 = 3'h1 == _T_354 ? 3'h4 : 3'h0; // @[Cat.scala 29:58]
  wire [2:0] _GEN_2 = 3'h2 == _T_354 ? 3'h6 : _GEN_1; // @[Cat.scala 29:58]
  wire [2:0] _GEN_3 = 3'h3 == _T_354 ? 3'h7 : _GEN_2; // @[Cat.scala 29:58]
  wire [2:0] _GEN_4 = 3'h4 == _T_354 ? 3'h0 : _GEN_3; // @[Cat.scala 29:58]
  wire [2:0] _GEN_5 = 3'h5 == _T_354 ? 3'h0 : _GEN_4; // @[Cat.scala 29:58]
  wire [2:0] _GEN_6 = 3'h6 == _T_354 ? 3'h2 : _GEN_5; // @[Cat.scala 29:58]
  wire [2:0] _GEN_7 = 3'h7 == _T_354 ? 3'h3 : _GEN_6; // @[Cat.scala 29:58]
  wire [24:0] _T_369 = {2'h1,io_in[4:2],2'h1,io_in[9:7],_GEN_7,2'h1,io_in[9:7],_T_359}; // @[Cat.scala 29:58]
  wire [30:0] _GEN_173 = {{6'd0}, _T_369}; // @[el2_ifu_compress.scala 101:43]
  wire [30:0] _T_370 = _GEN_173 | _T_357; // @[el2_ifu_compress.scala 101:43]
  wire [31:0] _T_371_0 = {{6'd0}, _T_325}; // @[el2_ifu_compress.scala 103:19 el2_ifu_compress.scala 103:19]
  wire [31:0] _T_371_1 = {{1'd0}, _T_337}; // @[el2_ifu_compress.scala 103:19 el2_ifu_compress.scala 103:19]
  wire [31:0] _GEN_9 = 2'h1 == io_in[11:10] ? _T_371_1 : _T_371_0; // @[el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_10 = 2'h2 == io_in[11:10] ? _T_350 : _GEN_9; // @[el2_ifu_compress.scala 18:14]
  wire [31:0] _T_371_3 = {{1'd0}, _T_370}; // @[el2_ifu_compress.scala 103:19 el2_ifu_compress.scala 103:19]
  wire [31:0] _GEN_11 = 2'h3 == io_in[11:10] ? _T_371_3 : _GEN_10; // @[el2_ifu_compress.scala 18:14]
  wire [9:0] _T_383 = io_in[12] ? 10'h3ff : 10'h0; // @[Bitwise.scala 72:12]
  wire [20:0] _T_398 = {_T_383,io_in[8],io_in[10:9],io_in[6],io_in[7],io_in[2],io_in[11],io_in[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_461 = {_T_398[20],_T_398[10:1],_T_398[11],_T_398[19:12],5'h0,7'h6f}; // @[Cat.scala 29:58]
  wire [4:0] _T_470 = io_in[12] ? 5'h1f : 5'h0; // @[Bitwise.scala 72:12]
  wire [12:0] _T_479 = {_T_470,io_in[6:5],io_in[2],io_in[11:10],io_in[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_528 = {_T_479[12],_T_479[10:5],5'h0,2'h1,io_in[9:7],3'h0,_T_479[4:1],_T_479[11],7'h63}; // @[Cat.scala 29:58]
  wire [31:0] _T_595 = {_T_479[12],_T_479[10:5],5'h0,2'h1,io_in[9:7],3'h1,_T_479[4:1],_T_479[11],7'h63}; // @[Cat.scala 29:58]
  wire [6:0] _T_602 = _T_221 ? 7'h3 : 7'h1f; // @[el2_ifu_compress.scala 109:23]
  wire [25:0] _T_611 = {io_in[12],io_in[6:2],io_in[11:7],3'h1,io_in[11:7],7'h13}; // @[Cat.scala 29:58]
  wire [28:0] _T_627 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],7'h7}; // @[Cat.scala 29:58]
  wire [27:0] _T_642 = {io_in[3:2],io_in[12],io_in[6:4],2'h0,5'h2,3'h2,io_in[11:7],_T_602}; // @[Cat.scala 29:58]
  wire [28:0] _T_657 = {io_in[4:2],io_in[12],io_in[6:5],3'h0,5'h2,3'h3,io_in[11:7],_T_602}; // @[Cat.scala 29:58]
  wire [24:0] _T_667 = {io_in[6:2],5'h0,3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_678 = {io_in[6:2],io_in[11:7],3'h0,io_in[11:7],7'h33}; // @[Cat.scala 29:58]
  wire [24:0] _T_689 = {io_in[6:2],io_in[11:7],3'h0,12'h67}; // @[Cat.scala 29:58]
  wire [24:0] _T_691 = {_T_689[24:7],7'h1f}; // @[Cat.scala 29:58]
  wire [24:0] _T_694 = _T_221 ? _T_689 : _T_691; // @[el2_ifu_compress.scala 130:33]
  wire  _T_700 = |io_in[6:2]; // @[el2_ifu_compress.scala 131:27]
  wire [31:0] _T_671_bits = {{7'd0}, _T_667}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _T_698_bits = {{7'd0}, _T_694}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _T_701_bits = _T_700 ? _T_671_bits : _T_698_bits; // @[el2_ifu_compress.scala 131:22]
  wire [4:0] _T_701_rd = _T_700 ? io_in[11:7] : 5'h0; // @[el2_ifu_compress.scala 131:22]
  wire [4:0] _T_701_rs1 = _T_700 ? 5'h0 : io_in[11:7]; // @[el2_ifu_compress.scala 131:22]
  wire [4:0] _T_701_rs2 = _T_700 ? io_in[6:2] : io_in[6:2]; // @[el2_ifu_compress.scala 131:22]
  wire [4:0] _T_701_rs3 = _T_700 ? io_in[31:27] : io_in[31:27]; // @[el2_ifu_compress.scala 131:22]
  wire [24:0] _T_707 = {io_in[6:2],io_in[11:7],3'h0,12'he7}; // @[Cat.scala 29:58]
  wire [24:0] _T_709 = {_T_689[24:7],7'h73}; // @[Cat.scala 29:58]
  wire [24:0] _T_710 = _T_709 | 25'h100000; // @[el2_ifu_compress.scala 133:46]
  wire [24:0] _T_713 = _T_221 ? _T_707 : _T_710; // @[el2_ifu_compress.scala 134:33]
  wire [31:0] _T_683_bits = {{7'd0}, _T_678}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _T_717_bits = {{7'd0}, _T_713}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _T_720_bits = _T_700 ? _T_683_bits : _T_717_bits; // @[el2_ifu_compress.scala 135:25]
  wire [4:0] _T_720_rd = _T_700 ? io_in[11:7] : 5'h1; // @[el2_ifu_compress.scala 135:25]
  wire [4:0] _T_720_rs1 = _T_700 ? io_in[11:7] : io_in[11:7]; // @[el2_ifu_compress.scala 135:25]
  wire [31:0] _T_722_bits = io_in[12] ? _T_720_bits : _T_701_bits; // @[el2_ifu_compress.scala 136:10]
  wire [4:0] _T_722_rd = io_in[12] ? _T_720_rd : _T_701_rd; // @[el2_ifu_compress.scala 136:10]
  wire [4:0] _T_722_rs1 = io_in[12] ? _T_720_rs1 : _T_701_rs1; // @[el2_ifu_compress.scala 136:10]
  wire [4:0] _T_722_rs2 = io_in[12] ? _T_701_rs2 : _T_701_rs2; // @[el2_ifu_compress.scala 136:10]
  wire [4:0] _T_722_rs3 = io_in[12] ? _T_701_rs3 : _T_701_rs3; // @[el2_ifu_compress.scala 136:10]
  wire [8:0] _T_726 = {io_in[9:7],io_in[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [28:0] _T_738 = {_T_726[8:5],io_in[6:2],5'h2,3'h3,_T_726[4:0],7'h27}; // @[Cat.scala 29:58]
  wire [7:0] _T_746 = {io_in[8:7],io_in[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [27:0] _T_758 = {_T_746[7:5],io_in[6:2],5'h2,3'h2,_T_746[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [28:0] _T_778 = {_T_726[8:5],io_in[6:2],5'h2,3'h3,_T_726[4:0],7'h23}; // @[Cat.scala 29:58]
  wire [4:0] _T_826 = {io_in[1:0],io_in[15:13]}; // @[Cat.scala 29:58]
  wire [31:0] _T_24_bits = {{2'd0}, _T_18}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _T_44_bits = {{4'd0}, _T_36}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_17 = 5'h1 == _T_826 ? _T_44_bits : _T_24_bits; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_18 = 5'h1 == _T_826 ? _T_14 : _T_14; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_19 = 5'h1 == _T_826 ? _T_30 : 5'h2; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_21 = 5'h1 == _T_826 ? io_in[31:27] : io_in[31:27]; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_66_bits = {{5'd0}, _T_58}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_22 = 5'h2 == _T_826 ? _T_66_bits : _GEN_17; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_23 = 5'h2 == _T_826 ? _T_14 : _GEN_18; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_24 = 5'h2 == _T_826 ? _T_30 : _GEN_19; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_26 = 5'h2 == _T_826 ? io_in[31:27] : _GEN_21; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_86_bits = {{4'd0}, _T_78}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_27 = 5'h3 == _T_826 ? _T_86_bits : _GEN_22; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_28 = 5'h3 == _T_826 ? _T_14 : _GEN_23; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_29 = 5'h3 == _T_826 ? _T_30 : _GEN_24; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_31 = 5'h3 == _T_826 ? io_in[31:27] : _GEN_26; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_117_bits = {{5'd0}, _T_109}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_32 = 5'h4 == _T_826 ? _T_117_bits : _GEN_27; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_33 = 5'h4 == _T_826 ? _T_14 : _GEN_28; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_34 = 5'h4 == _T_826 ? _T_30 : _GEN_29; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_36 = 5'h4 == _T_826 ? io_in[31:27] : _GEN_31; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_144_bits = {{4'd0}, _T_136}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_37 = 5'h5 == _T_826 ? _T_144_bits : _GEN_32; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_38 = 5'h5 == _T_826 ? _T_14 : _GEN_33; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_39 = 5'h5 == _T_826 ? _T_30 : _GEN_34; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_41 = 5'h5 == _T_826 ? io_in[31:27] : _GEN_36; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_175_bits = {{5'd0}, _T_167}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_42 = 5'h6 == _T_826 ? _T_175_bits : _GEN_37; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_43 = 5'h6 == _T_826 ? _T_14 : _GEN_38; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_44 = 5'h6 == _T_826 ? _T_30 : _GEN_39; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_46 = 5'h6 == _T_826 ? io_in[31:27] : _GEN_41; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_202_bits = {{4'd0}, _T_194}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_47 = 5'h7 == _T_826 ? _T_202_bits : _GEN_42; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_48 = 5'h7 == _T_826 ? _T_14 : _GEN_43; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_49 = 5'h7 == _T_826 ? _T_30 : _GEN_44; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_51 = 5'h7 == _T_826 ? io_in[31:27] : _GEN_46; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_52 = 5'h8 == _T_826 ? _T_213 : _GEN_47; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_53 = 5'h8 == _T_826 ? io_in[11:7] : _GEN_48; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_54 = 5'h8 == _T_826 ? io_in[11:7] : _GEN_49; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_55 = 5'h8 == _T_826 ? _T_14 : _GEN_48; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_56 = 5'h8 == _T_826 ? io_in[31:27] : _GEN_51; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_57 = 5'h9 == _T_826 ? _T_233 : _GEN_52; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_58 = 5'h9 == _T_826 ? io_in[11:7] : _GEN_53; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_59 = 5'h9 == _T_826 ? io_in[11:7] : _GEN_54; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_60 = 5'h9 == _T_826 ? _T_14 : _GEN_55; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_61 = 5'h9 == _T_826 ? io_in[31:27] : _GEN_56; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_62 = 5'ha == _T_826 ? _T_249 : _GEN_57; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_63 = 5'ha == _T_826 ? io_in[11:7] : _GEN_58; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_64 = 5'ha == _T_826 ? 5'h0 : _GEN_59; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_65 = 5'ha == _T_826 ? _T_14 : _GEN_60; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_66 = 5'ha == _T_826 ? io_in[31:27] : _GEN_61; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_67 = 5'hb == _T_826 ? _T_314_bits : _GEN_62; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_68 = 5'hb == _T_826 ? _T_314_rd : _GEN_63; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_69 = 5'hb == _T_826 ? _T_314_rd : _GEN_64; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_70 = 5'hb == _T_826 ? _T_314_rs2 : _GEN_65; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_71 = 5'hb == _T_826 ? _T_314_rs3 : _GEN_66; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_72 = 5'hc == _T_826 ? _GEN_11 : _GEN_67; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_73 = 5'hc == _T_826 ? _T_30 : _GEN_68; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_74 = 5'hc == _T_826 ? _T_30 : _GEN_69; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_75 = 5'hc == _T_826 ? _T_14 : _GEN_70; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_76 = 5'hc == _T_826 ? io_in[31:27] : _GEN_71; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_77 = 5'hd == _T_826 ? _T_461 : _GEN_72; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_78 = 5'hd == _T_826 ? 5'h0 : _GEN_73; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_79 = 5'hd == _T_826 ? _T_30 : _GEN_74; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_80 = 5'hd == _T_826 ? _T_14 : _GEN_75; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_81 = 5'hd == _T_826 ? io_in[31:27] : _GEN_76; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_82 = 5'he == _T_826 ? _T_528 : _GEN_77; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_83 = 5'he == _T_826 ? _T_30 : _GEN_78; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_84 = 5'he == _T_826 ? _T_30 : _GEN_79; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_85 = 5'he == _T_826 ? 5'h0 : _GEN_80; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_86 = 5'he == _T_826 ? io_in[31:27] : _GEN_81; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_87 = 5'hf == _T_826 ? _T_595 : _GEN_82; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_88 = 5'hf == _T_826 ? 5'h0 : _GEN_83; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_89 = 5'hf == _T_826 ? _T_30 : _GEN_84; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_90 = 5'hf == _T_826 ? 5'h0 : _GEN_85; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_91 = 5'hf == _T_826 ? io_in[31:27] : _GEN_86; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_616_bits = {{6'd0}, _T_611}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_92 = 5'h10 == _T_826 ? _T_616_bits : _GEN_87; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_93 = 5'h10 == _T_826 ? io_in[11:7] : _GEN_88; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_94 = 5'h10 == _T_826 ? io_in[11:7] : _GEN_89; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_95 = 5'h10 == _T_826 ? io_in[6:2] : _GEN_90; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_96 = 5'h10 == _T_826 ? io_in[31:27] : _GEN_91; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_631_bits = {{3'd0}, _T_627}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_97 = 5'h11 == _T_826 ? _T_631_bits : _GEN_92; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_98 = 5'h11 == _T_826 ? io_in[11:7] : _GEN_93; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_99 = 5'h11 == _T_826 ? 5'h2 : _GEN_94; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_100 = 5'h11 == _T_826 ? io_in[6:2] : _GEN_95; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_101 = 5'h11 == _T_826 ? io_in[31:27] : _GEN_96; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_646_bits = {{4'd0}, _T_642}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_102 = 5'h12 == _T_826 ? _T_646_bits : _GEN_97; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_103 = 5'h12 == _T_826 ? io_in[11:7] : _GEN_98; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_104 = 5'h12 == _T_826 ? 5'h2 : _GEN_99; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_105 = 5'h12 == _T_826 ? io_in[6:2] : _GEN_100; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_106 = 5'h12 == _T_826 ? io_in[31:27] : _GEN_101; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_661_bits = {{3'd0}, _T_657}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_107 = 5'h13 == _T_826 ? _T_661_bits : _GEN_102; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_108 = 5'h13 == _T_826 ? io_in[11:7] : _GEN_103; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_109 = 5'h13 == _T_826 ? 5'h2 : _GEN_104; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_110 = 5'h13 == _T_826 ? io_in[6:2] : _GEN_105; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_111 = 5'h13 == _T_826 ? io_in[31:27] : _GEN_106; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_112 = 5'h14 == _T_826 ? _T_722_bits : _GEN_107; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_113 = 5'h14 == _T_826 ? _T_722_rd : _GEN_108; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_114 = 5'h14 == _T_826 ? _T_722_rs1 : _GEN_109; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_115 = 5'h14 == _T_826 ? _T_722_rs2 : _GEN_110; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_116 = 5'h14 == _T_826 ? _T_722_rs3 : _GEN_111; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_742_bits = {{3'd0}, _T_738}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_117 = 5'h15 == _T_826 ? _T_742_bits : _GEN_112; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_118 = 5'h15 == _T_826 ? io_in[11:7] : _GEN_113; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_119 = 5'h15 == _T_826 ? 5'h2 : _GEN_114; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_120 = 5'h15 == _T_826 ? io_in[6:2] : _GEN_115; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_121 = 5'h15 == _T_826 ? io_in[31:27] : _GEN_116; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_762_bits = {{4'd0}, _T_758}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_122 = 5'h16 == _T_826 ? _T_762_bits : _GEN_117; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_123 = 5'h16 == _T_826 ? io_in[11:7] : _GEN_118; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_124 = 5'h16 == _T_826 ? 5'h2 : _GEN_119; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_125 = 5'h16 == _T_826 ? io_in[6:2] : _GEN_120; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_126 = 5'h16 == _T_826 ? io_in[31:27] : _GEN_121; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _T_782_bits = {{3'd0}, _T_778}; // @[el2_ifu_compress.scala 17:19 el2_ifu_compress.scala 18:14]
  wire [31:0] _GEN_127 = 5'h17 == _T_826 ? _T_782_bits : _GEN_122; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_128 = 5'h17 == _T_826 ? io_in[11:7] : _GEN_123; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_129 = 5'h17 == _T_826 ? 5'h2 : _GEN_124; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_130 = 5'h17 == _T_826 ? io_in[6:2] : _GEN_125; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_131 = 5'h17 == _T_826 ? io_in[31:27] : _GEN_126; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_132 = 5'h18 == _T_826 ? io_in : _GEN_127; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_133 = 5'h18 == _T_826 ? io_in[11:7] : _GEN_128; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_134 = 5'h18 == _T_826 ? io_in[19:15] : _GEN_129; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_135 = 5'h18 == _T_826 ? io_in[24:20] : _GEN_130; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_136 = 5'h18 == _T_826 ? io_in[31:27] : _GEN_131; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_137 = 5'h19 == _T_826 ? io_in : _GEN_132; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_138 = 5'h19 == _T_826 ? io_in[11:7] : _GEN_133; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_139 = 5'h19 == _T_826 ? io_in[19:15] : _GEN_134; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_140 = 5'h19 == _T_826 ? io_in[24:20] : _GEN_135; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_141 = 5'h19 == _T_826 ? io_in[31:27] : _GEN_136; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_142 = 5'h1a == _T_826 ? io_in : _GEN_137; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_143 = 5'h1a == _T_826 ? io_in[11:7] : _GEN_138; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_144 = 5'h1a == _T_826 ? io_in[19:15] : _GEN_139; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_145 = 5'h1a == _T_826 ? io_in[24:20] : _GEN_140; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_146 = 5'h1a == _T_826 ? io_in[31:27] : _GEN_141; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_147 = 5'h1b == _T_826 ? io_in : _GEN_142; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_148 = 5'h1b == _T_826 ? io_in[11:7] : _GEN_143; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_149 = 5'h1b == _T_826 ? io_in[19:15] : _GEN_144; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_150 = 5'h1b == _T_826 ? io_in[24:20] : _GEN_145; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_151 = 5'h1b == _T_826 ? io_in[31:27] : _GEN_146; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_152 = 5'h1c == _T_826 ? io_in : _GEN_147; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_153 = 5'h1c == _T_826 ? io_in[11:7] : _GEN_148; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_154 = 5'h1c == _T_826 ? io_in[19:15] : _GEN_149; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_155 = 5'h1c == _T_826 ? io_in[24:20] : _GEN_150; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_156 = 5'h1c == _T_826 ? io_in[31:27] : _GEN_151; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_157 = 5'h1d == _T_826 ? io_in : _GEN_152; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_158 = 5'h1d == _T_826 ? io_in[11:7] : _GEN_153; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_159 = 5'h1d == _T_826 ? io_in[19:15] : _GEN_154; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_160 = 5'h1d == _T_826 ? io_in[24:20] : _GEN_155; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_161 = 5'h1d == _T_826 ? io_in[31:27] : _GEN_156; // @[el2_ifu_compress.scala 195:12]
  wire [31:0] _GEN_162 = 5'h1e == _T_826 ? io_in : _GEN_157; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_163 = 5'h1e == _T_826 ? io_in[11:7] : _GEN_158; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_164 = 5'h1e == _T_826 ? io_in[19:15] : _GEN_159; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_165 = 5'h1e == _T_826 ? io_in[24:20] : _GEN_160; // @[el2_ifu_compress.scala 195:12]
  wire [4:0] _GEN_166 = 5'h1e == _T_826 ? io_in[31:27] : _GEN_161; // @[el2_ifu_compress.scala 195:12]
  assign io_out_bits = 5'h1f == _T_826 ? io_in : _GEN_162; // @[el2_ifu_compress.scala 195:12]
  assign io_out_rd = 5'h1f == _T_826 ? io_in[11:7] : _GEN_163; // @[el2_ifu_compress.scala 195:12]
  assign io_out_rs1 = 5'h1f == _T_826 ? io_in[19:15] : _GEN_164; // @[el2_ifu_compress.scala 195:12]
  assign io_out_rs2 = 5'h1f == _T_826 ? io_in[24:20] : _GEN_165; // @[el2_ifu_compress.scala 195:12]
  assign io_out_rs3 = 5'h1f == _T_826 ? io_in[31:27] : _GEN_166; // @[el2_ifu_compress.scala 195:12]
  assign io_rvc = io_in[1:0] != 2'h3; // @[el2_ifu_compress.scala 193:12]
endmodule
