// NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE NOTE
// This is an automatically generated file by awais.abbas on Tue Dec 29 15:11:49 PKT 2020
//
// cmd:    swerv -target=default 
//

`include "common_defines.vh"
`undef ASSERT_ON
`undef TEC_RV_ICG
`define TEC_RV_ICG HDBLVT16_CKGTPLT_V5_12
`define PHYSICAL 1
