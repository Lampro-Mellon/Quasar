module rvclkhdr(
  output  io_l1clk,
  input   io_clk,
  input   io_en,
  input   io_scan_mode
);
  wire  clkhdr_Q; // @[el2_lib.scala 452:26]
  wire  clkhdr_CK; // @[el2_lib.scala 452:26]
  wire  clkhdr_EN; // @[el2_lib.scala 452:26]
  wire  clkhdr_SE; // @[el2_lib.scala 452:26]
  TEC_RV_ICG clkhdr ( // @[el2_lib.scala 452:26]
    .Q(clkhdr_Q),
    .CK(clkhdr_CK),
    .EN(clkhdr_EN),
    .SE(clkhdr_SE)
  );
  assign io_l1clk = clkhdr_Q; // @[el2_lib.scala 453:14]
  assign clkhdr_CK = io_clk; // @[el2_lib.scala 454:18]
  assign clkhdr_EN = io_en; // @[el2_lib.scala 455:18]
  assign clkhdr_SE = io_scan_mode; // @[el2_lib.scala 456:18]
endmodule
module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [63:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
`endif // RANDOMIZE_REG_INIT
  wire  rvclkhdr_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_1_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_1_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_1_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_1_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_2_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_2_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_2_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_2_io_scan_mode; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_3_io_l1clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_3_io_clk; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_3_io_en; // @[el2_lib.scala 461:22]
  wire  rvclkhdr_3_io_scan_mode; // @[el2_lib.scala 461:22]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 185:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 321:36]
  wire  _T_319 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 322:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_319; // @[el2_ifu_mem_ctl.scala 322:42]
  wire  _T = io_ifc_fetch_req_bf_raw | ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 186:53]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 253:30]
  wire  _T_1 = _T | miss_pending; // @[el2_ifu_mem_ctl.scala 186:71]
  wire  _T_2 = _T_1 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 186:86]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 548:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_319; // @[el2_ifu_mem_ctl.scala 550:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 187:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 308:63]
  wire [4:0] _GEN_460 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 666:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_460 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 666:53]
  wire [1:0] _GEN_461 = {{1'd0}, _T_319}; // @[el2_ifu_mem_ctl.scala 669:91]
  wire [1:0] _T_3095 = ic_fetch_val_shift_right[3:2] & _GEN_461; // @[el2_ifu_mem_ctl.scala 669:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 323:60]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:46]
  wire [1:0] _GEN_462 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 669:113]
  wire [1:0] _T_3096 = _T_3095 & _GEN_462; // @[el2_ifu_mem_ctl.scala 669:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 655:59]
  wire [1:0] _GEN_463 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 669:130]
  wire [1:0] _T_3097 = _T_3096 | _GEN_463; // @[el2_ifu_mem_ctl.scala 669:130]
  wire  _T_3098 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 669:154]
  wire [1:0] _GEN_464 = {{1'd0}, _T_3098}; // @[el2_ifu_mem_ctl.scala 669:152]
  wire [1:0] _T_3099 = _T_3097 & _GEN_464; // @[el2_ifu_mem_ctl.scala 669:152]
  wire [1:0] _T_3088 = ic_fetch_val_shift_right[1:0] & _GEN_461; // @[el2_ifu_mem_ctl.scala 669:91]
  wire [1:0] _T_3089 = _T_3088 & _GEN_462; // @[el2_ifu_mem_ctl.scala 669:113]
  wire [1:0] _T_3090 = _T_3089 | _GEN_463; // @[el2_ifu_mem_ctl.scala 669:130]
  wire [1:0] _T_3092 = _T_3090 & _GEN_464; // @[el2_ifu_mem_ctl.scala 669:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3099,_T_3092}; // @[Cat.scala 29:58]
  wire  _T_3199 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 311:30]
  wire  _T_3200 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 311:44]
  wire  _T_3201 = _T_3199 ^ _T_3200; // @[el2_lib.scala 311:35]
  wire [5:0] _T_3209 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 311:76]
  wire  _T_3210 = ^_T_3209; // @[el2_lib.scala 311:83]
  wire  _T_3211 = io_iccm_rd_data_ecc[37] ^ _T_3210; // @[el2_lib.scala 311:71]
  wire [6:0] _T_3218 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 311:103]
  wire [14:0] _T_3226 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3218}; // @[el2_lib.scala 311:103]
  wire  _T_3227 = ^_T_3226; // @[el2_lib.scala 311:110]
  wire  _T_3228 = io_iccm_rd_data_ecc[36] ^ _T_3227; // @[el2_lib.scala 311:98]
  wire [6:0] _T_3235 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 311:130]
  wire [14:0] _T_3243 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3235}; // @[el2_lib.scala 311:130]
  wire  _T_3244 = ^_T_3243; // @[el2_lib.scala 311:137]
  wire  _T_3245 = io_iccm_rd_data_ecc[35] ^ _T_3244; // @[el2_lib.scala 311:125]
  wire [8:0] _T_3254 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 311:157]
  wire [17:0] _T_3263 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3254}; // @[el2_lib.scala 311:157]
  wire  _T_3264 = ^_T_3263; // @[el2_lib.scala 311:164]
  wire  _T_3265 = io_iccm_rd_data_ecc[34] ^ _T_3264; // @[el2_lib.scala 311:152]
  wire [8:0] _T_3274 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 311:184]
  wire [17:0] _T_3283 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3274}; // @[el2_lib.scala 311:184]
  wire  _T_3284 = ^_T_3283; // @[el2_lib.scala 311:191]
  wire  _T_3285 = io_iccm_rd_data_ecc[33] ^ _T_3284; // @[el2_lib.scala 311:179]
  wire [8:0] _T_3294 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 311:211]
  wire [17:0] _T_3303 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3294}; // @[el2_lib.scala 311:211]
  wire  _T_3304 = ^_T_3303; // @[el2_lib.scala 311:218]
  wire  _T_3305 = io_iccm_rd_data_ecc[32] ^ _T_3304; // @[el2_lib.scala 311:206]
  wire [6:0] _T_3311 = {_T_3201,_T_3211,_T_3228,_T_3245,_T_3265,_T_3285,_T_3305}; // @[Cat.scala 29:58]
  wire  _T_3312 = _T_3311 != 7'h0; // @[el2_lib.scala 312:44]
  wire  _T_3313 = iccm_ecc_word_enable[0] & _T_3312; // @[el2_lib.scala 312:32]
  wire  _T_3315 = _T_3313 & _T_3311[6]; // @[el2_lib.scala 312:53]
  wire  _T_3584 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 311:30]
  wire  _T_3585 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 311:44]
  wire  _T_3586 = _T_3584 ^ _T_3585; // @[el2_lib.scala 311:35]
  wire [5:0] _T_3594 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 311:76]
  wire  _T_3595 = ^_T_3594; // @[el2_lib.scala 311:83]
  wire  _T_3596 = io_iccm_rd_data_ecc[76] ^ _T_3595; // @[el2_lib.scala 311:71]
  wire [6:0] _T_3603 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 311:103]
  wire [14:0] _T_3611 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3603}; // @[el2_lib.scala 311:103]
  wire  _T_3612 = ^_T_3611; // @[el2_lib.scala 311:110]
  wire  _T_3613 = io_iccm_rd_data_ecc[75] ^ _T_3612; // @[el2_lib.scala 311:98]
  wire [6:0] _T_3620 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 311:130]
  wire [14:0] _T_3628 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3620}; // @[el2_lib.scala 311:130]
  wire  _T_3629 = ^_T_3628; // @[el2_lib.scala 311:137]
  wire  _T_3630 = io_iccm_rd_data_ecc[74] ^ _T_3629; // @[el2_lib.scala 311:125]
  wire [8:0] _T_3639 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 311:157]
  wire [17:0] _T_3648 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3639}; // @[el2_lib.scala 311:157]
  wire  _T_3649 = ^_T_3648; // @[el2_lib.scala 311:164]
  wire  _T_3650 = io_iccm_rd_data_ecc[73] ^ _T_3649; // @[el2_lib.scala 311:152]
  wire [8:0] _T_3659 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 311:184]
  wire [17:0] _T_3668 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3659}; // @[el2_lib.scala 311:184]
  wire  _T_3669 = ^_T_3668; // @[el2_lib.scala 311:191]
  wire  _T_3670 = io_iccm_rd_data_ecc[72] ^ _T_3669; // @[el2_lib.scala 311:179]
  wire [8:0] _T_3679 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 311:211]
  wire [17:0] _T_3688 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3679}; // @[el2_lib.scala 311:211]
  wire  _T_3689 = ^_T_3688; // @[el2_lib.scala 311:218]
  wire  _T_3690 = io_iccm_rd_data_ecc[71] ^ _T_3689; // @[el2_lib.scala 311:206]
  wire [6:0] _T_3696 = {_T_3586,_T_3596,_T_3613,_T_3630,_T_3650,_T_3670,_T_3690}; // @[Cat.scala 29:58]
  wire  _T_3697 = _T_3696 != 7'h0; // @[el2_lib.scala 312:44]
  wire  _T_3698 = iccm_ecc_word_enable[1] & _T_3697; // @[el2_lib.scala 312:32]
  wire  _T_3700 = _T_3698 & _T_3696[6]; // @[el2_lib.scala 312:53]
  wire [1:0] iccm_single_ecc_error = {_T_3315,_T_3700}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 190:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 632:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 192:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 477:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 192:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 192:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 192:72]
  wire  _T_2492 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2497 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2517 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 527:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 391:42]
  wire  _T_2519 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 527:79]
  wire  _T_2520 = _T_2517 | _T_2519; // @[el2_ifu_mem_ctl.scala 527:56]
  wire  _T_2521 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 527:122]
  wire  _T_2522 = ~_T_2521; // @[el2_ifu_mem_ctl.scala 527:101]
  wire  _T_2523 = _T_2520 & _T_2522; // @[el2_ifu_mem_ctl.scala 527:99]
  wire  _T_2524 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2538 = io_ifu_fetch_val[0] & _T_319; // @[el2_ifu_mem_ctl.scala 534:45]
  wire  _T_2539 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 534:69]
  wire  _T_2540 = _T_2538 & _T_2539; // @[el2_ifu_mem_ctl.scala 534:67]
  wire  _T_2541 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_2524 ? _T_2540 : _T_2541; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2497 ? _T_2523 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2492 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 192:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 194:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 194:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 283:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 283:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 701:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 283:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 274:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 274:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 325:71]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 274:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 274:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 283:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 283:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 283:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 283:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 547:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 589:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 616:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 310:62]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 597:56]
  wire  _T_2638 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 614:69]
  wire  _T_2639 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 614:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2638 : _T_2639; // @[el2_ifu_mem_ctl.scala 614:28]
  wire  _T_2590 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 593:68]
  wire  _T_2591 = ic_act_miss_f | _T_2590; // @[el2_ifu_mem_ctl.scala 593:48]
  wire  bus_reset_data_beat_cnt = _T_2591 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 593:91]
  wire  _T_2587 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 592:50]
  wire  _T_2588 = bus_ifu_wr_en_ff & _T_2587; // @[el2_ifu_mem_ctl.scala 592:48]
  wire  _T_2589 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 592:72]
  wire  bus_inc_data_beat_cnt = _T_2588 & _T_2589; // @[el2_ifu_mem_ctl.scala 592:70]
  wire [2:0] _T_2595 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 596:115]
  wire [2:0] _T_2597 = bus_inc_data_beat_cnt ? _T_2595 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2592 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 594:32]
  wire  _T_2593 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 594:57]
  wire  bus_hold_data_beat_cnt = _T_2592 & _T_2593; // @[el2_ifu_mem_ctl.scala 594:55]
  wire [2:0] _T_2598 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2597 | _T_2598; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 194:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 195:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 194:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 195:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_319; // @[el2_ifu_mem_ctl.scala 201:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 427:45]
  wire  _T_2122 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 448:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 404:60]
  wire  _T_2153 = _T_2122 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2126 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2154 = _T_2126 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2161 = _T_2153 | _T_2154; // @[Mux.scala 27:72]
  wire  _T_2130 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2155 = _T_2130 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2162 = _T_2161 | _T_2155; // @[Mux.scala 27:72]
  wire  _T_2134 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2156 = _T_2134 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2163 = _T_2162 | _T_2156; // @[Mux.scala 27:72]
  wire  _T_2138 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2157 = _T_2138 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2164 = _T_2163 | _T_2157; // @[Mux.scala 27:72]
  wire  _T_2142 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2158 = _T_2142 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2165 = _T_2164 | _T_2158; // @[Mux.scala 27:72]
  wire  _T_2146 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2159 = _T_2146 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2166 = _T_2165 | _T_2159; // @[Mux.scala 27:72]
  wire  _T_2150 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 448:127]
  wire  _T_2160 = _T_2150 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2166 | _T_2160; // @[Mux.scala 27:72]
  wire  _T_2208 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 450:69]
  wire  _T_2209 = ic_miss_buff_data_valid_bypass_index & _T_2208; // @[el2_ifu_mem_ctl.scala 450:67]
  wire  _T_2211 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 450:91]
  wire  _T_2212 = _T_2209 & _T_2211; // @[el2_ifu_mem_ctl.scala 450:89]
  wire  _T_2217 = _T_2209 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 451:65]
  wire  _T_2218 = _T_2212 | _T_2217; // @[el2_ifu_mem_ctl.scala 450:112]
  wire  _T_2220 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 452:43]
  wire  _T_2223 = _T_2220 & _T_2211; // @[el2_ifu_mem_ctl.scala 452:65]
  wire  _T_2224 = _T_2218 | _T_2223; // @[el2_ifu_mem_ctl.scala 451:88]
  wire  _T_2228 = _T_2220 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 453:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 430:75]
  wire  _T_2168 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2192 = _T_2168 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2171 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2193 = _T_2171 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2192 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2174 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2194 = _T_2174 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2177 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2195 = _T_2177 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2180 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2196 = _T_2180 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2183 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2197 = _T_2183 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2204 = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2186 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2198 = _T_2186 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2205 = _T_2204 | _T_2198; // @[Mux.scala 27:72]
  wire  _T_2189 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 449:110]
  wire  _T_2199 = _T_2189 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2205 | _T_2199; // @[Mux.scala 27:72]
  wire  _T_2229 = _T_2228 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 453:87]
  wire  _T_2230 = _T_2224 | _T_2229; // @[el2_ifu_mem_ctl.scala 452:88]
  wire  _T_2234 = ic_miss_buff_data_valid_bypass_index & _T_2150; // @[el2_ifu_mem_ctl.scala 454:43]
  wire  miss_buff_hit_unq_f = _T_2230 | _T_2234; // @[el2_ifu_mem_ctl.scala 453:131]
  wire  _T_2250 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 459:55]
  wire  _T_2251 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 459:87]
  wire  _T_2252 = _T_2250 | _T_2251; // @[el2_ifu_mem_ctl.scala 459:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2252; // @[el2_ifu_mem_ctl.scala 459:41]
  wire  _T_2235 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 456:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 311:49]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 447:51]
  wire  _T_2236 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 456:68]
  wire  _T_2237 = miss_buff_hit_unq_f & _T_2236; // @[el2_ifu_mem_ctl.scala 456:66]
  wire  stream_hit_f = _T_2235 & _T_2237; // @[el2_ifu_mem_ctl.scala 456:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 278:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 278:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 278:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 599:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 626:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 205:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 205:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 205:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 205:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:16]
  wire  _T_44 = _T_42 & _T_319; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 207:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 208:49]
  wire  _T_54 = ic_byp_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 209:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 209:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 209:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 197:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 209:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 209:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_319; // @[el2_ifu_mem_ctl.scala 210:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 210:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 210:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 210:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 211:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 212:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 209:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 208:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 207:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 206:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2247 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 458:60]
  wire  _T_2248 = _T_2247 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 458:94]
  wire  stream_eol_f = _T_2248 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 458:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 220:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 220:87]
  wire  _T_113 = _T_111 & _T_2589; // @[el2_ifu_mem_ctl.scala 220:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 220:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 224:48]
  wire  _T_126 = _T_124 & _T_2589; // @[el2_ifu_mem_ctl.scala 224:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 284:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 284:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 284:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 285:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 284:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 285:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 339:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 285:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 285:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 285:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:50]
  wire  _T_137 = _T_135 & _T_2589; // @[el2_ifu_mem_ctl.scala 228:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 286:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 287:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 287:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 286:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:35]
  wire  _T_143 = _T_141 & _T_2589; // @[el2_ifu_mem_ctl.scala 229:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 234:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 233:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 238:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 238:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 195:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 195:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 195:26]
  wire  scnd_miss_req_in = _T_22 & _T_319; // @[el2_ifu_mem_ctl.scala 195:91]
  wire  _T_30 = ic_act_miss_f & _T_2589; // @[el2_ifu_mem_ctl.scala 202:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 213:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 213:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 213:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 213:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 217:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 217:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 221:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 225:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 230:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 235:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 235:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 254:95]
  wire  _T_175 = _T_2250 & _T_174; // @[el2_ifu_mem_ctl.scala 254:93]
  wire  crit_wd_byp_ok_ff = _T_2251 | _T_175; // @[el2_ifu_mem_ctl.scala 254:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 255:36]
  wire  _T_180 = _T_2250 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 255:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 255:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 255:70]
  wire  _T_184 = _T_2250 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 256:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 256:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 255:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 256:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 257:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 257:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 256:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 259:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 259:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:64]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 733:14]
  wire  _T_4763 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_4891 = _T_4763 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4764 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_4892 = _T_4764 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_5019 = _T_4891 | _T_4892; // @[Mux.scala 27:72]
  wire  _T_4765 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_4893 = _T_4765 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_5020 = _T_5019 | _T_4893; // @[Mux.scala 27:72]
  wire  _T_4766 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_4894 = _T_4766 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_5021 = _T_5020 | _T_4894; // @[Mux.scala 27:72]
  wire  _T_4767 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_4895 = _T_4767 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_5022 = _T_5021 | _T_4895; // @[Mux.scala 27:72]
  wire  _T_4768 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_4896 = _T_4768 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_5023 = _T_5022 | _T_4896; // @[Mux.scala 27:72]
  wire  _T_4769 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_4897 = _T_4769 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_5024 = _T_5023 | _T_4897; // @[Mux.scala 27:72]
  wire  _T_4770 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_4898 = _T_4770 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_5025 = _T_5024 | _T_4898; // @[Mux.scala 27:72]
  wire  _T_4771 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_4899 = _T_4771 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_5026 = _T_5025 | _T_4899; // @[Mux.scala 27:72]
  wire  _T_4772 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_4900 = _T_4772 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_5027 = _T_5026 | _T_4900; // @[Mux.scala 27:72]
  wire  _T_4773 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_4901 = _T_4773 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_5028 = _T_5027 | _T_4901; // @[Mux.scala 27:72]
  wire  _T_4774 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_4902 = _T_4774 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_5029 = _T_5028 | _T_4902; // @[Mux.scala 27:72]
  wire  _T_4775 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_4903 = _T_4775 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_5030 = _T_5029 | _T_4903; // @[Mux.scala 27:72]
  wire  _T_4776 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_4904 = _T_4776 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_5031 = _T_5030 | _T_4904; // @[Mux.scala 27:72]
  wire  _T_4777 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_4905 = _T_4777 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_5032 = _T_5031 | _T_4905; // @[Mux.scala 27:72]
  wire  _T_4778 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_4906 = _T_4778 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_5033 = _T_5032 | _T_4906; // @[Mux.scala 27:72]
  wire  _T_4779 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_4907 = _T_4779 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_5034 = _T_5033 | _T_4907; // @[Mux.scala 27:72]
  wire  _T_4780 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_4908 = _T_4780 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_5035 = _T_5034 | _T_4908; // @[Mux.scala 27:72]
  wire  _T_4781 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_4909 = _T_4781 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_5036 = _T_5035 | _T_4909; // @[Mux.scala 27:72]
  wire  _T_4782 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_4910 = _T_4782 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_5037 = _T_5036 | _T_4910; // @[Mux.scala 27:72]
  wire  _T_4783 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_4911 = _T_4783 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_5038 = _T_5037 | _T_4911; // @[Mux.scala 27:72]
  wire  _T_4784 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_4912 = _T_4784 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_5039 = _T_5038 | _T_4912; // @[Mux.scala 27:72]
  wire  _T_4785 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_4913 = _T_4785 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_5040 = _T_5039 | _T_4913; // @[Mux.scala 27:72]
  wire  _T_4786 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_4914 = _T_4786 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_5041 = _T_5040 | _T_4914; // @[Mux.scala 27:72]
  wire  _T_4787 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_4915 = _T_4787 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_5042 = _T_5041 | _T_4915; // @[Mux.scala 27:72]
  wire  _T_4788 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_4916 = _T_4788 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_5043 = _T_5042 | _T_4916; // @[Mux.scala 27:72]
  wire  _T_4789 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_4917 = _T_4789 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_5044 = _T_5043 | _T_4917; // @[Mux.scala 27:72]
  wire  _T_4790 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_4918 = _T_4790 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_5045 = _T_5044 | _T_4918; // @[Mux.scala 27:72]
  wire  _T_4791 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_4919 = _T_4791 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_5046 = _T_5045 | _T_4919; // @[Mux.scala 27:72]
  wire  _T_4792 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_4920 = _T_4792 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_5047 = _T_5046 | _T_4920; // @[Mux.scala 27:72]
  wire  _T_4793 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_4921 = _T_4793 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_5048 = _T_5047 | _T_4921; // @[Mux.scala 27:72]
  wire  _T_4794 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_4922 = _T_4794 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_5049 = _T_5048 | _T_4922; // @[Mux.scala 27:72]
  wire  _T_4795 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_4923 = _T_4795 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_5050 = _T_5049 | _T_4923; // @[Mux.scala 27:72]
  wire  _T_4796 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_4924 = _T_4796 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_5051 = _T_5050 | _T_4924; // @[Mux.scala 27:72]
  wire  _T_4797 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_4925 = _T_4797 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_5052 = _T_5051 | _T_4925; // @[Mux.scala 27:72]
  wire  _T_4798 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_4926 = _T_4798 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_5053 = _T_5052 | _T_4926; // @[Mux.scala 27:72]
  wire  _T_4799 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_4927 = _T_4799 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_5054 = _T_5053 | _T_4927; // @[Mux.scala 27:72]
  wire  _T_4800 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_4928 = _T_4800 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_5055 = _T_5054 | _T_4928; // @[Mux.scala 27:72]
  wire  _T_4801 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_4929 = _T_4801 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_5056 = _T_5055 | _T_4929; // @[Mux.scala 27:72]
  wire  _T_4802 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_4930 = _T_4802 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_5057 = _T_5056 | _T_4930; // @[Mux.scala 27:72]
  wire  _T_4803 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_4931 = _T_4803 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_5058 = _T_5057 | _T_4931; // @[Mux.scala 27:72]
  wire  _T_4804 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_4932 = _T_4804 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_5059 = _T_5058 | _T_4932; // @[Mux.scala 27:72]
  wire  _T_4805 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_4933 = _T_4805 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_5060 = _T_5059 | _T_4933; // @[Mux.scala 27:72]
  wire  _T_4806 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_4934 = _T_4806 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_5061 = _T_5060 | _T_4934; // @[Mux.scala 27:72]
  wire  _T_4807 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_4935 = _T_4807 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_5062 = _T_5061 | _T_4935; // @[Mux.scala 27:72]
  wire  _T_4808 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_4936 = _T_4808 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_5063 = _T_5062 | _T_4936; // @[Mux.scala 27:72]
  wire  _T_4809 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_4937 = _T_4809 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_5064 = _T_5063 | _T_4937; // @[Mux.scala 27:72]
  wire  _T_4810 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_4938 = _T_4810 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_5065 = _T_5064 | _T_4938; // @[Mux.scala 27:72]
  wire  _T_4811 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_4939 = _T_4811 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_5066 = _T_5065 | _T_4939; // @[Mux.scala 27:72]
  wire  _T_4812 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_4940 = _T_4812 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_5067 = _T_5066 | _T_4940; // @[Mux.scala 27:72]
  wire  _T_4813 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_4941 = _T_4813 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_5068 = _T_5067 | _T_4941; // @[Mux.scala 27:72]
  wire  _T_4814 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_4942 = _T_4814 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_5069 = _T_5068 | _T_4942; // @[Mux.scala 27:72]
  wire  _T_4815 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_4943 = _T_4815 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_5070 = _T_5069 | _T_4943; // @[Mux.scala 27:72]
  wire  _T_4816 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_4944 = _T_4816 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_5071 = _T_5070 | _T_4944; // @[Mux.scala 27:72]
  wire  _T_4817 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_4945 = _T_4817 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_5072 = _T_5071 | _T_4945; // @[Mux.scala 27:72]
  wire  _T_4818 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_4946 = _T_4818 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_5073 = _T_5072 | _T_4946; // @[Mux.scala 27:72]
  wire  _T_4819 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_4947 = _T_4819 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_5074 = _T_5073 | _T_4947; // @[Mux.scala 27:72]
  wire  _T_4820 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_4948 = _T_4820 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_5075 = _T_5074 | _T_4948; // @[Mux.scala 27:72]
  wire  _T_4821 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_4949 = _T_4821 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_5076 = _T_5075 | _T_4949; // @[Mux.scala 27:72]
  wire  _T_4822 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_4950 = _T_4822 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_5077 = _T_5076 | _T_4950; // @[Mux.scala 27:72]
  wire  _T_4823 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_4951 = _T_4823 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_5078 = _T_5077 | _T_4951; // @[Mux.scala 27:72]
  wire  _T_4824 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_4952 = _T_4824 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_5079 = _T_5078 | _T_4952; // @[Mux.scala 27:72]
  wire  _T_4825 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_4953 = _T_4825 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_5080 = _T_5079 | _T_4953; // @[Mux.scala 27:72]
  wire  _T_4826 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_4954 = _T_4826 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_5081 = _T_5080 | _T_4954; // @[Mux.scala 27:72]
  wire  _T_4827 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_4955 = _T_4827 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_5082 = _T_5081 | _T_4955; // @[Mux.scala 27:72]
  wire  _T_4828 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_4956 = _T_4828 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_5083 = _T_5082 | _T_4956; // @[Mux.scala 27:72]
  wire  _T_4829 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_4957 = _T_4829 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_5084 = _T_5083 | _T_4957; // @[Mux.scala 27:72]
  wire  _T_4830 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_4958 = _T_4830 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_5085 = _T_5084 | _T_4958; // @[Mux.scala 27:72]
  wire  _T_4831 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_4959 = _T_4831 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_5086 = _T_5085 | _T_4959; // @[Mux.scala 27:72]
  wire  _T_4832 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_4960 = _T_4832 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_5087 = _T_5086 | _T_4960; // @[Mux.scala 27:72]
  wire  _T_4833 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_4961 = _T_4833 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_5088 = _T_5087 | _T_4961; // @[Mux.scala 27:72]
  wire  _T_4834 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_4962 = _T_4834 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_5089 = _T_5088 | _T_4962; // @[Mux.scala 27:72]
  wire  _T_4835 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_4963 = _T_4835 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_5090 = _T_5089 | _T_4963; // @[Mux.scala 27:72]
  wire  _T_4836 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_4964 = _T_4836 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_5091 = _T_5090 | _T_4964; // @[Mux.scala 27:72]
  wire  _T_4837 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_4965 = _T_4837 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_5092 = _T_5091 | _T_4965; // @[Mux.scala 27:72]
  wire  _T_4838 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_4966 = _T_4838 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_5093 = _T_5092 | _T_4966; // @[Mux.scala 27:72]
  wire  _T_4839 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_4967 = _T_4839 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_5094 = _T_5093 | _T_4967; // @[Mux.scala 27:72]
  wire  _T_4840 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_4968 = _T_4840 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_5095 = _T_5094 | _T_4968; // @[Mux.scala 27:72]
  wire  _T_4841 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_4969 = _T_4841 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_5096 = _T_5095 | _T_4969; // @[Mux.scala 27:72]
  wire  _T_4842 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_4970 = _T_4842 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_5097 = _T_5096 | _T_4970; // @[Mux.scala 27:72]
  wire  _T_4843 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_4971 = _T_4843 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_5098 = _T_5097 | _T_4971; // @[Mux.scala 27:72]
  wire  _T_4844 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_4972 = _T_4844 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_5099 = _T_5098 | _T_4972; // @[Mux.scala 27:72]
  wire  _T_4845 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_4973 = _T_4845 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_5100 = _T_5099 | _T_4973; // @[Mux.scala 27:72]
  wire  _T_4846 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_4974 = _T_4846 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_5101 = _T_5100 | _T_4974; // @[Mux.scala 27:72]
  wire  _T_4847 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_4975 = _T_4847 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_5102 = _T_5101 | _T_4975; // @[Mux.scala 27:72]
  wire  _T_4848 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_4976 = _T_4848 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_5103 = _T_5102 | _T_4976; // @[Mux.scala 27:72]
  wire  _T_4849 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_4977 = _T_4849 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_5104 = _T_5103 | _T_4977; // @[Mux.scala 27:72]
  wire  _T_4850 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_4978 = _T_4850 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_5105 = _T_5104 | _T_4978; // @[Mux.scala 27:72]
  wire  _T_4851 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_4979 = _T_4851 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_5106 = _T_5105 | _T_4979; // @[Mux.scala 27:72]
  wire  _T_4852 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_4980 = _T_4852 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_5107 = _T_5106 | _T_4980; // @[Mux.scala 27:72]
  wire  _T_4853 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_4981 = _T_4853 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_5108 = _T_5107 | _T_4981; // @[Mux.scala 27:72]
  wire  _T_4854 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_4982 = _T_4854 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_5109 = _T_5108 | _T_4982; // @[Mux.scala 27:72]
  wire  _T_4855 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_4983 = _T_4855 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_5110 = _T_5109 | _T_4983; // @[Mux.scala 27:72]
  wire  _T_4856 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_4984 = _T_4856 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_5111 = _T_5110 | _T_4984; // @[Mux.scala 27:72]
  wire  _T_4857 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_4985 = _T_4857 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_5112 = _T_5111 | _T_4985; // @[Mux.scala 27:72]
  wire  _T_4858 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_4986 = _T_4858 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_5113 = _T_5112 | _T_4986; // @[Mux.scala 27:72]
  wire  _T_4859 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_4987 = _T_4859 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_5114 = _T_5113 | _T_4987; // @[Mux.scala 27:72]
  wire  _T_4860 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_4988 = _T_4860 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_5115 = _T_5114 | _T_4988; // @[Mux.scala 27:72]
  wire  _T_4861 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_4989 = _T_4861 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_5116 = _T_5115 | _T_4989; // @[Mux.scala 27:72]
  wire  _T_4862 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_4990 = _T_4862 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_5117 = _T_5116 | _T_4990; // @[Mux.scala 27:72]
  wire  _T_4863 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_4991 = _T_4863 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_5118 = _T_5117 | _T_4991; // @[Mux.scala 27:72]
  wire  _T_4864 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_4992 = _T_4864 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_5119 = _T_5118 | _T_4992; // @[Mux.scala 27:72]
  wire  _T_4865 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_4993 = _T_4865 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_5120 = _T_5119 | _T_4993; // @[Mux.scala 27:72]
  wire  _T_4866 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_4994 = _T_4866 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_5121 = _T_5120 | _T_4994; // @[Mux.scala 27:72]
  wire  _T_4867 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_4995 = _T_4867 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_5122 = _T_5121 | _T_4995; // @[Mux.scala 27:72]
  wire  _T_4868 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_4996 = _T_4868 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_5123 = _T_5122 | _T_4996; // @[Mux.scala 27:72]
  wire  _T_4869 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_4997 = _T_4869 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_5124 = _T_5123 | _T_4997; // @[Mux.scala 27:72]
  wire  _T_4870 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_4998 = _T_4870 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_5125 = _T_5124 | _T_4998; // @[Mux.scala 27:72]
  wire  _T_4871 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_4999 = _T_4871 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_5126 = _T_5125 | _T_4999; // @[Mux.scala 27:72]
  wire  _T_4872 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_5000 = _T_4872 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_5127 = _T_5126 | _T_5000; // @[Mux.scala 27:72]
  wire  _T_4873 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_5001 = _T_4873 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_5128 = _T_5127 | _T_5001; // @[Mux.scala 27:72]
  wire  _T_4874 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_5002 = _T_4874 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_5129 = _T_5128 | _T_5002; // @[Mux.scala 27:72]
  wire  _T_4875 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_5003 = _T_4875 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_5130 = _T_5129 | _T_5003; // @[Mux.scala 27:72]
  wire  _T_4876 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_5004 = _T_4876 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_5131 = _T_5130 | _T_5004; // @[Mux.scala 27:72]
  wire  _T_4877 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_5005 = _T_4877 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_5132 = _T_5131 | _T_5005; // @[Mux.scala 27:72]
  wire  _T_4878 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_5006 = _T_4878 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_5133 = _T_5132 | _T_5006; // @[Mux.scala 27:72]
  wire  _T_4879 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_5007 = _T_4879 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_5134 = _T_5133 | _T_5007; // @[Mux.scala 27:72]
  wire  _T_4880 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_5008 = _T_4880 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_5135 = _T_5134 | _T_5008; // @[Mux.scala 27:72]
  wire  _T_4881 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_5009 = _T_4881 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_5136 = _T_5135 | _T_5009; // @[Mux.scala 27:72]
  wire  _T_4882 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_5010 = _T_4882 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_5137 = _T_5136 | _T_5010; // @[Mux.scala 27:72]
  wire  _T_4883 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_5011 = _T_4883 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_5138 = _T_5137 | _T_5011; // @[Mux.scala 27:72]
  wire  _T_4884 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_5012 = _T_4884 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_5139 = _T_5138 | _T_5012; // @[Mux.scala 27:72]
  wire  _T_4885 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_5013 = _T_4885 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_5140 = _T_5139 | _T_5013; // @[Mux.scala 27:72]
  wire  _T_4886 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_5014 = _T_4886 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_5141 = _T_5140 | _T_5014; // @[Mux.scala 27:72]
  wire  _T_4887 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_5015 = _T_4887 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_5142 = _T_5141 | _T_5015; // @[Mux.scala 27:72]
  wire  _T_4888 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_5016 = _T_4888 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5143 = _T_5142 | _T_5016; // @[Mux.scala 27:72]
  wire  _T_4889 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_5017 = _T_4889 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5144 = _T_5143 | _T_5017; // @[Mux.scala 27:72]
  wire  _T_4890 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 729:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_5018 = _T_4890 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5144 | _T_5018; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 262:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 262:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:58]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 264:67]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 266:54]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 271:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 276:59]
  wire  _T_214 = _T_212 | _T_2235; // @[el2_ifu_mem_ctl.scala 276:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 276:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 282:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 282:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 282:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 282:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 289:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 289:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 289:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 290:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 290:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 293:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 293:135]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2659 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 622:48]
  wire  _T_2660 = _T_2659 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 622:52]
  wire  bus_ifu_wr_data_error_ff = _T_2660 & miss_pending; // @[el2_ifu_mem_ctl.scala 622:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 367:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 366:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 293:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 293:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 296:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 296:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 317:59]
  wire  _T_10352 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 785:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 318:53]
  wire  _T_10354 = _T_10352 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 785:51]
  wire  _T_10356 = _T_10354 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 785:67]
  wire  _T_10358 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 785:86]
  wire  replace_way_mb_any_0 = _T_10356 | _T_10358; // @[el2_ifu_mem_ctl.scala 785:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10361 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:50]
  wire  _T_10363 = _T_10361 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:66]
  wire  _T_10365 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:85]
  wire  _T_10367 = _T_10365 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:100]
  wire  replace_way_mb_any_1 = _T_10363 | _T_10367; // @[el2_ifu_mem_ctl.scala 786:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 301:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 301:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 302:56]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 305:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 305:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 305:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 305:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 307:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 316:48]
  wire  _T_309 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 315:57]
  wire  _T_315 = _T_2250 & flush_final_f; // @[el2_ifu_mem_ctl.scala 320:87]
  wire  _T_316 = ~_T_315; // @[el2_ifu_mem_ctl.scala 320:55]
  wire  _T_317 = io_ifc_fetch_req_bf & _T_316; // @[el2_ifu_mem_ctl.scala 320:53]
  wire  _T_2242 = ~_T_2237; // @[el2_ifu_mem_ctl.scala 457:46]
  wire  _T_2243 = _T_2235 & _T_2242; // @[el2_ifu_mem_ctl.scala 457:44]
  wire  stream_miss_f = _T_2243 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 457:84]
  wire  _T_318 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 320:106]
  wire  ifc_fetch_req_qual_bf = _T_317 & _T_318; // @[el2_ifu_mem_ctl.scala 320:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 326:68]
  reg [2:0] bus_rd_addr_count; // @[el2_ifu_mem_ctl.scala 604:55]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_325 = _T_239 | _T_2235; // @[el2_ifu_mem_ctl.scala 328:55]
  wire  _T_328 = _T_325 & _T_56; // @[el2_ifu_mem_ctl.scala 328:82]
  wire  _T_2256 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 462:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2256}; // @[Cat.scala 29:58]
  wire  _T_2257 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2281 = _T_2257 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2260 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2282 = _T_2260 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2281 | _T_2282; // @[Mux.scala 27:72]
  wire  _T_2263 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2283 = _T_2263 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2289 | _T_2283; // @[Mux.scala 27:72]
  wire  _T_2266 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2284 = _T_2266 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2290 | _T_2284; // @[Mux.scala 27:72]
  wire  _T_2269 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2285 = _T_2269 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2291 | _T_2285; // @[Mux.scala 27:72]
  wire  _T_2272 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2286 = _T_2272 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2293 = _T_2292 | _T_2286; // @[Mux.scala 27:72]
  wire  _T_2275 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2287 = _T_2275 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2294 = _T_2293 | _T_2287; // @[Mux.scala 27:72]
  wire  _T_2278 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 463:81]
  wire  _T_2288 = _T_2278 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2294 | _T_2288; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 464:46]
  wire  _T_332 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 332:35]
  wire  _T_334 = _T_332 & _T_17; // @[el2_ifu_mem_ctl.scala 332:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 619:61]
  wire  _T_2653 = ic_act_miss_f_delayed & _T_2251; // @[el2_ifu_mem_ctl.scala 620:53]
  wire  reset_tag_valid_for_miss = _T_2653 & _T_17; // @[el2_ifu_mem_ctl.scala 620:84]
  wire  sel_mb_addr = _T_334 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 332:79]
  wire [30:0] _T_338 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_339 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 334:37]
  wire [30:0] _T_340 = sel_mb_addr ? _T_338 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_341 = _T_339 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_340 | _T_341; // @[Mux.scala 27:72]
  wire  _T_346 = _T_334 & last_beat; // @[el2_ifu_mem_ctl.scala 336:84]
  wire  _T_2647 = ~_T_2659; // @[el2_ifu_mem_ctl.scala 617:84]
  wire  _T_2648 = _T_100 & _T_2647; // @[el2_ifu_mem_ctl.scala 617:82]
  wire  bus_ifu_wr_en_ff_q = _T_2648 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 617:108]
  wire  sel_mb_status_addr = _T_346 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 336:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_338 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 337:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_569 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 394:13]
  wire  _T_570 = ^_T_569; // @[el2_lib.scala 394:20]
  wire [6:0] _T_576 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 394:30]
  wire [7:0] _T_583 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 394:30]
  wire [14:0] _T_584 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_576}; // @[el2_lib.scala 394:30]
  wire [7:0] _T_591 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 394:30]
  wire [30:0] _T_600 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_584}; // @[el2_lib.scala 394:30]
  wire  _T_601 = ^_T_600; // @[el2_lib.scala 394:37]
  wire [6:0] _T_607 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 394:47]
  wire [14:0] _T_615 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_607}; // @[el2_lib.scala 394:47]
  wire [30:0] _T_631 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_591,_T_615}; // @[el2_lib.scala 394:47]
  wire  _T_632 = ^_T_631; // @[el2_lib.scala 394:54]
  wire [6:0] _T_638 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 394:64]
  wire [14:0] _T_646 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_638}; // @[el2_lib.scala 394:64]
  wire [30:0] _T_662 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_583,_T_646}; // @[el2_lib.scala 394:64]
  wire  _T_663 = ^_T_662; // @[el2_lib.scala 394:71]
  wire [7:0] _T_670 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 394:81]
  wire [16:0] _T_679 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_670}; // @[el2_lib.scala 394:81]
  wire [8:0] _T_687 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 394:81]
  wire [17:0] _T_696 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_687}; // @[el2_lib.scala 394:81]
  wire [34:0] _T_697 = {_T_696,_T_679}; // @[el2_lib.scala 394:81]
  wire  _T_698 = ^_T_697; // @[el2_lib.scala 394:88]
  wire [7:0] _T_705 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 394:98]
  wire [16:0] _T_714 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_705}; // @[el2_lib.scala 394:98]
  wire [8:0] _T_722 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 394:98]
  wire [17:0] _T_731 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_722}; // @[el2_lib.scala 394:98]
  wire [34:0] _T_732 = {_T_731,_T_714}; // @[el2_lib.scala 394:98]
  wire  _T_733 = ^_T_732; // @[el2_lib.scala 394:105]
  wire [7:0] _T_740 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 394:115]
  wire [16:0] _T_749 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_740}; // @[el2_lib.scala 394:115]
  wire [8:0] _T_757 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 394:115]
  wire [17:0] _T_766 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_757}; // @[el2_lib.scala 394:115]
  wire [34:0] _T_767 = {_T_766,_T_749}; // @[el2_lib.scala 394:115]
  wire  _T_768 = ^_T_767; // @[el2_lib.scala 394:122]
  wire [3:0] _T_2297 = {ifu_bus_rid_ff[2:1],_T_2256,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2298 = _T_2297 == 4'h0; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2345 = _T_2298 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2301 = _T_2297 == 4'h1; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2346 = _T_2301 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2345 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2304 = _T_2297 == 4'h2; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2347 = _T_2304 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire  _T_2307 = _T_2297 == 4'h3; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2348 = _T_2307 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2363 = _T_2362 | _T_2348; // @[Mux.scala 27:72]
  wire  _T_2310 = _T_2297 == 4'h4; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2349 = _T_2310 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2364 = _T_2363 | _T_2349; // @[Mux.scala 27:72]
  wire  _T_2313 = _T_2297 == 4'h5; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2350 = _T_2313 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2365 = _T_2364 | _T_2350; // @[Mux.scala 27:72]
  wire  _T_2316 = _T_2297 == 4'h6; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2351 = _T_2316 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2366 = _T_2365 | _T_2351; // @[Mux.scala 27:72]
  wire  _T_2319 = _T_2297 == 4'h7; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2352 = _T_2319 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2367 = _T_2366 | _T_2352; // @[Mux.scala 27:72]
  wire  _T_2322 = _T_2297 == 4'h8; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2353 = _T_2322 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2368 = _T_2367 | _T_2353; // @[Mux.scala 27:72]
  wire  _T_2325 = _T_2297 == 4'h9; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2354 = _T_2325 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2369 = _T_2368 | _T_2354; // @[Mux.scala 27:72]
  wire  _T_2328 = _T_2297 == 4'ha; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2355 = _T_2328 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 27:72]
  wire  _T_2331 = _T_2297 == 4'hb; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2356 = _T_2331 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2371 = _T_2370 | _T_2356; // @[Mux.scala 27:72]
  wire  _T_2334 = _T_2297 == 4'hc; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2357 = _T_2334 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2372 = _T_2371 | _T_2357; // @[Mux.scala 27:72]
  wire  _T_2337 = _T_2297 == 4'hd; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2358 = _T_2337 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2373 = _T_2372 | _T_2358; // @[Mux.scala 27:72]
  wire  _T_2340 = _T_2297 == 4'he; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2359 = _T_2340 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2374 = _T_2373 | _T_2359; // @[Mux.scala 27:72]
  wire  _T_2343 = _T_2297 == 4'hf; // @[el2_ifu_mem_ctl.scala 465:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2360 = _T_2343 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2375 = _T_2374 | _T_2360; // @[Mux.scala 27:72]
  wire [3:0] _T_2377 = {ifu_bus_rid_ff[2:1],_T_2256,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2378 = _T_2377 == 4'h0; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2425 = _T_2378 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2381 = _T_2377 == 4'h1; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2426 = _T_2381 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2441 = _T_2425 | _T_2426; // @[Mux.scala 27:72]
  wire  _T_2384 = _T_2377 == 4'h2; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2427 = _T_2384 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2442 = _T_2441 | _T_2427; // @[Mux.scala 27:72]
  wire  _T_2387 = _T_2377 == 4'h3; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2428 = _T_2387 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2443 = _T_2442 | _T_2428; // @[Mux.scala 27:72]
  wire  _T_2390 = _T_2377 == 4'h4; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2429 = _T_2390 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2444 = _T_2443 | _T_2429; // @[Mux.scala 27:72]
  wire  _T_2393 = _T_2377 == 4'h5; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2430 = _T_2393 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2445 = _T_2444 | _T_2430; // @[Mux.scala 27:72]
  wire  _T_2396 = _T_2377 == 4'h6; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2431 = _T_2396 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2446 = _T_2445 | _T_2431; // @[Mux.scala 27:72]
  wire  _T_2399 = _T_2377 == 4'h7; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2432 = _T_2399 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2447 = _T_2446 | _T_2432; // @[Mux.scala 27:72]
  wire  _T_2402 = _T_2377 == 4'h8; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2433 = _T_2402 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2448 = _T_2447 | _T_2433; // @[Mux.scala 27:72]
  wire  _T_2405 = _T_2377 == 4'h9; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2434 = _T_2405 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2449 = _T_2448 | _T_2434; // @[Mux.scala 27:72]
  wire  _T_2408 = _T_2377 == 4'ha; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2435 = _T_2408 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2450 = _T_2449 | _T_2435; // @[Mux.scala 27:72]
  wire  _T_2411 = _T_2377 == 4'hb; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2436 = _T_2411 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2451 = _T_2450 | _T_2436; // @[Mux.scala 27:72]
  wire  _T_2414 = _T_2377 == 4'hc; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2437 = _T_2414 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2452 = _T_2451 | _T_2437; // @[Mux.scala 27:72]
  wire  _T_2417 = _T_2377 == 4'hd; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2438 = _T_2417 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2453 = _T_2452 | _T_2438; // @[Mux.scala 27:72]
  wire  _T_2420 = _T_2377 == 4'he; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2439 = _T_2420 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2454 = _T_2453 | _T_2439; // @[Mux.scala 27:72]
  wire  _T_2423 = _T_2377 == 4'hf; // @[el2_ifu_mem_ctl.scala 466:66]
  wire [31:0] _T_2440 = _T_2423 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2455 = _T_2454 | _T_2440; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2375,_T_2455}; // @[Cat.scala 29:58]
  wire [6:0] _T_991 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 394:13]
  wire  _T_992 = ^_T_991; // @[el2_lib.scala 394:20]
  wire [6:0] _T_998 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 394:30]
  wire [7:0] _T_1005 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 394:30]
  wire [14:0] _T_1006 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_998}; // @[el2_lib.scala 394:30]
  wire [7:0] _T_1013 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 394:30]
  wire [30:0] _T_1022 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1006}; // @[el2_lib.scala 394:30]
  wire  _T_1023 = ^_T_1022; // @[el2_lib.scala 394:37]
  wire [6:0] _T_1029 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 394:47]
  wire [14:0] _T_1037 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1029}; // @[el2_lib.scala 394:47]
  wire [30:0] _T_1053 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1013,_T_1037}; // @[el2_lib.scala 394:47]
  wire  _T_1054 = ^_T_1053; // @[el2_lib.scala 394:54]
  wire [6:0] _T_1060 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 394:64]
  wire [14:0] _T_1068 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1060}; // @[el2_lib.scala 394:64]
  wire [30:0] _T_1084 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1005,_T_1068}; // @[el2_lib.scala 394:64]
  wire  _T_1085 = ^_T_1084; // @[el2_lib.scala 394:71]
  wire [7:0] _T_1092 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 394:81]
  wire [16:0] _T_1101 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1092}; // @[el2_lib.scala 394:81]
  wire [8:0] _T_1109 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 394:81]
  wire [17:0] _T_1118 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1109}; // @[el2_lib.scala 394:81]
  wire [34:0] _T_1119 = {_T_1118,_T_1101}; // @[el2_lib.scala 394:81]
  wire  _T_1120 = ^_T_1119; // @[el2_lib.scala 394:88]
  wire [7:0] _T_1127 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 394:98]
  wire [16:0] _T_1136 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1127}; // @[el2_lib.scala 394:98]
  wire [8:0] _T_1144 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 394:98]
  wire [17:0] _T_1153 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1144}; // @[el2_lib.scala 394:98]
  wire [34:0] _T_1154 = {_T_1153,_T_1136}; // @[el2_lib.scala 394:98]
  wire  _T_1155 = ^_T_1154; // @[el2_lib.scala 394:105]
  wire [7:0] _T_1162 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 394:115]
  wire [16:0] _T_1171 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1162}; // @[el2_lib.scala 394:115]
  wire [8:0] _T_1179 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 394:115]
  wire [17:0] _T_1188 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1179}; // @[el2_lib.scala 394:115]
  wire [34:0] _T_1189 = {_T_1188,_T_1171}; // @[el2_lib.scala 394:115]
  wire  _T_1190 = ^_T_1189; // @[el2_lib.scala 394:122]
  wire [70:0] _T_1235 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1234 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2375,_T_2455}; // @[Cat.scala 29:58]
  wire [141:0] _T_1236 = {_T_570,_T_601,_T_632,_T_663,_T_698,_T_733,_T_768,ifu_bus_rdata_ff,_T_1234}; // @[Cat.scala 29:58]
  wire [141:0] _T_1239 = {_T_992,_T_1023,_T_1054,_T_1085,_T_1120,_T_1155,_T_1190,_T_2375,_T_2455,_T_1235}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1236 : _T_1239; // @[el2_ifu_mem_ctl.scala 358:28]
  wire  _T_1198 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 348:56]
  wire  _T_1199 = _T_1198 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 348:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 412:28]
  wire  _T_1415 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 615:35]
  wire  _T_1284 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1341 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 403:118]
  wire  _T_1342 = ic_miss_buff_data_valid[0] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1342; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1438 = _T_1415 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1418 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1345 = ic_miss_buff_data_valid[1] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1345; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1439 = _T_1418 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1438 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1421 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1348 = ic_miss_buff_data_valid[2] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1348; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1440 = _T_1421 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1424 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1351 = ic_miss_buff_data_valid[3] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1351; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1441 = _T_1424 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1427 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1354 = ic_miss_buff_data_valid[4] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1354; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1442 = _T_1427 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1430 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1357 = ic_miss_buff_data_valid[5] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1357; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1443 = _T_1430 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1450 = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1433 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1290 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1290; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1360 = ic_miss_buff_data_valid[6] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1360; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1444 = _T_1433 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1451 = _T_1450 | _T_1444; // @[Mux.scala 27:72]
  wire  _T_1436 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 414:114]
  wire  _T_1291 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 397:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1291; // @[el2_ifu_mem_ctl.scala 397:73]
  wire  _T_1363 = ic_miss_buff_data_valid[7] & _T_1341; // @[el2_ifu_mem_ctl.scala 403:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1363; // @[el2_ifu_mem_ctl.scala 403:88]
  wire  _T_1445 = _T_1436 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1451 | _T_1445; // @[Mux.scala 27:72]
  wire  _T_1454 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 415:58]
  wire  _T_1455 = bypass_valid_value_check & _T_1454; // @[el2_ifu_mem_ctl.scala 415:56]
  wire  _T_1457 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 415:77]
  wire  _T_1458 = _T_1455 & _T_1457; // @[el2_ifu_mem_ctl.scala 415:75]
  wire  _T_1463 = _T_1455 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 416:75]
  wire  _T_1464 = _T_1458 | _T_1463; // @[el2_ifu_mem_ctl.scala 415:95]
  wire  _T_1466 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 417:56]
  wire  _T_1469 = _T_1466 & _T_1457; // @[el2_ifu_mem_ctl.scala 417:74]
  wire  _T_1470 = _T_1464 | _T_1469; // @[el2_ifu_mem_ctl.scala 416:94]
  wire  _T_1474 = _T_1466 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 418:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 413:70]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1491 = _T_1475 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1492 = _T_1477 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1491 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1479 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1493 = _T_1479 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1499 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1481 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1494 = _T_1481 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1500 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1483 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1495 = _T_1483 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1501 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1485 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1496 = _T_1485 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1502 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1487 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1497 = _T_1487 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1504 = _T_1503 | _T_1497; // @[Mux.scala 27:72]
  wire  _T_1489 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 418:132]
  wire  _T_1498 = _T_1489 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1504 | _T_1498; // @[Mux.scala 27:72]
  wire  _T_1507 = _T_1474 & _T_1505; // @[el2_ifu_mem_ctl.scala 418:69]
  wire  _T_1508 = _T_1470 | _T_1507; // @[el2_ifu_mem_ctl.scala 417:94]
  wire [4:0] _GEN_469 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 419:95]
  wire  _T_1511 = _GEN_469 == 5'h1f; // @[el2_ifu_mem_ctl.scala 419:95]
  wire  _T_1512 = bypass_valid_value_check & _T_1511; // @[el2_ifu_mem_ctl.scala 419:56]
  wire  bypass_data_ready_in = _T_1508 | _T_1512; // @[el2_ifu_mem_ctl.scala 418:181]
  wire  _T_1513 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 423:53]
  wire  _T_1514 = _T_1513 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 423:73]
  wire  _T_1516 = _T_1514 & _T_319; // @[el2_ifu_mem_ctl.scala 423:96]
  wire  _T_1518 = _T_1516 & _T_58; // @[el2_ifu_mem_ctl.scala 423:118]
  wire  _T_1520 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 424:73]
  wire  _T_1522 = _T_1520 & _T_319; // @[el2_ifu_mem_ctl.scala 424:96]
  wire  _T_1524 = _T_1522 & _T_58; // @[el2_ifu_mem_ctl.scala 424:118]
  wire  _T_1525 = _T_1518 | _T_1524; // @[el2_ifu_mem_ctl.scala 423:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 426:58]
  wire  _T_1526 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 425:54]
  wire  _T_1527 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 425:76]
  wire  _T_1528 = _T_1526 & _T_1527; // @[el2_ifu_mem_ctl.scala 425:74]
  wire  _T_1530 = _T_1528 & _T_319; // @[el2_ifu_mem_ctl.scala 425:96]
  wire  ic_crit_wd_rdy_new_in = _T_1525 | _T_1530; // @[el2_ifu_mem_ctl.scala 424:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 625:43]
  wire  _T_1251 = ic_crit_wd_rdy | _T_2235; // @[el2_ifu_mem_ctl.scala 371:38]
  wire  _T_1253 = _T_1251 | _T_2251; // @[el2_ifu_mem_ctl.scala 371:64]
  wire  _T_1254 = ~_T_1253; // @[el2_ifu_mem_ctl.scala 371:21]
  wire  _T_1255 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 371:98]
  wire  sel_ic_data = _T_1254 & _T_1255; // @[el2_ifu_mem_ctl.scala 371:96]
  wire  _T_2458 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 470:44]
  wire  _T_1624 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 437:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 409:60]
  wire  _T_1568 = _T_1415 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1418 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1568 | _T_1569; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1421 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1570; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1424 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1571; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1427 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1572; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1430 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1580 = _T_1579 | _T_1573; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1433 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1581 = _T_1580 | _T_1574; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1436 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1581 | _T_1575; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_2168 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1608 = _T_2171 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1615 = _T_1607 | _T_1608; // @[Mux.scala 27:72]
  wire  _T_1609 = _T_2174 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1616 = _T_1615 | _T_1609; // @[Mux.scala 27:72]
  wire  _T_1610 = _T_2177 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1617 = _T_1616 | _T_1610; // @[Mux.scala 27:72]
  wire  _T_1611 = _T_2180 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1618 = _T_1617 | _T_1611; // @[Mux.scala 27:72]
  wire  _T_1612 = _T_2183 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1619 = _T_1618 | _T_1612; // @[Mux.scala 27:72]
  wire  _T_1613 = _T_2186 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1620 = _T_1619 | _T_1613; // @[Mux.scala 27:72]
  wire  _T_1614 = _T_2189 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1620 | _T_1614; // @[Mux.scala 27:72]
  wire  _T_1625 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 439:70]
  wire  ifu_byp_data_err_new = _T_1624 ? ic_miss_buff_data_error_bypass : _T_1625; // @[el2_ifu_mem_ctl.scala 437:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 382:42]
  wire  _T_2459 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 470:91]
  wire  _T_2460 = ~_T_2459; // @[el2_ifu_mem_ctl.scala 470:60]
  wire  ic_rd_parity_final_err = _T_2458 & _T_2460; // @[el2_ifu_mem_ctl.scala 470:58]
  reg  ic_debug_ict_array_sel_ff; // @[el2_ifu_mem_ctl.scala 833:63]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9970 = _T_4763 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 760:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9972 = _T_4764 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10225 = _T_9970 | _T_9972; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9974 = _T_4765 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10226 = _T_10225 | _T_9974; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9976 = _T_4766 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10227 = _T_10226 | _T_9976; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9978 = _T_4767 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10228 = _T_10227 | _T_9978; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9980 = _T_4768 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10229 = _T_10228 | _T_9980; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9982 = _T_4769 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10230 = _T_10229 | _T_9982; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9984 = _T_4770 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10231 = _T_10230 | _T_9984; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9986 = _T_4771 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10232 = _T_10231 | _T_9986; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9988 = _T_4772 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10233 = _T_10232 | _T_9988; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9990 = _T_4773 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10234 = _T_10233 | _T_9990; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9992 = _T_4774 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10235 = _T_10234 | _T_9992; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9994 = _T_4775 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10236 = _T_10235 | _T_9994; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9996 = _T_4776 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10237 = _T_10236 | _T_9996; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9998 = _T_4777 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10238 = _T_10237 | _T_9998; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_10000 = _T_4778 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10239 = _T_10238 | _T_10000; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_10002 = _T_4779 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10240 = _T_10239 | _T_10002; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_10004 = _T_4780 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10241 = _T_10240 | _T_10004; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_10006 = _T_4781 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10242 = _T_10241 | _T_10006; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_10008 = _T_4782 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10243 = _T_10242 | _T_10008; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_10010 = _T_4783 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10244 = _T_10243 | _T_10010; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_10012 = _T_4784 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10245 = _T_10244 | _T_10012; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_10014 = _T_4785 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10246 = _T_10245 | _T_10014; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_10016 = _T_4786 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10247 = _T_10246 | _T_10016; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_10018 = _T_4787 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10248 = _T_10247 | _T_10018; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_10020 = _T_4788 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10249 = _T_10248 | _T_10020; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_10022 = _T_4789 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10250 = _T_10249 | _T_10022; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_10024 = _T_4790 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10251 = _T_10250 | _T_10024; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_10026 = _T_4791 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10252 = _T_10251 | _T_10026; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_10028 = _T_4792 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10253 = _T_10252 | _T_10028; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_10030 = _T_4793 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10254 = _T_10253 | _T_10030; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_10032 = _T_4794 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10255 = _T_10254 | _T_10032; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_10034 = _T_4795 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10256 = _T_10255 | _T_10034; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_10036 = _T_4796 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10257 = _T_10256 | _T_10036; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_10038 = _T_4797 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10258 = _T_10257 | _T_10038; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_10040 = _T_4798 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10259 = _T_10258 | _T_10040; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_10042 = _T_4799 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10260 = _T_10259 | _T_10042; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_10044 = _T_4800 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10261 = _T_10260 | _T_10044; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_10046 = _T_4801 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10262 = _T_10261 | _T_10046; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_10048 = _T_4802 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10263 = _T_10262 | _T_10048; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_10050 = _T_4803 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10264 = _T_10263 | _T_10050; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_10052 = _T_4804 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10265 = _T_10264 | _T_10052; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_10054 = _T_4805 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10266 = _T_10265 | _T_10054; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_10056 = _T_4806 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10267 = _T_10266 | _T_10056; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_10058 = _T_4807 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10268 = _T_10267 | _T_10058; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_10060 = _T_4808 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10269 = _T_10268 | _T_10060; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_10062 = _T_4809 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10270 = _T_10269 | _T_10062; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_10064 = _T_4810 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10271 = _T_10270 | _T_10064; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_10066 = _T_4811 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10272 = _T_10271 | _T_10066; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_10068 = _T_4812 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10273 = _T_10272 | _T_10068; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_10070 = _T_4813 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10274 = _T_10273 | _T_10070; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_10072 = _T_4814 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10275 = _T_10274 | _T_10072; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_10074 = _T_4815 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10276 = _T_10275 | _T_10074; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_10076 = _T_4816 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10277 = _T_10276 | _T_10076; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_10078 = _T_4817 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10278 = _T_10277 | _T_10078; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_10080 = _T_4818 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10279 = _T_10278 | _T_10080; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_10082 = _T_4819 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10280 = _T_10279 | _T_10082; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_10084 = _T_4820 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10281 = _T_10280 | _T_10084; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_10086 = _T_4821 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10282 = _T_10281 | _T_10086; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_10088 = _T_4822 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10283 = _T_10282 | _T_10088; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_10090 = _T_4823 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10284 = _T_10283 | _T_10090; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_10092 = _T_4824 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10285 = _T_10284 | _T_10092; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_10094 = _T_4825 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10286 = _T_10285 | _T_10094; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_10096 = _T_4826 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10287 = _T_10286 | _T_10096; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_10098 = _T_4827 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10288 = _T_10287 | _T_10098; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_10100 = _T_4828 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10289 = _T_10288 | _T_10100; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_10102 = _T_4829 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10290 = _T_10289 | _T_10102; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_10104 = _T_4830 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10291 = _T_10290 | _T_10104; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_10106 = _T_4831 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10292 = _T_10291 | _T_10106; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_10108 = _T_4832 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10293 = _T_10292 | _T_10108; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_10110 = _T_4833 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10294 = _T_10293 | _T_10110; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_10112 = _T_4834 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10295 = _T_10294 | _T_10112; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_10114 = _T_4835 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10296 = _T_10295 | _T_10114; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_10116 = _T_4836 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10297 = _T_10296 | _T_10116; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_10118 = _T_4837 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10298 = _T_10297 | _T_10118; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_10120 = _T_4838 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10299 = _T_10298 | _T_10120; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_10122 = _T_4839 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10300 = _T_10299 | _T_10122; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_10124 = _T_4840 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10301 = _T_10300 | _T_10124; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_10126 = _T_4841 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10302 = _T_10301 | _T_10126; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_10128 = _T_4842 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10303 = _T_10302 | _T_10128; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_10130 = _T_4843 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10304 = _T_10303 | _T_10130; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_10132 = _T_4844 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10305 = _T_10304 | _T_10132; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_10134 = _T_4845 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10306 = _T_10305 | _T_10134; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_10136 = _T_4846 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10307 = _T_10306 | _T_10136; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_10138 = _T_4847 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10308 = _T_10307 | _T_10138; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_10140 = _T_4848 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10309 = _T_10308 | _T_10140; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_10142 = _T_4849 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10310 = _T_10309 | _T_10142; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_10144 = _T_4850 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10311 = _T_10310 | _T_10144; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_10146 = _T_4851 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10312 = _T_10311 | _T_10146; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_10148 = _T_4852 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10313 = _T_10312 | _T_10148; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_10150 = _T_4853 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10314 = _T_10313 | _T_10150; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_10152 = _T_4854 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10315 = _T_10314 | _T_10152; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_10154 = _T_4855 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10316 = _T_10315 | _T_10154; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_10156 = _T_4856 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10317 = _T_10316 | _T_10156; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_10158 = _T_4857 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10318 = _T_10317 | _T_10158; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_10160 = _T_4858 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10319 = _T_10318 | _T_10160; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_10162 = _T_4859 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10320 = _T_10319 | _T_10162; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_10164 = _T_4860 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10321 = _T_10320 | _T_10164; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_10166 = _T_4861 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10322 = _T_10321 | _T_10166; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_10168 = _T_4862 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10323 = _T_10322 | _T_10168; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_10170 = _T_4863 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10324 = _T_10323 | _T_10170; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_10172 = _T_4864 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10325 = _T_10324 | _T_10172; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_10174 = _T_4865 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10326 = _T_10325 | _T_10174; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_10176 = _T_4866 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10327 = _T_10326 | _T_10176; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_10178 = _T_4867 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10328 = _T_10327 | _T_10178; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_10180 = _T_4868 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10329 = _T_10328 | _T_10180; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_10182 = _T_4869 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10330 = _T_10329 | _T_10182; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_10184 = _T_4870 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10331 = _T_10330 | _T_10184; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_10186 = _T_4871 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10332 = _T_10331 | _T_10186; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_10188 = _T_4872 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10333 = _T_10332 | _T_10188; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_10190 = _T_4873 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10334 = _T_10333 | _T_10190; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_10192 = _T_4874 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10335 = _T_10334 | _T_10192; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_10194 = _T_4875 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10336 = _T_10335 | _T_10194; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_10196 = _T_4876 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10337 = _T_10336 | _T_10196; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_10198 = _T_4877 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10338 = _T_10337 | _T_10198; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_10200 = _T_4878 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10339 = _T_10338 | _T_10200; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_10202 = _T_4879 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10340 = _T_10339 | _T_10202; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_10204 = _T_4880 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10341 = _T_10340 | _T_10204; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_10206 = _T_4881 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10342 = _T_10341 | _T_10206; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_10208 = _T_4882 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10343 = _T_10342 | _T_10208; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_10210 = _T_4883 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10344 = _T_10343 | _T_10210; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_10212 = _T_4884 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10345 = _T_10344 | _T_10212; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_10214 = _T_4885 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10346 = _T_10345 | _T_10214; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_10216 = _T_4886 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10347 = _T_10346 | _T_10216; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_10218 = _T_4887 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10348 = _T_10347 | _T_10218; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_10220 = _T_4888 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10349 = _T_10348 | _T_10220; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_10222 = _T_4889 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10350 = _T_10349 | _T_10222; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_10224 = _T_4890 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_10351 = _T_10350 | _T_10224; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9587 = _T_4763 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 760:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9589 = _T_4764 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9842 = _T_9587 | _T_9589; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9591 = _T_4765 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9843 = _T_9842 | _T_9591; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9593 = _T_4766 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9844 = _T_9843 | _T_9593; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9595 = _T_4767 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9845 = _T_9844 | _T_9595; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9597 = _T_4768 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9846 = _T_9845 | _T_9597; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9599 = _T_4769 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9847 = _T_9846 | _T_9599; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9601 = _T_4770 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9848 = _T_9847 | _T_9601; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9603 = _T_4771 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9849 = _T_9848 | _T_9603; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9605 = _T_4772 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9850 = _T_9849 | _T_9605; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9607 = _T_4773 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9851 = _T_9850 | _T_9607; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9609 = _T_4774 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9852 = _T_9851 | _T_9609; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9611 = _T_4775 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9853 = _T_9852 | _T_9611; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9613 = _T_4776 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9854 = _T_9853 | _T_9613; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9615 = _T_4777 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9855 = _T_9854 | _T_9615; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9617 = _T_4778 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9856 = _T_9855 | _T_9617; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9619 = _T_4779 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9857 = _T_9856 | _T_9619; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9621 = _T_4780 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9858 = _T_9857 | _T_9621; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9623 = _T_4781 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9859 = _T_9858 | _T_9623; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9625 = _T_4782 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9860 = _T_9859 | _T_9625; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9627 = _T_4783 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9861 = _T_9860 | _T_9627; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9629 = _T_4784 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9862 = _T_9861 | _T_9629; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9631 = _T_4785 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9863 = _T_9862 | _T_9631; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9633 = _T_4786 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9864 = _T_9863 | _T_9633; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9635 = _T_4787 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9865 = _T_9864 | _T_9635; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9637 = _T_4788 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9866 = _T_9865 | _T_9637; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9639 = _T_4789 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9867 = _T_9866 | _T_9639; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9641 = _T_4790 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9868 = _T_9867 | _T_9641; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9643 = _T_4791 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9869 = _T_9868 | _T_9643; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9645 = _T_4792 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9870 = _T_9869 | _T_9645; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9647 = _T_4793 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9871 = _T_9870 | _T_9647; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9649 = _T_4794 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9872 = _T_9871 | _T_9649; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9651 = _T_4795 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9873 = _T_9872 | _T_9651; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9653 = _T_4796 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9874 = _T_9873 | _T_9653; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9655 = _T_4797 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9875 = _T_9874 | _T_9655; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9657 = _T_4798 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9876 = _T_9875 | _T_9657; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9659 = _T_4799 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9877 = _T_9876 | _T_9659; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9661 = _T_4800 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9878 = _T_9877 | _T_9661; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9663 = _T_4801 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9879 = _T_9878 | _T_9663; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9665 = _T_4802 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9880 = _T_9879 | _T_9665; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9667 = _T_4803 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9881 = _T_9880 | _T_9667; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9669 = _T_4804 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9882 = _T_9881 | _T_9669; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9671 = _T_4805 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9883 = _T_9882 | _T_9671; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9673 = _T_4806 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9884 = _T_9883 | _T_9673; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9675 = _T_4807 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9885 = _T_9884 | _T_9675; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9677 = _T_4808 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9886 = _T_9885 | _T_9677; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9679 = _T_4809 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9887 = _T_9886 | _T_9679; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9681 = _T_4810 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9888 = _T_9887 | _T_9681; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9683 = _T_4811 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9889 = _T_9888 | _T_9683; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9685 = _T_4812 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9890 = _T_9889 | _T_9685; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9687 = _T_4813 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9891 = _T_9890 | _T_9687; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9689 = _T_4814 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9892 = _T_9891 | _T_9689; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9691 = _T_4815 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9893 = _T_9892 | _T_9691; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9693 = _T_4816 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9894 = _T_9893 | _T_9693; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9695 = _T_4817 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9895 = _T_9894 | _T_9695; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9697 = _T_4818 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9896 = _T_9895 | _T_9697; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9699 = _T_4819 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9897 = _T_9896 | _T_9699; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9701 = _T_4820 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9898 = _T_9897 | _T_9701; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9703 = _T_4821 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9899 = _T_9898 | _T_9703; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9705 = _T_4822 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9900 = _T_9899 | _T_9705; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9707 = _T_4823 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9901 = _T_9900 | _T_9707; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9709 = _T_4824 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9902 = _T_9901 | _T_9709; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9711 = _T_4825 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9903 = _T_9902 | _T_9711; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9713 = _T_4826 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9904 = _T_9903 | _T_9713; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9715 = _T_4827 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9905 = _T_9904 | _T_9715; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9717 = _T_4828 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9906 = _T_9905 | _T_9717; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9719 = _T_4829 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9907 = _T_9906 | _T_9719; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9721 = _T_4830 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9908 = _T_9907 | _T_9721; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9723 = _T_4831 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9909 = _T_9908 | _T_9723; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9725 = _T_4832 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9910 = _T_9909 | _T_9725; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9727 = _T_4833 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9911 = _T_9910 | _T_9727; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9729 = _T_4834 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9912 = _T_9911 | _T_9729; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9731 = _T_4835 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9913 = _T_9912 | _T_9731; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9733 = _T_4836 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9914 = _T_9913 | _T_9733; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9735 = _T_4837 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9915 = _T_9914 | _T_9735; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9737 = _T_4838 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9916 = _T_9915 | _T_9737; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9739 = _T_4839 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9917 = _T_9916 | _T_9739; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9741 = _T_4840 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9918 = _T_9917 | _T_9741; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9743 = _T_4841 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9919 = _T_9918 | _T_9743; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9745 = _T_4842 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9920 = _T_9919 | _T_9745; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9747 = _T_4843 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9921 = _T_9920 | _T_9747; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9749 = _T_4844 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9922 = _T_9921 | _T_9749; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9751 = _T_4845 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9923 = _T_9922 | _T_9751; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9753 = _T_4846 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9924 = _T_9923 | _T_9753; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9755 = _T_4847 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9925 = _T_9924 | _T_9755; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9757 = _T_4848 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9926 = _T_9925 | _T_9757; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9759 = _T_4849 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9927 = _T_9926 | _T_9759; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9761 = _T_4850 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9928 = _T_9927 | _T_9761; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9763 = _T_4851 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9929 = _T_9928 | _T_9763; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9765 = _T_4852 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9930 = _T_9929 | _T_9765; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9767 = _T_4853 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9931 = _T_9930 | _T_9767; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9769 = _T_4854 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9932 = _T_9931 | _T_9769; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9771 = _T_4855 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9933 = _T_9932 | _T_9771; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9773 = _T_4856 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9934 = _T_9933 | _T_9773; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9775 = _T_4857 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9935 = _T_9934 | _T_9775; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9777 = _T_4858 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9936 = _T_9935 | _T_9777; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9779 = _T_4859 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9937 = _T_9936 | _T_9779; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9781 = _T_4860 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9938 = _T_9937 | _T_9781; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9783 = _T_4861 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9939 = _T_9938 | _T_9783; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9785 = _T_4862 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9940 = _T_9939 | _T_9785; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9787 = _T_4863 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9941 = _T_9940 | _T_9787; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9789 = _T_4864 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9942 = _T_9941 | _T_9789; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9791 = _T_4865 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9943 = _T_9942 | _T_9791; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9793 = _T_4866 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9944 = _T_9943 | _T_9793; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9795 = _T_4867 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9945 = _T_9944 | _T_9795; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9797 = _T_4868 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9946 = _T_9945 | _T_9797; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9799 = _T_4869 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9947 = _T_9946 | _T_9799; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9801 = _T_4870 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9948 = _T_9947 | _T_9801; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9803 = _T_4871 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9949 = _T_9948 | _T_9803; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9805 = _T_4872 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9950 = _T_9949 | _T_9805; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9807 = _T_4873 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9951 = _T_9950 | _T_9807; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9809 = _T_4874 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9952 = _T_9951 | _T_9809; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9811 = _T_4875 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9953 = _T_9952 | _T_9811; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9813 = _T_4876 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9954 = _T_9953 | _T_9813; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9815 = _T_4877 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9955 = _T_9954 | _T_9815; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9817 = _T_4878 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9956 = _T_9955 | _T_9817; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9819 = _T_4879 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9957 = _T_9956 | _T_9819; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9821 = _T_4880 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9958 = _T_9957 | _T_9821; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9823 = _T_4881 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9959 = _T_9958 | _T_9823; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9825 = _T_4882 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9960 = _T_9959 | _T_9825; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9827 = _T_4883 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9961 = _T_9960 | _T_9827; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9829 = _T_4884 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9962 = _T_9961 | _T_9829; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9831 = _T_4885 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9963 = _T_9962 | _T_9831; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9833 = _T_4886 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9964 = _T_9963 | _T_9833; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9835 = _T_4887 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9965 = _T_9964 | _T_9835; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9837 = _T_4888 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9966 = _T_9965 | _T_9837; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9839 = _T_4889 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9967 = _T_9966 | _T_9839; // @[el2_ifu_mem_ctl.scala 760:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9841 = _T_4890 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 760:10]
  wire  _T_9968 = _T_9967 | _T_9841; // @[el2_ifu_mem_ctl.scala 760:91]
  wire [1:0] ic_tag_valid_unq = {_T_10351,_T_9968}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[el2_ifu_mem_ctl.scala 832:53]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 834:54]
  wire [1:0] _T_10391 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10392 = ic_debug_way_ff & _T_10391; // @[el2_ifu_mem_ctl.scala 815:67]
  wire [1:0] _T_10393 = ic_tag_valid_unq & _T_10392; // @[el2_ifu_mem_ctl.scala 815:48]
  wire  ic_debug_tag_val_rd_out = |_T_10393; // @[el2_ifu_mem_ctl.scala 815:115]
  wire [65:0] _T_1210 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1211; // @[el2_ifu_mem_ctl.scala 354:63]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2593; // @[el2_ifu_mem_ctl.scala 365:80]
  wire  _T_1249 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 370:98]
  wire  sel_byp_data = _T_1253 & _T_1249; // @[el2_ifu_mem_ctl.scala 370:96]
  wire [63:0] _T_1260 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1261 = _T_1260 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 377:69]
  wire [63:0] _T_1263 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2115 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 445:31]
  wire  _T_1628 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 441:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1629 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1677 = _T_1629 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1632 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1678 = _T_1632 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1677 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1635 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1679 = _T_1635 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire  _T_1638 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1680 = _T_1638 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1695 = _T_1694 | _T_1680; // @[Mux.scala 27:72]
  wire  _T_1641 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1681 = _T_1641 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1696 = _T_1695 | _T_1681; // @[Mux.scala 27:72]
  wire  _T_1644 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1682 = _T_1644 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1697 = _T_1696 | _T_1682; // @[Mux.scala 27:72]
  wire  _T_1647 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1683 = _T_1647 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1698 = _T_1697 | _T_1683; // @[Mux.scala 27:72]
  wire  _T_1650 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1684 = _T_1650 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1699 = _T_1698 | _T_1684; // @[Mux.scala 27:72]
  wire  _T_1653 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1685 = _T_1653 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1700 = _T_1699 | _T_1685; // @[Mux.scala 27:72]
  wire  _T_1656 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1686 = _T_1656 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1701 = _T_1700 | _T_1686; // @[Mux.scala 27:72]
  wire  _T_1659 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1687 = _T_1659 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1702 = _T_1701 | _T_1687; // @[Mux.scala 27:72]
  wire  _T_1662 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1688 = _T_1662 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1703 = _T_1702 | _T_1688; // @[Mux.scala 27:72]
  wire  _T_1665 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1689 = _T_1665 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1704 = _T_1703 | _T_1689; // @[Mux.scala 27:72]
  wire  _T_1668 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1690 = _T_1668 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1705 = _T_1704 | _T_1690; // @[Mux.scala 27:72]
  wire  _T_1671 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1691 = _T_1671 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1706 = _T_1705 | _T_1691; // @[Mux.scala 27:72]
  wire  _T_1674 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1692 = _T_1674 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1707 = _T_1706 | _T_1692; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1709 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1757 = _T_1709 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1712 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1758 = _T_1712 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1757 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1715 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1759 = _T_1715 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1718 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1760 = _T_1718 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1775 = _T_1774 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1721 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1761 = _T_1721 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1776 = _T_1775 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1724 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1762 = _T_1724 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1777 = _T_1776 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1727 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1763 = _T_1727 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1778 = _T_1777 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1730 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1764 = _T_1730 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1779 = _T_1778 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1733 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1765 = _T_1733 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1780 = _T_1779 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1736 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1766 = _T_1736 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1781 = _T_1780 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1739 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1767 = _T_1739 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1782 = _T_1781 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1742 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1768 = _T_1742 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1783 = _T_1782 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1745 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1769 = _T_1745 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1784 = _T_1783 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1748 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1770 = _T_1748 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1785 = _T_1784 | _T_1770; // @[Mux.scala 27:72]
  wire  _T_1751 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1771 = _T_1751 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1786 = _T_1785 | _T_1771; // @[Mux.scala 27:72]
  wire  _T_1754 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:179]
  wire [31:0] _T_1772 = _T_1754 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1787 = _T_1786 | _T_1772; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1789 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1837 = _T_1789 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1792 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1838 = _T_1792 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1837 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1795 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1839 = _T_1795 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire  _T_1798 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1840 = _T_1798 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1855 = _T_1854 | _T_1840; // @[Mux.scala 27:72]
  wire  _T_1801 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1841 = _T_1801 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1856 = _T_1855 | _T_1841; // @[Mux.scala 27:72]
  wire  _T_1804 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1842 = _T_1804 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1857 = _T_1856 | _T_1842; // @[Mux.scala 27:72]
  wire  _T_1807 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1843 = _T_1807 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1858 = _T_1857 | _T_1843; // @[Mux.scala 27:72]
  wire  _T_1810 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1844 = _T_1810 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1859 = _T_1858 | _T_1844; // @[Mux.scala 27:72]
  wire  _T_1813 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1845 = _T_1813 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1860 = _T_1859 | _T_1845; // @[Mux.scala 27:72]
  wire  _T_1816 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1846 = _T_1816 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1861 = _T_1860 | _T_1846; // @[Mux.scala 27:72]
  wire  _T_1819 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1847 = _T_1819 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1862 = _T_1861 | _T_1847; // @[Mux.scala 27:72]
  wire  _T_1822 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1848 = _T_1822 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1863 = _T_1862 | _T_1848; // @[Mux.scala 27:72]
  wire  _T_1825 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1849 = _T_1825 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1864 = _T_1863 | _T_1849; // @[Mux.scala 27:72]
  wire  _T_1828 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1850 = _T_1828 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1865 = _T_1864 | _T_1850; // @[Mux.scala 27:72]
  wire  _T_1831 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1851 = _T_1831 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1866 = _T_1865 | _T_1851; // @[Mux.scala 27:72]
  wire  _T_1834 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:285]
  wire [31:0] _T_1852 = _T_1834 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1867 = _T_1866 | _T_1852; // @[Mux.scala 27:72]
  wire [79:0] _T_1870 = {_T_1707,_T_1787,_T_1867}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1871 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1919 = _T_1871 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1874 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1920 = _T_1874 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1919 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1877 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1921 = _T_1877 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire  _T_1880 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1922 = _T_1880 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1937 = _T_1936 | _T_1922; // @[Mux.scala 27:72]
  wire  _T_1883 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1923 = _T_1883 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1938 = _T_1937 | _T_1923; // @[Mux.scala 27:72]
  wire  _T_1886 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1924 = _T_1886 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1939 = _T_1938 | _T_1924; // @[Mux.scala 27:72]
  wire  _T_1889 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1925 = _T_1889 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1940 = _T_1939 | _T_1925; // @[Mux.scala 27:72]
  wire  _T_1892 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1926 = _T_1892 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1941 = _T_1940 | _T_1926; // @[Mux.scala 27:72]
  wire  _T_1895 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1927 = _T_1895 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1942 = _T_1941 | _T_1927; // @[Mux.scala 27:72]
  wire  _T_1898 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1928 = _T_1898 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1943 = _T_1942 | _T_1928; // @[Mux.scala 27:72]
  wire  _T_1901 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1929 = _T_1901 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1944 = _T_1943 | _T_1929; // @[Mux.scala 27:72]
  wire  _T_1904 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1930 = _T_1904 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1945 = _T_1944 | _T_1930; // @[Mux.scala 27:72]
  wire  _T_1907 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1931 = _T_1907 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1946 = _T_1945 | _T_1931; // @[Mux.scala 27:72]
  wire  _T_1910 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1932 = _T_1910 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1947 = _T_1946 | _T_1932; // @[Mux.scala 27:72]
  wire  _T_1913 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1933 = _T_1913 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1948 = _T_1947 | _T_1933; // @[Mux.scala 27:72]
  wire  _T_1916 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 443:73]
  wire [15:0] _T_1934 = _T_1916 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1949 = _T_1948 | _T_1934; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1629 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1632 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_1999 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1635 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1638 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2017 = _T_2016 | _T_2002; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_1641 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2018 = _T_2017 | _T_2003; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_1644 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2019 = _T_2018 | _T_2004; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_1647 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2020 = _T_2019 | _T_2005; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_1650 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2021 = _T_2020 | _T_2006; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_1653 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2022 = _T_2021 | _T_2007; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_1656 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2023 = _T_2022 | _T_2008; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_1659 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2024 = _T_2023 | _T_2009; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_1662 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2025 = _T_2024 | _T_2010; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_1665 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2026 = _T_2025 | _T_2011; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_1668 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2027 = _T_2026 | _T_2012; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_1671 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2028 = _T_2027 | _T_2013; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_1674 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2029 = _T_2028 | _T_2014; // @[Mux.scala 27:72]
  wire [79:0] _T_2112 = {_T_1949,_T_2029,_T_1787}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1628 ? _T_1870 : _T_2112; // @[el2_ifu_mem_ctl.scala 441:37]
  wire [79:0] _T_2117 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2115 ? ic_byp_data_only_pre_new : _T_2117; // @[el2_ifu_mem_ctl.scala 445:30]
  wire [79:0] _GEN_470 = {{16'd0}, _T_1263}; // @[el2_ifu_mem_ctl.scala 377:114]
  wire [79:0] _T_1264 = _GEN_470 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 377:114]
  wire [79:0] _GEN_471 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 377:88]
  wire [79:0] ic_premux_data_temp = _GEN_471 | _T_1264; // @[el2_ifu_mem_ctl.scala 377:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_319; // @[el2_ifu_mem_ctl.scala 384:38]
  wire [1:0] _T_1273 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 388:8]
  wire  _T_1275 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 390:45]
  wire  _T_1277 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 390:80]
  wire  _T_1278 = ~_T_1277; // @[el2_ifu_mem_ctl.scala 390:71]
  wire  _T_1279 = _T_1275 & _T_1278; // @[el2_ifu_mem_ctl.scala 390:69]
  wire  _T_1280 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 390:131]
  wire  _T_1281 = _T_1279 & _T_1280; // @[el2_ifu_mem_ctl.scala 390:114]
  wire [7:0] _T_1370 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1375 = ic_miss_buff_data_error[0] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  _T_2656 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 621:47]
  wire  _T_2657 = _T_2656 & _T_13; // @[el2_ifu_mem_ctl.scala 621:50]
  wire  bus_ifu_wr_data_error = _T_2657 & miss_pending; // @[el2_ifu_mem_ctl.scala 621:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1375; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1379 = ic_miss_buff_data_error[1] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1379; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1383 = ic_miss_buff_data_error[2] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1383; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1387 = ic_miss_buff_data_error[3] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1387; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1391 = ic_miss_buff_data_error[4] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1391; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1395 = ic_miss_buff_data_error[5] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1395; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1399 = ic_miss_buff_data_error[6] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1399; // @[el2_ifu_mem_ctl.scala 407:72]
  wire  _T_1403 = ic_miss_buff_data_error[7] & _T_1341; // @[el2_ifu_mem_ctl.scala 408:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1403; // @[el2_ifu_mem_ctl.scala 407:72]
  wire [7:0] _T_1410 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2467 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2475 = _T_6 & _T_319; // @[el2_ifu_mem_ctl.scala 490:65]
  wire  _T_2476 = _T_2475 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 490:88]
  wire  _T_2478 = _T_2476 & _T_2589; // @[el2_ifu_mem_ctl.scala 490:112]
  wire  _T_2479 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2480 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 495:50]
  wire  _T_2482 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2488 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2490 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2488 | _T_2490; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2482 ? _T_2480 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2479 ? _T_2480 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2467 ? _T_2478 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2467 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2481 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 496:56]
  wire  _GEN_43 = _T_2479 & _T_2481; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2467 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 481:58]
  wire  _T_2464 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 480:49]
  wire  _T_2469 = io_ic_error_start & _T_319; // @[el2_ifu_mem_ctl.scala 489:87]
  wire  _T_2483 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 499:54]
  wire  _T_2484 = _T_2483 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 499:84]
  wire  _T_2493 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 520:66]
  wire  _T_2494 = io_dec_tlu_flush_err_wb & _T_2493; // @[el2_ifu_mem_ctl.scala 520:52]
  wire  _T_2496 = _T_2494 & _T_2589; // @[el2_ifu_mem_ctl.scala 520:81]
  wire  _T_2498 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 523:59]
  wire  _T_2499 = _T_2498 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 523:86]
  wire  _T_2513 = _T_2498 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 526:81]
  wire  _T_2514 = _T_2513 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 526:103]
  wire  _T_2515 = _T_2514 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 526:126]
  wire  _T_2535 = _T_2513 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 533:103]
  wire  _T_2542 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 538:62]
  wire  _T_2543 = io_dec_tlu_flush_lower_wb & _T_2542; // @[el2_ifu_mem_ctl.scala 538:60]
  wire  _T_2544 = _T_2543 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 538:88]
  wire  _T_2545 = _T_2544 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 538:115]
  wire  _GEN_50 = _T_2541 & _T_2499; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_2524 ? _T_2535 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_2524 | _T_2541; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_2497 ? _T_2515 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2497 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2492 ? _T_2496 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2557 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 555:64]
  wire  _T_2559 = _T_2557 & _T_2589; // @[el2_ifu_mem_ctl.scala 555:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2561 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 555:133]
  wire  _T_2562 = _T_2561 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 555:164]
  wire  _T_2563 = _T_2562 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 555:184]
  wire  _T_2564 = _T_2563 & miss_pending; // @[el2_ifu_mem_ctl.scala 555:204]
  wire  _T_2565 = ~_T_2564; // @[el2_ifu_mem_ctl.scala 555:112]
  wire  ifc_bus_ic_req_ff_in = _T_2559 & _T_2565; // @[el2_ifu_mem_ctl.scala 555:110]
  wire  _T_2566 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 556:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 587:45]
  wire  _T_2583 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 590:35]
  wire  _T_2584 = _T_2583 & miss_pending; // @[el2_ifu_mem_ctl.scala 590:53]
  wire  bus_cmd_sent = _T_2584 & _T_2589; // @[el2_ifu_mem_ctl.scala 590:68]
  wire [2:0] _T_2574 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2576 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2578 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 588:51]
  wire  _T_2604 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 598:73]
  wire  _T_2605 = _T_2590 & _T_2604; // @[el2_ifu_mem_ctl.scala 598:71]
  wire  _T_2607 = last_data_recieved_ff & _T_1341; // @[el2_ifu_mem_ctl.scala 598:114]
  wire  last_data_recieved_in = _T_2605 | _T_2607; // @[el2_ifu_mem_ctl.scala 598:89]
  wire [2:0] _T_2613 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 603:45]
  wire  _T_2617 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 606:48]
  wire  _T_2618 = _T_2617 & miss_pending; // @[el2_ifu_mem_ctl.scala 606:68]
  wire  bus_inc_cmd_beat_cnt = _T_2618 & _T_2589; // @[el2_ifu_mem_ctl.scala 606:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 608:57]
  wire  _T_2622 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 609:31]
  wire  _T_2623 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 609:71]
  wire  _T_2624 = _T_2623 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 609:87]
  wire  _T_2625 = ~_T_2624; // @[el2_ifu_mem_ctl.scala 609:55]
  wire  bus_hold_cmd_beat_cnt = _T_2622 & _T_2625; // @[el2_ifu_mem_ctl.scala 609:53]
  wire  _T_2626 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 610:46]
  wire  bus_cmd_beat_en = _T_2626 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 610:62]
  wire [2:0] _T_2629 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 612:46]
  wire [2:0] _T_2631 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2632 = bus_inc_cmd_beat_cnt ? _T_2629 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2633 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2635 = _T_2631 | _T_2632; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2635 | _T_2633; // @[Mux.scala 27:72]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 624:62]
  wire  _T_2664 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 629:50]
  wire  _T_2665 = io_ifc_dma_access_ok & _T_2664; // @[el2_ifu_mem_ctl.scala 629:47]
  wire  _T_2666 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 629:70]
  wire  ifc_dma_access_ok_d = _T_2665 & _T_2666; // @[el2_ifu_mem_ctl.scala 629:68]
  wire  _T_2670 = _T_2665 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 630:72]
  wire  _T_2671 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 630:111]
  wire  _T_2672 = _T_2670 & _T_2671; // @[el2_ifu_mem_ctl.scala 630:97]
  wire  ifc_dma_access_q_ok = _T_2672 & _T_2666; // @[el2_ifu_mem_ctl.scala 630:127]
  wire  _T_2675 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 633:40]
  wire  _T_2676 = _T_2675 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 633:58]
  wire  _T_2679 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 634:60]
  wire  _T_2680 = _T_2675 & _T_2679; // @[el2_ifu_mem_ctl.scala 634:58]
  wire  _T_2681 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 634:104]
  wire [2:0] _T_2686 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2707 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[33]; // @[el2_lib.scala 237:74]
  wire  _T_2708 = _T_2707 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 237:74]
  wire  _T_2709 = _T_2708 ^ io_dma_mem_wdata[36]; // @[el2_lib.scala 237:74]
  wire  _T_2710 = _T_2709 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 237:74]
  wire  _T_2711 = _T_2710 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 237:74]
  wire  _T_2712 = _T_2711 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 237:74]
  wire  _T_2713 = _T_2712 ^ io_dma_mem_wdata[43]; // @[el2_lib.scala 237:74]
  wire  _T_2714 = _T_2713 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 237:74]
  wire  _T_2715 = _T_2714 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 237:74]
  wire  _T_2716 = _T_2715 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 237:74]
  wire  _T_2717 = _T_2716 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 237:74]
  wire  _T_2718 = _T_2717 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 237:74]
  wire  _T_2719 = _T_2718 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 237:74]
  wire  _T_2720 = _T_2719 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 237:74]
  wire  _T_2721 = _T_2720 ^ io_dma_mem_wdata[58]; // @[el2_lib.scala 237:74]
  wire  _T_2722 = _T_2721 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 237:74]
  wire  _T_2723 = _T_2722 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 237:74]
  wire  _T_2742 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 237:74]
  wire  _T_2743 = _T_2742 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 237:74]
  wire  _T_2744 = _T_2743 ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 237:74]
  wire  _T_2745 = _T_2744 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 237:74]
  wire  _T_2746 = _T_2745 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 237:74]
  wire  _T_2747 = _T_2746 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 237:74]
  wire  _T_2748 = _T_2747 ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 237:74]
  wire  _T_2749 = _T_2748 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 237:74]
  wire  _T_2750 = _T_2749 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 237:74]
  wire  _T_2751 = _T_2750 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 237:74]
  wire  _T_2752 = _T_2751 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 237:74]
  wire  _T_2753 = _T_2752 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 237:74]
  wire  _T_2754 = _T_2753 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 237:74]
  wire  _T_2755 = _T_2754 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 237:74]
  wire  _T_2756 = _T_2755 ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 237:74]
  wire  _T_2757 = _T_2756 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 237:74]
  wire  _T_2758 = _T_2757 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 237:74]
  wire  _T_2777 = io_dma_mem_wdata[33] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 237:74]
  wire  _T_2778 = _T_2777 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 237:74]
  wire  _T_2779 = _T_2778 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 237:74]
  wire  _T_2780 = _T_2779 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 237:74]
  wire  _T_2781 = _T_2780 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 237:74]
  wire  _T_2782 = _T_2781 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 237:74]
  wire  _T_2783 = _T_2782 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 237:74]
  wire  _T_2784 = _T_2783 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 237:74]
  wire  _T_2785 = _T_2784 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 237:74]
  wire  _T_2786 = _T_2785 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 237:74]
  wire  _T_2787 = _T_2786 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 237:74]
  wire  _T_2788 = _T_2787 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 237:74]
  wire  _T_2789 = _T_2788 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 237:74]
  wire  _T_2790 = _T_2789 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 237:74]
  wire  _T_2791 = _T_2790 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 237:74]
  wire  _T_2792 = _T_2791 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 237:74]
  wire  _T_2793 = _T_2792 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 237:74]
  wire  _T_2809 = io_dma_mem_wdata[36] ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 237:74]
  wire  _T_2810 = _T_2809 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 237:74]
  wire  _T_2811 = _T_2810 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 237:74]
  wire  _T_2812 = _T_2811 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 237:74]
  wire  _T_2813 = _T_2812 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 237:74]
  wire  _T_2814 = _T_2813 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 237:74]
  wire  _T_2815 = _T_2814 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 237:74]
  wire  _T_2816 = _T_2815 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 237:74]
  wire  _T_2817 = _T_2816 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 237:74]
  wire  _T_2818 = _T_2817 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 237:74]
  wire  _T_2819 = _T_2818 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 237:74]
  wire  _T_2820 = _T_2819 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 237:74]
  wire  _T_2821 = _T_2820 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 237:74]
  wire  _T_2822 = _T_2821 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 237:74]
  wire  _T_2838 = io_dma_mem_wdata[43] ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 237:74]
  wire  _T_2839 = _T_2838 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 237:74]
  wire  _T_2840 = _T_2839 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 237:74]
  wire  _T_2841 = _T_2840 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 237:74]
  wire  _T_2842 = _T_2841 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 237:74]
  wire  _T_2843 = _T_2842 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 237:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 237:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 237:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 237:74]
  wire  _T_2847 = _T_2846 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 237:74]
  wire  _T_2848 = _T_2847 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 237:74]
  wire  _T_2849 = _T_2848 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 237:74]
  wire  _T_2850 = _T_2849 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 237:74]
  wire  _T_2851 = _T_2850 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 237:74]
  wire  _T_2858 = io_dma_mem_wdata[58] ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 237:74]
  wire  _T_2859 = _T_2858 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 237:74]
  wire  _T_2860 = _T_2859 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 237:74]
  wire  _T_2861 = _T_2860 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 237:74]
  wire  _T_2862 = _T_2861 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 237:74]
  wire [5:0] _T_2867 = {_T_2862,_T_2851,_T_2822,_T_2793,_T_2758,_T_2723}; // @[Cat.scala 29:58]
  wire  _T_2868 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 245:13]
  wire  _T_2869 = ^_T_2867; // @[el2_lib.scala 245:23]
  wire  _T_2870 = _T_2868 ^ _T_2869; // @[el2_lib.scala 245:18]
  wire  _T_2891 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[1]; // @[el2_lib.scala 237:74]
  wire  _T_2892 = _T_2891 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 237:74]
  wire  _T_2893 = _T_2892 ^ io_dma_mem_wdata[4]; // @[el2_lib.scala 237:74]
  wire  _T_2894 = _T_2893 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 237:74]
  wire  _T_2895 = _T_2894 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 237:74]
  wire  _T_2896 = _T_2895 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 237:74]
  wire  _T_2897 = _T_2896 ^ io_dma_mem_wdata[11]; // @[el2_lib.scala 237:74]
  wire  _T_2898 = _T_2897 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 237:74]
  wire  _T_2899 = _T_2898 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 237:74]
  wire  _T_2900 = _T_2899 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 237:74]
  wire  _T_2901 = _T_2900 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 237:74]
  wire  _T_2902 = _T_2901 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 237:74]
  wire  _T_2903 = _T_2902 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 237:74]
  wire  _T_2904 = _T_2903 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 237:74]
  wire  _T_2905 = _T_2904 ^ io_dma_mem_wdata[26]; // @[el2_lib.scala 237:74]
  wire  _T_2906 = _T_2905 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 237:74]
  wire  _T_2907 = _T_2906 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 237:74]
  wire  _T_2926 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 237:74]
  wire  _T_2927 = _T_2926 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 237:74]
  wire  _T_2928 = _T_2927 ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 237:74]
  wire  _T_2929 = _T_2928 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 237:74]
  wire  _T_2930 = _T_2929 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 237:74]
  wire  _T_2931 = _T_2930 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 237:74]
  wire  _T_2932 = _T_2931 ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 237:74]
  wire  _T_2933 = _T_2932 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 237:74]
  wire  _T_2934 = _T_2933 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 237:74]
  wire  _T_2935 = _T_2934 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 237:74]
  wire  _T_2936 = _T_2935 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 237:74]
  wire  _T_2937 = _T_2936 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 237:74]
  wire  _T_2938 = _T_2937 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 237:74]
  wire  _T_2939 = _T_2938 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 237:74]
  wire  _T_2940 = _T_2939 ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 237:74]
  wire  _T_2941 = _T_2940 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 237:74]
  wire  _T_2942 = _T_2941 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 237:74]
  wire  _T_2961 = io_dma_mem_wdata[1] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 237:74]
  wire  _T_2962 = _T_2961 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 237:74]
  wire  _T_2963 = _T_2962 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 237:74]
  wire  _T_2964 = _T_2963 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 237:74]
  wire  _T_2965 = _T_2964 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 237:74]
  wire  _T_2966 = _T_2965 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 237:74]
  wire  _T_2967 = _T_2966 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 237:74]
  wire  _T_2968 = _T_2967 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 237:74]
  wire  _T_2969 = _T_2968 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 237:74]
  wire  _T_2970 = _T_2969 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 237:74]
  wire  _T_2971 = _T_2970 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 237:74]
  wire  _T_2972 = _T_2971 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 237:74]
  wire  _T_2973 = _T_2972 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 237:74]
  wire  _T_2974 = _T_2973 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 237:74]
  wire  _T_2975 = _T_2974 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 237:74]
  wire  _T_2976 = _T_2975 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 237:74]
  wire  _T_2977 = _T_2976 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 237:74]
  wire  _T_2993 = io_dma_mem_wdata[4] ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 237:74]
  wire  _T_2994 = _T_2993 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 237:74]
  wire  _T_2995 = _T_2994 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 237:74]
  wire  _T_2996 = _T_2995 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 237:74]
  wire  _T_2997 = _T_2996 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 237:74]
  wire  _T_2998 = _T_2997 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 237:74]
  wire  _T_2999 = _T_2998 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 237:74]
  wire  _T_3000 = _T_2999 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 237:74]
  wire  _T_3001 = _T_3000 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 237:74]
  wire  _T_3002 = _T_3001 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 237:74]
  wire  _T_3003 = _T_3002 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 237:74]
  wire  _T_3004 = _T_3003 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 237:74]
  wire  _T_3005 = _T_3004 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 237:74]
  wire  _T_3006 = _T_3005 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 237:74]
  wire  _T_3022 = io_dma_mem_wdata[11] ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 237:74]
  wire  _T_3023 = _T_3022 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 237:74]
  wire  _T_3024 = _T_3023 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 237:74]
  wire  _T_3025 = _T_3024 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 237:74]
  wire  _T_3026 = _T_3025 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 237:74]
  wire  _T_3027 = _T_3026 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 237:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 237:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 237:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 237:74]
  wire  _T_3031 = _T_3030 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 237:74]
  wire  _T_3032 = _T_3031 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 237:74]
  wire  _T_3033 = _T_3032 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 237:74]
  wire  _T_3034 = _T_3033 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 237:74]
  wire  _T_3035 = _T_3034 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 237:74]
  wire  _T_3042 = io_dma_mem_wdata[26] ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 237:74]
  wire  _T_3043 = _T_3042 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 237:74]
  wire  _T_3044 = _T_3043 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 237:74]
  wire  _T_3045 = _T_3044 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 237:74]
  wire  _T_3046 = _T_3045 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 237:74]
  wire [5:0] _T_3051 = {_T_3046,_T_3035,_T_3006,_T_2977,_T_2942,_T_2907}; // @[Cat.scala 29:58]
  wire  _T_3052 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 245:13]
  wire  _T_3053 = ^_T_3051; // @[el2_lib.scala 245:23]
  wire  _T_3054 = _T_3052 ^ _T_3053; // @[el2_lib.scala 245:18]
  wire [6:0] _T_3055 = {_T_3054,_T_3046,_T_3035,_T_3006,_T_2977,_T_2942,_T_2907}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2870,_T_2862,_T_2851,_T_2822,_T_2793,_T_2758,_T_2723,_T_3055}; // @[Cat.scala 29:58]
  wire  _T_3057 = ~_T_2675; // @[el2_ifu_mem_ctl.scala 640:45]
  wire  _T_3058 = iccm_correct_ecc & _T_3057; // @[el2_ifu_mem_ctl.scala 640:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3059 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3066 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 654:53]
  wire  _T_3399 = _T_3311[5:0] == 6'h27; // @[el2_lib.scala 317:41]
  wire  _T_3397 = _T_3311[5:0] == 6'h26; // @[el2_lib.scala 317:41]
  wire  _T_3395 = _T_3311[5:0] == 6'h25; // @[el2_lib.scala 317:41]
  wire  _T_3393 = _T_3311[5:0] == 6'h24; // @[el2_lib.scala 317:41]
  wire  _T_3391 = _T_3311[5:0] == 6'h23; // @[el2_lib.scala 317:41]
  wire  _T_3389 = _T_3311[5:0] == 6'h22; // @[el2_lib.scala 317:41]
  wire  _T_3387 = _T_3311[5:0] == 6'h21; // @[el2_lib.scala 317:41]
  wire  _T_3385 = _T_3311[5:0] == 6'h20; // @[el2_lib.scala 317:41]
  wire  _T_3383 = _T_3311[5:0] == 6'h1f; // @[el2_lib.scala 317:41]
  wire  _T_3381 = _T_3311[5:0] == 6'h1e; // @[el2_lib.scala 317:41]
  wire [9:0] _T_3457 = {_T_3399,_T_3397,_T_3395,_T_3393,_T_3391,_T_3389,_T_3387,_T_3385,_T_3383,_T_3381}; // @[el2_lib.scala 320:69]
  wire  _T_3379 = _T_3311[5:0] == 6'h1d; // @[el2_lib.scala 317:41]
  wire  _T_3377 = _T_3311[5:0] == 6'h1c; // @[el2_lib.scala 317:41]
  wire  _T_3375 = _T_3311[5:0] == 6'h1b; // @[el2_lib.scala 317:41]
  wire  _T_3373 = _T_3311[5:0] == 6'h1a; // @[el2_lib.scala 317:41]
  wire  _T_3371 = _T_3311[5:0] == 6'h19; // @[el2_lib.scala 317:41]
  wire  _T_3369 = _T_3311[5:0] == 6'h18; // @[el2_lib.scala 317:41]
  wire  _T_3367 = _T_3311[5:0] == 6'h17; // @[el2_lib.scala 317:41]
  wire  _T_3365 = _T_3311[5:0] == 6'h16; // @[el2_lib.scala 317:41]
  wire  _T_3363 = _T_3311[5:0] == 6'h15; // @[el2_lib.scala 317:41]
  wire  _T_3361 = _T_3311[5:0] == 6'h14; // @[el2_lib.scala 317:41]
  wire [9:0] _T_3448 = {_T_3379,_T_3377,_T_3375,_T_3373,_T_3371,_T_3369,_T_3367,_T_3365,_T_3363,_T_3361}; // @[el2_lib.scala 320:69]
  wire  _T_3359 = _T_3311[5:0] == 6'h13; // @[el2_lib.scala 317:41]
  wire  _T_3357 = _T_3311[5:0] == 6'h12; // @[el2_lib.scala 317:41]
  wire  _T_3355 = _T_3311[5:0] == 6'h11; // @[el2_lib.scala 317:41]
  wire  _T_3353 = _T_3311[5:0] == 6'h10; // @[el2_lib.scala 317:41]
  wire  _T_3351 = _T_3311[5:0] == 6'hf; // @[el2_lib.scala 317:41]
  wire  _T_3349 = _T_3311[5:0] == 6'he; // @[el2_lib.scala 317:41]
  wire  _T_3347 = _T_3311[5:0] == 6'hd; // @[el2_lib.scala 317:41]
  wire  _T_3345 = _T_3311[5:0] == 6'hc; // @[el2_lib.scala 317:41]
  wire  _T_3343 = _T_3311[5:0] == 6'hb; // @[el2_lib.scala 317:41]
  wire  _T_3341 = _T_3311[5:0] == 6'ha; // @[el2_lib.scala 317:41]
  wire [9:0] _T_3438 = {_T_3359,_T_3357,_T_3355,_T_3353,_T_3351,_T_3349,_T_3347,_T_3345,_T_3343,_T_3341}; // @[el2_lib.scala 320:69]
  wire  _T_3339 = _T_3311[5:0] == 6'h9; // @[el2_lib.scala 317:41]
  wire  _T_3337 = _T_3311[5:0] == 6'h8; // @[el2_lib.scala 317:41]
  wire  _T_3335 = _T_3311[5:0] == 6'h7; // @[el2_lib.scala 317:41]
  wire  _T_3333 = _T_3311[5:0] == 6'h6; // @[el2_lib.scala 317:41]
  wire  _T_3331 = _T_3311[5:0] == 6'h5; // @[el2_lib.scala 317:41]
  wire  _T_3329 = _T_3311[5:0] == 6'h4; // @[el2_lib.scala 317:41]
  wire  _T_3327 = _T_3311[5:0] == 6'h3; // @[el2_lib.scala 317:41]
  wire  _T_3325 = _T_3311[5:0] == 6'h2; // @[el2_lib.scala 317:41]
  wire  _T_3323 = _T_3311[5:0] == 6'h1; // @[el2_lib.scala 317:41]
  wire [18:0] _T_3439 = {_T_3438,_T_3339,_T_3337,_T_3335,_T_3333,_T_3331,_T_3329,_T_3327,_T_3325,_T_3323}; // @[el2_lib.scala 320:69]
  wire [38:0] _T_3459 = {_T_3457,_T_3448,_T_3439}; // @[el2_lib.scala 320:69]
  wire [7:0] _T_3414 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3420 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3414}; // @[Cat.scala 29:58]
  wire [38:0] _T_3460 = _T_3459 ^ _T_3420; // @[el2_lib.scala 320:76]
  wire [38:0] _T_3461 = _T_3315 ? _T_3460 : _T_3420; // @[el2_lib.scala 320:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3461[37:32],_T_3461[30:16],_T_3461[14:8],_T_3461[6:4],_T_3461[2]}; // @[Cat.scala 29:58]
  wire  _T_3784 = _T_3696[5:0] == 6'h27; // @[el2_lib.scala 317:41]
  wire  _T_3782 = _T_3696[5:0] == 6'h26; // @[el2_lib.scala 317:41]
  wire  _T_3780 = _T_3696[5:0] == 6'h25; // @[el2_lib.scala 317:41]
  wire  _T_3778 = _T_3696[5:0] == 6'h24; // @[el2_lib.scala 317:41]
  wire  _T_3776 = _T_3696[5:0] == 6'h23; // @[el2_lib.scala 317:41]
  wire  _T_3774 = _T_3696[5:0] == 6'h22; // @[el2_lib.scala 317:41]
  wire  _T_3772 = _T_3696[5:0] == 6'h21; // @[el2_lib.scala 317:41]
  wire  _T_3770 = _T_3696[5:0] == 6'h20; // @[el2_lib.scala 317:41]
  wire  _T_3768 = _T_3696[5:0] == 6'h1f; // @[el2_lib.scala 317:41]
  wire  _T_3766 = _T_3696[5:0] == 6'h1e; // @[el2_lib.scala 317:41]
  wire [9:0] _T_3842 = {_T_3784,_T_3782,_T_3780,_T_3778,_T_3776,_T_3774,_T_3772,_T_3770,_T_3768,_T_3766}; // @[el2_lib.scala 320:69]
  wire  _T_3764 = _T_3696[5:0] == 6'h1d; // @[el2_lib.scala 317:41]
  wire  _T_3762 = _T_3696[5:0] == 6'h1c; // @[el2_lib.scala 317:41]
  wire  _T_3760 = _T_3696[5:0] == 6'h1b; // @[el2_lib.scala 317:41]
  wire  _T_3758 = _T_3696[5:0] == 6'h1a; // @[el2_lib.scala 317:41]
  wire  _T_3756 = _T_3696[5:0] == 6'h19; // @[el2_lib.scala 317:41]
  wire  _T_3754 = _T_3696[5:0] == 6'h18; // @[el2_lib.scala 317:41]
  wire  _T_3752 = _T_3696[5:0] == 6'h17; // @[el2_lib.scala 317:41]
  wire  _T_3750 = _T_3696[5:0] == 6'h16; // @[el2_lib.scala 317:41]
  wire  _T_3748 = _T_3696[5:0] == 6'h15; // @[el2_lib.scala 317:41]
  wire  _T_3746 = _T_3696[5:0] == 6'h14; // @[el2_lib.scala 317:41]
  wire [9:0] _T_3833 = {_T_3764,_T_3762,_T_3760,_T_3758,_T_3756,_T_3754,_T_3752,_T_3750,_T_3748,_T_3746}; // @[el2_lib.scala 320:69]
  wire  _T_3744 = _T_3696[5:0] == 6'h13; // @[el2_lib.scala 317:41]
  wire  _T_3742 = _T_3696[5:0] == 6'h12; // @[el2_lib.scala 317:41]
  wire  _T_3740 = _T_3696[5:0] == 6'h11; // @[el2_lib.scala 317:41]
  wire  _T_3738 = _T_3696[5:0] == 6'h10; // @[el2_lib.scala 317:41]
  wire  _T_3736 = _T_3696[5:0] == 6'hf; // @[el2_lib.scala 317:41]
  wire  _T_3734 = _T_3696[5:0] == 6'he; // @[el2_lib.scala 317:41]
  wire  _T_3732 = _T_3696[5:0] == 6'hd; // @[el2_lib.scala 317:41]
  wire  _T_3730 = _T_3696[5:0] == 6'hc; // @[el2_lib.scala 317:41]
  wire  _T_3728 = _T_3696[5:0] == 6'hb; // @[el2_lib.scala 317:41]
  wire  _T_3726 = _T_3696[5:0] == 6'ha; // @[el2_lib.scala 317:41]
  wire [9:0] _T_3823 = {_T_3744,_T_3742,_T_3740,_T_3738,_T_3736,_T_3734,_T_3732,_T_3730,_T_3728,_T_3726}; // @[el2_lib.scala 320:69]
  wire  _T_3724 = _T_3696[5:0] == 6'h9; // @[el2_lib.scala 317:41]
  wire  _T_3722 = _T_3696[5:0] == 6'h8; // @[el2_lib.scala 317:41]
  wire  _T_3720 = _T_3696[5:0] == 6'h7; // @[el2_lib.scala 317:41]
  wire  _T_3718 = _T_3696[5:0] == 6'h6; // @[el2_lib.scala 317:41]
  wire  _T_3716 = _T_3696[5:0] == 6'h5; // @[el2_lib.scala 317:41]
  wire  _T_3714 = _T_3696[5:0] == 6'h4; // @[el2_lib.scala 317:41]
  wire  _T_3712 = _T_3696[5:0] == 6'h3; // @[el2_lib.scala 317:41]
  wire  _T_3710 = _T_3696[5:0] == 6'h2; // @[el2_lib.scala 317:41]
  wire  _T_3708 = _T_3696[5:0] == 6'h1; // @[el2_lib.scala 317:41]
  wire [18:0] _T_3824 = {_T_3823,_T_3724,_T_3722,_T_3720,_T_3718,_T_3716,_T_3714,_T_3712,_T_3710,_T_3708}; // @[el2_lib.scala 320:69]
  wire [38:0] _T_3844 = {_T_3842,_T_3833,_T_3824}; // @[el2_lib.scala 320:69]
  wire [7:0] _T_3799 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3805 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3799}; // @[Cat.scala 29:58]
  wire [38:0] _T_3845 = _T_3844 ^ _T_3805; // @[el2_lib.scala 320:76]
  wire [38:0] _T_3846 = _T_3700 ? _T_3845 : _T_3805; // @[el2_lib.scala 320:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3846[37:32],_T_3846[30:16],_T_3846[14:8],_T_3846[6:4],_T_3846[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 646:35]
  wire  _T_3319 = ~_T_3311[6]; // @[el2_lib.scala 313:55]
  wire  _T_3320 = _T_3313 & _T_3319; // @[el2_lib.scala 313:53]
  wire  _T_3704 = ~_T_3696[6]; // @[el2_lib.scala 313:55]
  wire  _T_3705 = _T_3698 & _T_3704; // @[el2_lib.scala 313:53]
  wire [1:0] iccm_double_ecc_error = {_T_3320,_T_3705}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 648:53]
  wire [63:0] _T_3070 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3071 = {iccm_dma_rdata_1_muxed,_T_3461[37:32],_T_3461[30:16],_T_3461[14:8],_T_3461[6:4],_T_3461[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 650:54]
  reg [2:0] iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 651:74]
  reg  iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 656:76]
  reg [63:0] iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 660:75]
  wire  _T_3076 = _T_2675 & _T_2664; // @[el2_ifu_mem_ctl.scala 663:65]
  wire  _T_3080 = _T_3057 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 664:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3081 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [14:0] _T_3083 = _T_3080 ? _T_3081 : io_ifc_fetch_addr_bf[14:0]; // @[el2_ifu_mem_ctl.scala 664:8]
  wire  _T_3473 = _T_3311 == 7'h40; // @[el2_lib.scala 323:62]
  wire  _T_3474 = _T_3461[38] ^ _T_3473; // @[el2_lib.scala 323:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3474,_T_3461[31],_T_3461[15],_T_3461[7],_T_3461[3],_T_3461[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3858 = _T_3696 == 7'h40; // @[el2_lib.scala 323:62]
  wire  _T_3859 = _T_3846[38] ^ _T_3858; // @[el2_lib.scala 323:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3859,_T_3846[31],_T_3846[15],_T_3846[7],_T_3846[3],_T_3846[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3875 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 676:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 678:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 679:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 687:62]
  wire  _T_3883 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 681:76]
  wire  _T_3884 = io_iccm_rd_ecc_single_err & _T_3883; // @[el2_ifu_mem_ctl.scala 681:74]
  wire  _T_3886 = _T_3884 & _T_319; // @[el2_ifu_mem_ctl.scala 681:104]
  wire  iccm_ecc_write_status = _T_3886 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 681:127]
  wire  _T_3887 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 682:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3887 & _T_319; // @[el2_ifu_mem_ctl.scala 682:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 686:51]
  wire [13:0] _T_3892 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 685:102]
  wire [38:0] _T_3896 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3901 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 690:41]
  wire  _T_3902 = io_ifc_fetch_req_bf & _T_3901; // @[el2_ifu_mem_ctl.scala 690:39]
  wire  _T_3903 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 690:72]
  wire  _T_3904 = _T_3902 & _T_3903; // @[el2_ifu_mem_ctl.scala 690:70]
  wire  _T_3906 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 691:34]
  wire  _T_3907 = _T_2235 & _T_3906; // @[el2_ifu_mem_ctl.scala 691:32]
  wire  _T_3910 = _T_2251 & _T_3906; // @[el2_ifu_mem_ctl.scala 692:37]
  wire  _T_3911 = _T_3907 | _T_3910; // @[el2_ifu_mem_ctl.scala 691:88]
  wire  _T_3912 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 693:19]
  wire  _T_3914 = _T_3912 & _T_3906; // @[el2_ifu_mem_ctl.scala 693:41]
  wire  _T_3915 = _T_3911 | _T_3914; // @[el2_ifu_mem_ctl.scala 692:88]
  wire  _T_3916 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 694:19]
  wire  _T_3918 = _T_3916 & _T_3906; // @[el2_ifu_mem_ctl.scala 694:35]
  wire  _T_3919 = _T_3915 | _T_3918; // @[el2_ifu_mem_ctl.scala 693:88]
  wire  _T_3922 = _T_2250 & _T_3906; // @[el2_ifu_mem_ctl.scala 695:38]
  wire  _T_3923 = _T_3919 | _T_3922; // @[el2_ifu_mem_ctl.scala 694:88]
  wire  _T_3925 = _T_2251 & miss_state_en; // @[el2_ifu_mem_ctl.scala 696:37]
  wire  _T_3926 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 696:71]
  wire  _T_3927 = _T_3925 & _T_3926; // @[el2_ifu_mem_ctl.scala 696:54]
  wire  _T_3928 = _T_3923 | _T_3927; // @[el2_ifu_mem_ctl.scala 695:57]
  wire  _T_3929 = ~_T_3928; // @[el2_ifu_mem_ctl.scala 691:5]
  wire  _T_3930 = _T_3904 & _T_3929; // @[el2_ifu_mem_ctl.scala 690:96]
  wire  _T_3931 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 697:28]
  wire  _T_3933 = _T_3931 & _T_3901; // @[el2_ifu_mem_ctl.scala 697:50]
  wire  _T_3935 = _T_3933 & _T_3903; // @[el2_ifu_mem_ctl.scala 697:81]
  wire [1:0] _T_3938 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10376 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 792:74]
  wire  bus_wren_1 = _T_10376 & miss_pending; // @[el2_ifu_mem_ctl.scala 792:98]
  wire  _T_10375 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 792:74]
  wire  bus_wren_0 = _T_10375 & miss_pending; // @[el2_ifu_mem_ctl.scala 792:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_3944 = ~_T_108; // @[el2_ifu_mem_ctl.scala 700:106]
  wire  _T_3945 = _T_2235 & _T_3944; // @[el2_ifu_mem_ctl.scala 700:104]
  wire  _T_3946 = _T_2251 | _T_3945; // @[el2_ifu_mem_ctl.scala 700:77]
  wire  _T_3950 = ~_T_51; // @[el2_ifu_mem_ctl.scala 700:172]
  wire  _T_3951 = _T_3946 & _T_3950; // @[el2_ifu_mem_ctl.scala 700:170]
  wire  _T_3952 = ~_T_3951; // @[el2_ifu_mem_ctl.scala 700:44]
  wire  _T_3956 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 703:64]
  wire  _T_3957 = ~_T_3956; // @[el2_ifu_mem_ctl.scala 703:50]
  wire  _T_3958 = _T_276 & _T_3957; // @[el2_ifu_mem_ctl.scala 703:48]
  wire  _T_3959 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 703:81]
  wire  ic_valid = _T_3958 & _T_3959; // @[el2_ifu_mem_ctl.scala 703:79]
  wire  _T_3961 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 704:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 707:14]
  wire  _T_3964 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 710:74]
  wire  _T_10373 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 791:45]
  wire  way_status_wr_en = _T_10373 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 791:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3964; // @[el2_ifu_mem_ctl.scala 710:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 712:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 787:41]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 718:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 720:132]
  wire  _T_3984 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_3985 = _T_3984 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_3986 = _T_3985 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_3989 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_3990 = _T_3989 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_3991 = _T_3990 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_3994 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_3995 = _T_3994 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_3996 = _T_3995 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_3999 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_4000 = _T_3999 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_4001 = _T_4000 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4004 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_4005 = _T_4004 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_4006 = _T_4005 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4009 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_4010 = _T_4009 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_4011 = _T_4010 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4014 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_4015 = _T_4014 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_4016 = _T_4015 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4019 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 724:100]
  wire  _T_4020 = _T_4019 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:108]
  wire  _T_4021 = _T_4020 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4026 = _T_3985 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4031 = _T_3990 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4036 = _T_3995 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4041 = _T_4000 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4046 = _T_4005 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4051 = _T_4010 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4056 = _T_4015 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4061 = _T_4020 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4066 = _T_3985 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4071 = _T_3990 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4076 = _T_3995 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4081 = _T_4000 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4086 = _T_4005 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4091 = _T_4010 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4096 = _T_4015 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4101 = _T_4020 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4106 = _T_3985 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4111 = _T_3990 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4116 = _T_3995 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4121 = _T_4000 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4126 = _T_4005 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4131 = _T_4010 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4136 = _T_4015 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4141 = _T_4020 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4146 = _T_3985 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4151 = _T_3990 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4156 = _T_3995 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4161 = _T_4000 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4166 = _T_4005 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4171 = _T_4010 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4176 = _T_4015 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4181 = _T_4020 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4186 = _T_3985 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4191 = _T_3990 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4196 = _T_3995 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4201 = _T_4000 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4206 = _T_4005 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4211 = _T_4010 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4216 = _T_4015 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4221 = _T_4020 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4226 = _T_3985 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4231 = _T_3990 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4236 = _T_3995 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4241 = _T_4000 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4246 = _T_4005 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4251 = _T_4010 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4256 = _T_4015 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4261 = _T_4020 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4266 = _T_3985 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4271 = _T_3990 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4276 = _T_3995 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4281 = _T_4000 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4286 = _T_4005 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4291 = _T_4010 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4296 = _T_4015 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4301 = _T_4020 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4306 = _T_3985 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4311 = _T_3990 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4316 = _T_3995 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4321 = _T_4000 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4326 = _T_4005 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4331 = _T_4010 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4336 = _T_4015 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4341 = _T_4020 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4346 = _T_3985 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4351 = _T_3990 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4356 = _T_3995 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4361 = _T_4000 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4366 = _T_4005 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4371 = _T_4010 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4376 = _T_4015 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4381 = _T_4020 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4386 = _T_3985 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4391 = _T_3990 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4396 = _T_3995 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4401 = _T_4000 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4406 = _T_4005 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4411 = _T_4010 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4416 = _T_4015 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4421 = _T_4020 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4426 = _T_3985 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4431 = _T_3990 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4436 = _T_3995 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4441 = _T_4000 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4446 = _T_4005 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4451 = _T_4010 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4456 = _T_4015 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4461 = _T_4020 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4466 = _T_3985 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4471 = _T_3990 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4476 = _T_3995 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4481 = _T_4000 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4486 = _T_4005 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4491 = _T_4010 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4496 = _T_4015 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4501 = _T_4020 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4506 = _T_3985 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4511 = _T_3990 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4516 = _T_3995 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4521 = _T_4000 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4526 = _T_4005 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4531 = _T_4010 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4536 = _T_4015 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4541 = _T_4020 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4546 = _T_3985 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4551 = _T_3990 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4556 = _T_3995 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4561 = _T_4000 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4566 = _T_4005 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4571 = _T_4010 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4576 = _T_4015 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4581 = _T_4020 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4586 = _T_3985 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4591 = _T_3990 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4596 = _T_3995 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4601 = _T_4000 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4606 = _T_4005 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4611 = _T_4010 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4616 = _T_4015 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_4621 = _T_4020 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 724:131]
  wire  _T_10379 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 794:84]
  wire  _T_10380 = _T_10379 & miss_pending; // @[el2_ifu_mem_ctl.scala 794:108]
  wire  bus_wren_last_1 = _T_10380 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 794:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_10382 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 796:73]
  wire  _T_10377 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 794:84]
  wire  _T_10378 = _T_10377 & miss_pending; // @[el2_ifu_mem_ctl.scala 794:108]
  wire  bus_wren_last_0 = _T_10378 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 794:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_10381 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 796:73]
  wire [1:0] ifu_tag_wren = {_T_10382,_T_10381}; // @[Cat.scala 29:58]
  wire [1:0] _T_10417 = _T_3964 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10417 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 830:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 737:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 739:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 743:14]
  wire  _T_5155 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 747:78]
  wire  _T_5157 = _T_5155 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5159 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 748:70]
  wire  _T_5161 = _T_5159 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5162 = _T_5157 | _T_5161; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5163 = _T_5162 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire  _T_5167 = _T_5155 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5171 = _T_5159 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5172 = _T_5167 | _T_5171; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5173 = _T_5172 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire [1:0] tag_valid_clken_0 = {_T_5173,_T_5163}; // @[Cat.scala 29:58]
  wire  _T_5175 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 747:78]
  wire  _T_5177 = _T_5175 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5179 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 748:70]
  wire  _T_5181 = _T_5179 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5182 = _T_5177 | _T_5181; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5183 = _T_5182 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire  _T_5187 = _T_5175 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5191 = _T_5179 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5192 = _T_5187 | _T_5191; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5193 = _T_5192 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire [1:0] tag_valid_clken_1 = {_T_5193,_T_5183}; // @[Cat.scala 29:58]
  wire  _T_5195 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 747:78]
  wire  _T_5197 = _T_5195 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5199 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 748:70]
  wire  _T_5201 = _T_5199 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5202 = _T_5197 | _T_5201; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5203 = _T_5202 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire  _T_5207 = _T_5195 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5211 = _T_5199 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5212 = _T_5207 | _T_5211; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5213 = _T_5212 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire [1:0] tag_valid_clken_2 = {_T_5213,_T_5203}; // @[Cat.scala 29:58]
  wire  _T_5215 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 747:78]
  wire  _T_5217 = _T_5215 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5219 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 748:70]
  wire  _T_5221 = _T_5219 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5222 = _T_5217 | _T_5221; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5223 = _T_5222 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire  _T_5227 = _T_5215 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 747:87]
  wire  _T_5231 = _T_5219 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 748:79]
  wire  _T_5232 = _T_5227 | _T_5231; // @[el2_ifu_mem_ctl.scala 747:109]
  wire  _T_5233 = _T_5232 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 748:102]
  wire [1:0] tag_valid_clken_3 = {_T_5233,_T_5223}; // @[Cat.scala 29:58]
  wire  _T_5236 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 756:66]
  wire  _T_5237 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 756:93]
  wire  _T_5238 = _T_5236 & _T_5237; // @[el2_ifu_mem_ctl.scala 756:91]
  wire  _T_5241 = _T_4763 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5242 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5244 = _T_5242 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5245 = _T_5241 | _T_5244; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5246 = _T_5245 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5248 = _T_5246 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5258 = _T_4764 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5259 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5261 = _T_5259 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5262 = _T_5258 | _T_5261; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5263 = _T_5262 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5265 = _T_5263 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5275 = _T_4765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5276 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5278 = _T_5276 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5279 = _T_5275 | _T_5278; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5280 = _T_5279 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5282 = _T_5280 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5292 = _T_4766 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5293 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5295 = _T_5293 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5296 = _T_5292 | _T_5295; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5297 = _T_5296 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5299 = _T_5297 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5309 = _T_4767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5310 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5312 = _T_5310 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5313 = _T_5309 | _T_5312; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5314 = _T_5313 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5316 = _T_5314 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5326 = _T_4768 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5327 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5329 = _T_5327 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5330 = _T_5326 | _T_5329; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5331 = _T_5330 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5333 = _T_5331 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5343 = _T_4769 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5344 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5346 = _T_5344 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5347 = _T_5343 | _T_5346; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5348 = _T_5347 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5350 = _T_5348 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5360 = _T_4770 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5361 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5363 = _T_5361 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5364 = _T_5360 | _T_5363; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5365 = _T_5364 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5367 = _T_5365 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5377 = _T_4771 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5378 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5380 = _T_5378 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5381 = _T_5377 | _T_5380; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5382 = _T_5381 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5384 = _T_5382 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5394 = _T_4772 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5395 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5397 = _T_5395 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5398 = _T_5394 | _T_5397; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5399 = _T_5398 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5401 = _T_5399 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5411 = _T_4773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5412 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5414 = _T_5412 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5415 = _T_5411 | _T_5414; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5416 = _T_5415 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5418 = _T_5416 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5428 = _T_4774 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5429 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5431 = _T_5429 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5432 = _T_5428 | _T_5431; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5433 = _T_5432 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5435 = _T_5433 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5445 = _T_4775 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5446 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5448 = _T_5446 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5449 = _T_5445 | _T_5448; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5450 = _T_5449 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5452 = _T_5450 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5462 = _T_4776 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5463 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5465 = _T_5463 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5466 = _T_5462 | _T_5465; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5467 = _T_5466 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5469 = _T_5467 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5479 = _T_4777 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5480 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5482 = _T_5480 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5483 = _T_5479 | _T_5482; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5484 = _T_5483 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5486 = _T_5484 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5496 = _T_4778 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5497 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5499 = _T_5497 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5500 = _T_5496 | _T_5499; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5501 = _T_5500 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5503 = _T_5501 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5513 = _T_4779 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5514 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5516 = _T_5514 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5517 = _T_5513 | _T_5516; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5518 = _T_5517 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5520 = _T_5518 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5530 = _T_4780 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5531 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5533 = _T_5531 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5534 = _T_5530 | _T_5533; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5535 = _T_5534 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5537 = _T_5535 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5547 = _T_4781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5548 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5550 = _T_5548 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5551 = _T_5547 | _T_5550; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5552 = _T_5551 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5554 = _T_5552 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5564 = _T_4782 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5565 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5567 = _T_5565 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5568 = _T_5564 | _T_5567; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5569 = _T_5568 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5571 = _T_5569 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5581 = _T_4783 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5582 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5584 = _T_5582 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5585 = _T_5581 | _T_5584; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5586 = _T_5585 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5588 = _T_5586 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5598 = _T_4784 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5599 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5601 = _T_5599 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5602 = _T_5598 | _T_5601; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5603 = _T_5602 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5605 = _T_5603 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5615 = _T_4785 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5616 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5618 = _T_5616 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5619 = _T_5615 | _T_5618; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5620 = _T_5619 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5622 = _T_5620 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5632 = _T_4786 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5633 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5635 = _T_5633 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5636 = _T_5632 | _T_5635; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5637 = _T_5636 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5639 = _T_5637 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5649 = _T_4787 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5650 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5652 = _T_5650 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5653 = _T_5649 | _T_5652; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5654 = _T_5653 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5656 = _T_5654 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5666 = _T_4788 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5667 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5669 = _T_5667 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5670 = _T_5666 | _T_5669; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5671 = _T_5670 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5673 = _T_5671 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5683 = _T_4789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5684 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5686 = _T_5684 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5687 = _T_5683 | _T_5686; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5688 = _T_5687 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5690 = _T_5688 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5700 = _T_4790 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5701 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5703 = _T_5701 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5704 = _T_5700 | _T_5703; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5705 = _T_5704 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5707 = _T_5705 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5717 = _T_4791 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5718 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5720 = _T_5718 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5721 = _T_5717 | _T_5720; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5722 = _T_5721 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5724 = _T_5722 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5734 = _T_4792 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5735 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5737 = _T_5735 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5738 = _T_5734 | _T_5737; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5739 = _T_5738 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5741 = _T_5739 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5751 = _T_4793 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5752 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5754 = _T_5752 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5755 = _T_5751 | _T_5754; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5756 = _T_5755 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5758 = _T_5756 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5768 = _T_4794 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5769 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_5771 = _T_5769 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5772 = _T_5768 | _T_5771; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5773 = _T_5772 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5775 = _T_5773 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5785 = _T_4763 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5788 = _T_5242 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5789 = _T_5785 | _T_5788; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5790 = _T_5789 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5792 = _T_5790 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5802 = _T_4764 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5805 = _T_5259 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5806 = _T_5802 | _T_5805; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5807 = _T_5806 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5809 = _T_5807 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5819 = _T_4765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5822 = _T_5276 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5823 = _T_5819 | _T_5822; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5824 = _T_5823 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5826 = _T_5824 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5836 = _T_4766 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5839 = _T_5293 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5840 = _T_5836 | _T_5839; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5841 = _T_5840 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5843 = _T_5841 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5853 = _T_4767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5856 = _T_5310 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5857 = _T_5853 | _T_5856; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5858 = _T_5857 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5860 = _T_5858 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5870 = _T_4768 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5873 = _T_5327 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5874 = _T_5870 | _T_5873; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5875 = _T_5874 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5877 = _T_5875 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5887 = _T_4769 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5890 = _T_5344 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5891 = _T_5887 | _T_5890; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5892 = _T_5891 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5894 = _T_5892 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5904 = _T_4770 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5907 = _T_5361 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5908 = _T_5904 | _T_5907; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5909 = _T_5908 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5911 = _T_5909 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5921 = _T_4771 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5924 = _T_5378 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5925 = _T_5921 | _T_5924; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5926 = _T_5925 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5928 = _T_5926 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5938 = _T_4772 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5941 = _T_5395 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5942 = _T_5938 | _T_5941; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5943 = _T_5942 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5945 = _T_5943 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5955 = _T_4773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5958 = _T_5412 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5959 = _T_5955 | _T_5958; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5960 = _T_5959 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5962 = _T_5960 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5972 = _T_4774 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5975 = _T_5429 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5976 = _T_5972 | _T_5975; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5977 = _T_5976 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5979 = _T_5977 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_5989 = _T_4775 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_5992 = _T_5446 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_5993 = _T_5989 | _T_5992; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_5994 = _T_5993 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_5996 = _T_5994 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6006 = _T_4776 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6009 = _T_5463 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6010 = _T_6006 | _T_6009; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6011 = _T_6010 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6013 = _T_6011 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6023 = _T_4777 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6026 = _T_5480 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6027 = _T_6023 | _T_6026; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6028 = _T_6027 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6030 = _T_6028 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6040 = _T_4778 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6043 = _T_5497 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6044 = _T_6040 | _T_6043; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6045 = _T_6044 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6047 = _T_6045 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6057 = _T_4779 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6060 = _T_5514 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6061 = _T_6057 | _T_6060; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6062 = _T_6061 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6064 = _T_6062 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6074 = _T_4780 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6077 = _T_5531 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6078 = _T_6074 | _T_6077; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6079 = _T_6078 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6081 = _T_6079 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6091 = _T_4781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6094 = _T_5548 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6095 = _T_6091 | _T_6094; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6096 = _T_6095 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6098 = _T_6096 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6108 = _T_4782 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6111 = _T_5565 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6112 = _T_6108 | _T_6111; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6113 = _T_6112 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6115 = _T_6113 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6125 = _T_4783 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6128 = _T_5582 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6129 = _T_6125 | _T_6128; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6130 = _T_6129 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6132 = _T_6130 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6142 = _T_4784 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6145 = _T_5599 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6146 = _T_6142 | _T_6145; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6147 = _T_6146 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6149 = _T_6147 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6159 = _T_4785 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6162 = _T_5616 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6163 = _T_6159 | _T_6162; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6164 = _T_6163 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6166 = _T_6164 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6176 = _T_4786 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6179 = _T_5633 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6180 = _T_6176 | _T_6179; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6181 = _T_6180 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6183 = _T_6181 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6193 = _T_4787 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6196 = _T_5650 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6197 = _T_6193 | _T_6196; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6198 = _T_6197 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6200 = _T_6198 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6210 = _T_4788 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6213 = _T_5667 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6214 = _T_6210 | _T_6213; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6215 = _T_6214 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6217 = _T_6215 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6227 = _T_4789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6230 = _T_5684 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6231 = _T_6227 | _T_6230; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6232 = _T_6231 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6234 = _T_6232 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6244 = _T_4790 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6247 = _T_5701 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6248 = _T_6244 | _T_6247; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6249 = _T_6248 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6251 = _T_6249 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6261 = _T_4791 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6264 = _T_5718 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6265 = _T_6261 | _T_6264; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6266 = _T_6265 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6268 = _T_6266 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6278 = _T_4792 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6281 = _T_5735 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6282 = _T_6278 | _T_6281; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6283 = _T_6282 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6285 = _T_6283 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6295 = _T_4793 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6298 = _T_5752 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6299 = _T_6295 | _T_6298; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6300 = _T_6299 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6302 = _T_6300 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6312 = _T_4794 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6315 = _T_5769 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6316 = _T_6312 | _T_6315; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6317 = _T_6316 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6319 = _T_6317 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6329 = _T_4795 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6330 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6332 = _T_6330 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6333 = _T_6329 | _T_6332; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6334 = _T_6333 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6336 = _T_6334 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6346 = _T_4796 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6347 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6349 = _T_6347 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6350 = _T_6346 | _T_6349; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6351 = _T_6350 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6353 = _T_6351 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6363 = _T_4797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6364 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6366 = _T_6364 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6367 = _T_6363 | _T_6366; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6368 = _T_6367 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6370 = _T_6368 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6380 = _T_4798 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6381 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6383 = _T_6381 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6384 = _T_6380 | _T_6383; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6385 = _T_6384 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6387 = _T_6385 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6397 = _T_4799 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6398 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6400 = _T_6398 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6401 = _T_6397 | _T_6400; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6402 = _T_6401 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6404 = _T_6402 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6414 = _T_4800 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6415 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6417 = _T_6415 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6418 = _T_6414 | _T_6417; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6419 = _T_6418 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6421 = _T_6419 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6431 = _T_4801 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6432 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6434 = _T_6432 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6435 = _T_6431 | _T_6434; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6436 = _T_6435 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6438 = _T_6436 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6448 = _T_4802 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6449 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6451 = _T_6449 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6452 = _T_6448 | _T_6451; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6453 = _T_6452 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6455 = _T_6453 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6465 = _T_4803 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6466 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6468 = _T_6466 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6469 = _T_6465 | _T_6468; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6470 = _T_6469 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6472 = _T_6470 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6482 = _T_4804 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6483 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6485 = _T_6483 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6486 = _T_6482 | _T_6485; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6487 = _T_6486 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6489 = _T_6487 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6499 = _T_4805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6500 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6502 = _T_6500 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6503 = _T_6499 | _T_6502; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6504 = _T_6503 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6506 = _T_6504 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6516 = _T_4806 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6517 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6519 = _T_6517 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6520 = _T_6516 | _T_6519; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6521 = _T_6520 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6523 = _T_6521 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6533 = _T_4807 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6534 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6536 = _T_6534 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6537 = _T_6533 | _T_6536; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6538 = _T_6537 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6540 = _T_6538 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6550 = _T_4808 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6551 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6553 = _T_6551 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6554 = _T_6550 | _T_6553; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6555 = _T_6554 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6557 = _T_6555 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6567 = _T_4809 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6568 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6570 = _T_6568 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6571 = _T_6567 | _T_6570; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6572 = _T_6571 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6574 = _T_6572 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6584 = _T_4810 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6585 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6587 = _T_6585 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6588 = _T_6584 | _T_6587; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6589 = _T_6588 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6591 = _T_6589 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6601 = _T_4811 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6602 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6604 = _T_6602 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6605 = _T_6601 | _T_6604; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6606 = _T_6605 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6608 = _T_6606 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6618 = _T_4812 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6619 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6621 = _T_6619 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6622 = _T_6618 | _T_6621; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6623 = _T_6622 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6625 = _T_6623 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6635 = _T_4813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6636 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6638 = _T_6636 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6639 = _T_6635 | _T_6638; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6640 = _T_6639 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6642 = _T_6640 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6652 = _T_4814 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6653 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6655 = _T_6653 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6656 = _T_6652 | _T_6655; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6657 = _T_6656 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6659 = _T_6657 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6669 = _T_4815 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6670 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6672 = _T_6670 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6673 = _T_6669 | _T_6672; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6674 = _T_6673 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6676 = _T_6674 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6686 = _T_4816 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6687 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6689 = _T_6687 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6690 = _T_6686 | _T_6689; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6691 = _T_6690 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6693 = _T_6691 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6703 = _T_4817 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6704 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6706 = _T_6704 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6707 = _T_6703 | _T_6706; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6708 = _T_6707 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6710 = _T_6708 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6720 = _T_4818 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6721 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6723 = _T_6721 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6724 = _T_6720 | _T_6723; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6725 = _T_6724 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6727 = _T_6725 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6737 = _T_4819 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6738 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6740 = _T_6738 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6741 = _T_6737 | _T_6740; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6742 = _T_6741 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6744 = _T_6742 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6754 = _T_4820 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6755 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6757 = _T_6755 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6758 = _T_6754 | _T_6757; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6759 = _T_6758 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6761 = _T_6759 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6771 = _T_4821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6772 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6774 = _T_6772 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6775 = _T_6771 | _T_6774; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6776 = _T_6775 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6778 = _T_6776 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6788 = _T_4822 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6789 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6791 = _T_6789 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6792 = _T_6788 | _T_6791; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6793 = _T_6792 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6795 = _T_6793 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6805 = _T_4823 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6806 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6808 = _T_6806 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6809 = _T_6805 | _T_6808; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6810 = _T_6809 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6812 = _T_6810 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6822 = _T_4824 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6823 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6825 = _T_6823 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6826 = _T_6822 | _T_6825; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6827 = _T_6826 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6829 = _T_6827 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6839 = _T_4825 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6840 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6842 = _T_6840 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6843 = _T_6839 | _T_6842; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6844 = _T_6843 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6846 = _T_6844 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6856 = _T_4826 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6857 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_6859 = _T_6857 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6860 = _T_6856 | _T_6859; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6861 = _T_6860 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6863 = _T_6861 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6873 = _T_4795 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6876 = _T_6330 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6877 = _T_6873 | _T_6876; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6878 = _T_6877 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6880 = _T_6878 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6890 = _T_4796 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6893 = _T_6347 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6894 = _T_6890 | _T_6893; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6895 = _T_6894 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6897 = _T_6895 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6907 = _T_4797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6910 = _T_6364 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6911 = _T_6907 | _T_6910; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6912 = _T_6911 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6914 = _T_6912 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6924 = _T_4798 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6927 = _T_6381 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6928 = _T_6924 | _T_6927; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6929 = _T_6928 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6931 = _T_6929 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6941 = _T_4799 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6944 = _T_6398 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6945 = _T_6941 | _T_6944; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6946 = _T_6945 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6948 = _T_6946 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6958 = _T_4800 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6961 = _T_6415 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6962 = _T_6958 | _T_6961; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6963 = _T_6962 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6965 = _T_6963 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6975 = _T_4801 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6978 = _T_6432 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6979 = _T_6975 | _T_6978; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6980 = _T_6979 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6982 = _T_6980 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_6992 = _T_4802 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_6995 = _T_6449 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_6996 = _T_6992 | _T_6995; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_6997 = _T_6996 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_6999 = _T_6997 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7009 = _T_4803 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7012 = _T_6466 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7013 = _T_7009 | _T_7012; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7014 = _T_7013 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7016 = _T_7014 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7026 = _T_4804 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7029 = _T_6483 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7030 = _T_7026 | _T_7029; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7031 = _T_7030 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7033 = _T_7031 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7043 = _T_4805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7046 = _T_6500 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7047 = _T_7043 | _T_7046; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7048 = _T_7047 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7050 = _T_7048 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7060 = _T_4806 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7063 = _T_6517 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7064 = _T_7060 | _T_7063; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7065 = _T_7064 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7067 = _T_7065 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7077 = _T_4807 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7080 = _T_6534 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7081 = _T_7077 | _T_7080; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7082 = _T_7081 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7084 = _T_7082 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7094 = _T_4808 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7097 = _T_6551 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7098 = _T_7094 | _T_7097; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7099 = _T_7098 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7101 = _T_7099 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7111 = _T_4809 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7114 = _T_6568 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7115 = _T_7111 | _T_7114; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7116 = _T_7115 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7118 = _T_7116 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7128 = _T_4810 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7131 = _T_6585 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7132 = _T_7128 | _T_7131; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7133 = _T_7132 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7135 = _T_7133 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7145 = _T_4811 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7148 = _T_6602 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7149 = _T_7145 | _T_7148; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7150 = _T_7149 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7152 = _T_7150 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7162 = _T_4812 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7165 = _T_6619 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7166 = _T_7162 | _T_7165; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7167 = _T_7166 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7169 = _T_7167 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7179 = _T_4813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7182 = _T_6636 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7183 = _T_7179 | _T_7182; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7184 = _T_7183 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7186 = _T_7184 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7196 = _T_4814 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7199 = _T_6653 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7200 = _T_7196 | _T_7199; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7201 = _T_7200 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7203 = _T_7201 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7213 = _T_4815 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7216 = _T_6670 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7217 = _T_7213 | _T_7216; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7218 = _T_7217 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7220 = _T_7218 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7230 = _T_4816 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7233 = _T_6687 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7234 = _T_7230 | _T_7233; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7235 = _T_7234 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7237 = _T_7235 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7247 = _T_4817 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7250 = _T_6704 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7251 = _T_7247 | _T_7250; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7252 = _T_7251 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7254 = _T_7252 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7264 = _T_4818 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7267 = _T_6721 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7268 = _T_7264 | _T_7267; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7269 = _T_7268 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7271 = _T_7269 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7281 = _T_4819 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7284 = _T_6738 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7285 = _T_7281 | _T_7284; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7286 = _T_7285 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7288 = _T_7286 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7298 = _T_4820 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7301 = _T_6755 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7302 = _T_7298 | _T_7301; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7303 = _T_7302 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7305 = _T_7303 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7315 = _T_4821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7318 = _T_6772 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7319 = _T_7315 | _T_7318; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7320 = _T_7319 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7322 = _T_7320 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7332 = _T_4822 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7335 = _T_6789 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7336 = _T_7332 | _T_7335; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7337 = _T_7336 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7339 = _T_7337 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7349 = _T_4823 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7352 = _T_6806 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7353 = _T_7349 | _T_7352; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7354 = _T_7353 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7356 = _T_7354 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7366 = _T_4824 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7369 = _T_6823 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7370 = _T_7366 | _T_7369; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7371 = _T_7370 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7373 = _T_7371 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7383 = _T_4825 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7386 = _T_6840 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7387 = _T_7383 | _T_7386; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7388 = _T_7387 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7390 = _T_7388 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7400 = _T_4826 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7403 = _T_6857 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7404 = _T_7400 | _T_7403; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7405 = _T_7404 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7407 = _T_7405 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7417 = _T_4827 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7418 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7420 = _T_7418 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7421 = _T_7417 | _T_7420; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7422 = _T_7421 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7424 = _T_7422 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7434 = _T_4828 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7435 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7437 = _T_7435 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7438 = _T_7434 | _T_7437; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7439 = _T_7438 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7441 = _T_7439 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7451 = _T_4829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7452 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7454 = _T_7452 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7455 = _T_7451 | _T_7454; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7456 = _T_7455 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7458 = _T_7456 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7468 = _T_4830 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7469 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7471 = _T_7469 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7472 = _T_7468 | _T_7471; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7473 = _T_7472 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7475 = _T_7473 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7485 = _T_4831 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7486 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7488 = _T_7486 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7489 = _T_7485 | _T_7488; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7490 = _T_7489 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7492 = _T_7490 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7502 = _T_4832 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7503 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7505 = _T_7503 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7506 = _T_7502 | _T_7505; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7507 = _T_7506 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7509 = _T_7507 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7519 = _T_4833 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7520 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7522 = _T_7520 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7523 = _T_7519 | _T_7522; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7524 = _T_7523 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7526 = _T_7524 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7536 = _T_4834 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7537 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7539 = _T_7537 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7540 = _T_7536 | _T_7539; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7541 = _T_7540 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7543 = _T_7541 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7553 = _T_4835 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7554 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7556 = _T_7554 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7557 = _T_7553 | _T_7556; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7558 = _T_7557 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7560 = _T_7558 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7570 = _T_4836 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7571 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7573 = _T_7571 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7574 = _T_7570 | _T_7573; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7575 = _T_7574 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7577 = _T_7575 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7587 = _T_4837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7588 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7590 = _T_7588 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7591 = _T_7587 | _T_7590; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7592 = _T_7591 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7594 = _T_7592 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7604 = _T_4838 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7605 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7607 = _T_7605 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7608 = _T_7604 | _T_7607; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7609 = _T_7608 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7611 = _T_7609 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7621 = _T_4839 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7622 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7624 = _T_7622 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7625 = _T_7621 | _T_7624; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7626 = _T_7625 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7628 = _T_7626 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7638 = _T_4840 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7639 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7641 = _T_7639 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7642 = _T_7638 | _T_7641; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7643 = _T_7642 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7645 = _T_7643 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7655 = _T_4841 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7656 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7658 = _T_7656 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7659 = _T_7655 | _T_7658; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7660 = _T_7659 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7662 = _T_7660 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7672 = _T_4842 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7673 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7675 = _T_7673 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7676 = _T_7672 | _T_7675; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7677 = _T_7676 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7679 = _T_7677 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7689 = _T_4843 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7690 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7692 = _T_7690 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7693 = _T_7689 | _T_7692; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7694 = _T_7693 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7696 = _T_7694 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7706 = _T_4844 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7707 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7709 = _T_7707 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7710 = _T_7706 | _T_7709; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7711 = _T_7710 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7713 = _T_7711 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7723 = _T_4845 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7724 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7726 = _T_7724 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7727 = _T_7723 | _T_7726; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7728 = _T_7727 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7730 = _T_7728 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7740 = _T_4846 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7741 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7743 = _T_7741 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7744 = _T_7740 | _T_7743; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7745 = _T_7744 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7747 = _T_7745 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7757 = _T_4847 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7758 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7760 = _T_7758 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7761 = _T_7757 | _T_7760; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7762 = _T_7761 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7764 = _T_7762 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7774 = _T_4848 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7775 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7777 = _T_7775 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7778 = _T_7774 | _T_7777; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7779 = _T_7778 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7781 = _T_7779 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7791 = _T_4849 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7792 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7794 = _T_7792 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7795 = _T_7791 | _T_7794; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7796 = _T_7795 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7798 = _T_7796 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7808 = _T_4850 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7809 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7811 = _T_7809 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7812 = _T_7808 | _T_7811; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7813 = _T_7812 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7815 = _T_7813 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7825 = _T_4851 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7826 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7828 = _T_7826 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7829 = _T_7825 | _T_7828; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7830 = _T_7829 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7832 = _T_7830 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7842 = _T_4852 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7843 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7845 = _T_7843 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7846 = _T_7842 | _T_7845; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7847 = _T_7846 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7849 = _T_7847 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7859 = _T_4853 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7860 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7862 = _T_7860 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7863 = _T_7859 | _T_7862; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7864 = _T_7863 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7866 = _T_7864 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7876 = _T_4854 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7877 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7879 = _T_7877 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7880 = _T_7876 | _T_7879; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7881 = _T_7880 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7883 = _T_7881 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7893 = _T_4855 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7894 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7896 = _T_7894 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7897 = _T_7893 | _T_7896; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7898 = _T_7897 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7900 = _T_7898 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7910 = _T_4856 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7911 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7913 = _T_7911 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7914 = _T_7910 | _T_7913; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7915 = _T_7914 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7917 = _T_7915 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7927 = _T_4857 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7928 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7930 = _T_7928 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7931 = _T_7927 | _T_7930; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7932 = _T_7931 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7934 = _T_7932 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7944 = _T_4858 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7945 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_7947 = _T_7945 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7948 = _T_7944 | _T_7947; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7949 = _T_7948 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7951 = _T_7949 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7961 = _T_4827 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7964 = _T_7418 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7965 = _T_7961 | _T_7964; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7966 = _T_7965 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7968 = _T_7966 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7978 = _T_4828 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7981 = _T_7435 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7982 = _T_7978 | _T_7981; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_7983 = _T_7982 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_7985 = _T_7983 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_7995 = _T_4829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_7998 = _T_7452 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_7999 = _T_7995 | _T_7998; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8000 = _T_7999 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8002 = _T_8000 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8012 = _T_4830 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8015 = _T_7469 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8016 = _T_8012 | _T_8015; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8017 = _T_8016 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8019 = _T_8017 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8029 = _T_4831 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8032 = _T_7486 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8033 = _T_8029 | _T_8032; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8034 = _T_8033 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8036 = _T_8034 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8046 = _T_4832 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8049 = _T_7503 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8050 = _T_8046 | _T_8049; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8051 = _T_8050 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8053 = _T_8051 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8063 = _T_4833 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8066 = _T_7520 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8067 = _T_8063 | _T_8066; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8068 = _T_8067 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8070 = _T_8068 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8080 = _T_4834 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8083 = _T_7537 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8084 = _T_8080 | _T_8083; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8085 = _T_8084 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8087 = _T_8085 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8097 = _T_4835 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8100 = _T_7554 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8101 = _T_8097 | _T_8100; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8102 = _T_8101 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8104 = _T_8102 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8114 = _T_4836 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8117 = _T_7571 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8118 = _T_8114 | _T_8117; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8119 = _T_8118 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8121 = _T_8119 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8131 = _T_4837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8134 = _T_7588 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8135 = _T_8131 | _T_8134; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8136 = _T_8135 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8138 = _T_8136 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8148 = _T_4838 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8151 = _T_7605 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8152 = _T_8148 | _T_8151; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8153 = _T_8152 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8155 = _T_8153 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8165 = _T_4839 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8168 = _T_7622 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8169 = _T_8165 | _T_8168; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8170 = _T_8169 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8172 = _T_8170 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8182 = _T_4840 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8185 = _T_7639 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8186 = _T_8182 | _T_8185; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8187 = _T_8186 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8189 = _T_8187 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8199 = _T_4841 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8202 = _T_7656 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8203 = _T_8199 | _T_8202; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8204 = _T_8203 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8206 = _T_8204 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8216 = _T_4842 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8219 = _T_7673 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8220 = _T_8216 | _T_8219; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8221 = _T_8220 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8223 = _T_8221 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8233 = _T_4843 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8236 = _T_7690 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8237 = _T_8233 | _T_8236; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8238 = _T_8237 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8240 = _T_8238 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8250 = _T_4844 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8253 = _T_7707 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8254 = _T_8250 | _T_8253; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8255 = _T_8254 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8257 = _T_8255 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8267 = _T_4845 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8270 = _T_7724 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8271 = _T_8267 | _T_8270; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8272 = _T_8271 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8274 = _T_8272 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8284 = _T_4846 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8287 = _T_7741 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8288 = _T_8284 | _T_8287; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8289 = _T_8288 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8291 = _T_8289 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8301 = _T_4847 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8304 = _T_7758 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8305 = _T_8301 | _T_8304; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8306 = _T_8305 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8308 = _T_8306 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8318 = _T_4848 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8321 = _T_7775 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8322 = _T_8318 | _T_8321; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8323 = _T_8322 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8325 = _T_8323 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8335 = _T_4849 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8338 = _T_7792 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8339 = _T_8335 | _T_8338; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8340 = _T_8339 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8342 = _T_8340 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8352 = _T_4850 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8355 = _T_7809 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8356 = _T_8352 | _T_8355; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8357 = _T_8356 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8359 = _T_8357 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8369 = _T_4851 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8372 = _T_7826 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8373 = _T_8369 | _T_8372; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8374 = _T_8373 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8376 = _T_8374 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8386 = _T_4852 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8389 = _T_7843 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8390 = _T_8386 | _T_8389; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8391 = _T_8390 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8393 = _T_8391 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8403 = _T_4853 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8406 = _T_7860 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8407 = _T_8403 | _T_8406; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8408 = _T_8407 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8410 = _T_8408 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8420 = _T_4854 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8423 = _T_7877 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8424 = _T_8420 | _T_8423; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8425 = _T_8424 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8427 = _T_8425 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8437 = _T_4855 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8440 = _T_7894 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8441 = _T_8437 | _T_8440; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8442 = _T_8441 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8444 = _T_8442 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8454 = _T_4856 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8457 = _T_7911 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8458 = _T_8454 | _T_8457; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8459 = _T_8458 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8461 = _T_8459 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8471 = _T_4857 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8474 = _T_7928 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8475 = _T_8471 | _T_8474; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8476 = _T_8475 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8478 = _T_8476 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8488 = _T_4858 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8491 = _T_7945 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8492 = _T_8488 | _T_8491; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8493 = _T_8492 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8495 = _T_8493 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8505 = _T_4859 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8506 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8508 = _T_8506 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8509 = _T_8505 | _T_8508; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8510 = _T_8509 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8512 = _T_8510 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8522 = _T_4860 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8523 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8525 = _T_8523 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8526 = _T_8522 | _T_8525; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8527 = _T_8526 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8529 = _T_8527 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8539 = _T_4861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8540 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8542 = _T_8540 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8543 = _T_8539 | _T_8542; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8544 = _T_8543 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8546 = _T_8544 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8556 = _T_4862 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8557 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8559 = _T_8557 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8560 = _T_8556 | _T_8559; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8561 = _T_8560 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8563 = _T_8561 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8573 = _T_4863 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8574 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8576 = _T_8574 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8577 = _T_8573 | _T_8576; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8578 = _T_8577 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8580 = _T_8578 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8590 = _T_4864 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8591 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8593 = _T_8591 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8594 = _T_8590 | _T_8593; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8595 = _T_8594 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8597 = _T_8595 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8607 = _T_4865 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8608 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8610 = _T_8608 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8611 = _T_8607 | _T_8610; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8612 = _T_8611 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8614 = _T_8612 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8624 = _T_4866 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8625 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8627 = _T_8625 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8628 = _T_8624 | _T_8627; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8629 = _T_8628 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8631 = _T_8629 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8641 = _T_4867 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8642 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8644 = _T_8642 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8645 = _T_8641 | _T_8644; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8646 = _T_8645 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8648 = _T_8646 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8658 = _T_4868 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8659 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8661 = _T_8659 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8662 = _T_8658 | _T_8661; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8663 = _T_8662 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8665 = _T_8663 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8675 = _T_4869 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8676 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8678 = _T_8676 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8679 = _T_8675 | _T_8678; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8680 = _T_8679 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8682 = _T_8680 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8692 = _T_4870 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8693 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8695 = _T_8693 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8696 = _T_8692 | _T_8695; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8697 = _T_8696 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8699 = _T_8697 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8709 = _T_4871 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8710 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8712 = _T_8710 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8713 = _T_8709 | _T_8712; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8714 = _T_8713 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8716 = _T_8714 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8726 = _T_4872 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8727 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8729 = _T_8727 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8730 = _T_8726 | _T_8729; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8731 = _T_8730 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8733 = _T_8731 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8743 = _T_4873 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8744 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8746 = _T_8744 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8747 = _T_8743 | _T_8746; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8748 = _T_8747 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8750 = _T_8748 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8760 = _T_4874 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8761 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8763 = _T_8761 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8764 = _T_8760 | _T_8763; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8765 = _T_8764 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8767 = _T_8765 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8777 = _T_4875 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8778 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8780 = _T_8778 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8781 = _T_8777 | _T_8780; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8782 = _T_8781 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8784 = _T_8782 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8794 = _T_4876 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8795 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8797 = _T_8795 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8798 = _T_8794 | _T_8797; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8799 = _T_8798 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8801 = _T_8799 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8811 = _T_4877 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8812 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8814 = _T_8812 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8815 = _T_8811 | _T_8814; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8816 = _T_8815 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8818 = _T_8816 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8828 = _T_4878 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8829 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8831 = _T_8829 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8832 = _T_8828 | _T_8831; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8833 = _T_8832 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8835 = _T_8833 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8845 = _T_4879 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8846 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8848 = _T_8846 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8849 = _T_8845 | _T_8848; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8850 = _T_8849 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8852 = _T_8850 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8862 = _T_4880 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8863 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8865 = _T_8863 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8866 = _T_8862 | _T_8865; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8867 = _T_8866 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8869 = _T_8867 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8879 = _T_4881 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8880 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8882 = _T_8880 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8883 = _T_8879 | _T_8882; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8884 = _T_8883 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8886 = _T_8884 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8896 = _T_4882 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8897 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8899 = _T_8897 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8900 = _T_8896 | _T_8899; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8901 = _T_8900 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8903 = _T_8901 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8913 = _T_4883 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8914 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8916 = _T_8914 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8917 = _T_8913 | _T_8916; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8918 = _T_8917 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8920 = _T_8918 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8930 = _T_4884 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8931 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8933 = _T_8931 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8934 = _T_8930 | _T_8933; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8935 = _T_8934 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8937 = _T_8935 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8947 = _T_4885 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8948 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8950 = _T_8948 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8951 = _T_8947 | _T_8950; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8952 = _T_8951 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8954 = _T_8952 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8964 = _T_4886 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8965 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8967 = _T_8965 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8968 = _T_8964 | _T_8967; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8969 = _T_8968 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8971 = _T_8969 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8981 = _T_4887 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8982 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_8984 = _T_8982 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_8985 = _T_8981 | _T_8984; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_8986 = _T_8985 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_8988 = _T_8986 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_8998 = _T_4888 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_8999 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_9001 = _T_8999 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9002 = _T_8998 | _T_9001; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9003 = _T_9002 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9005 = _T_9003 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9015 = _T_4889 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9016 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_9018 = _T_9016 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9019 = _T_9015 | _T_9018; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9020 = _T_9019 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9022 = _T_9020 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9032 = _T_4890 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9033 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 757:102]
  wire  _T_9035 = _T_9033 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9036 = _T_9032 | _T_9035; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9037 = _T_9036 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9039 = _T_9037 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9049 = _T_4859 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9052 = _T_8506 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9053 = _T_9049 | _T_9052; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9054 = _T_9053 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9056 = _T_9054 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9066 = _T_4860 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9069 = _T_8523 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9070 = _T_9066 | _T_9069; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9071 = _T_9070 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9073 = _T_9071 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9083 = _T_4861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9086 = _T_8540 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9087 = _T_9083 | _T_9086; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9088 = _T_9087 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9090 = _T_9088 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9100 = _T_4862 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9103 = _T_8557 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9104 = _T_9100 | _T_9103; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9105 = _T_9104 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9107 = _T_9105 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9117 = _T_4863 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9120 = _T_8574 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9121 = _T_9117 | _T_9120; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9122 = _T_9121 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9124 = _T_9122 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9134 = _T_4864 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9137 = _T_8591 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9138 = _T_9134 | _T_9137; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9139 = _T_9138 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9141 = _T_9139 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9151 = _T_4865 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9154 = _T_8608 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9155 = _T_9151 | _T_9154; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9156 = _T_9155 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9158 = _T_9156 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9168 = _T_4866 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9171 = _T_8625 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9172 = _T_9168 | _T_9171; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9173 = _T_9172 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9175 = _T_9173 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9185 = _T_4867 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9188 = _T_8642 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9189 = _T_9185 | _T_9188; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9190 = _T_9189 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9192 = _T_9190 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9202 = _T_4868 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9205 = _T_8659 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9206 = _T_9202 | _T_9205; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9207 = _T_9206 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9209 = _T_9207 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9219 = _T_4869 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9222 = _T_8676 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9223 = _T_9219 | _T_9222; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9224 = _T_9223 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9226 = _T_9224 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9236 = _T_4870 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9239 = _T_8693 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9240 = _T_9236 | _T_9239; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9241 = _T_9240 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9243 = _T_9241 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9253 = _T_4871 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9256 = _T_8710 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9257 = _T_9253 | _T_9256; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9258 = _T_9257 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9260 = _T_9258 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9270 = _T_4872 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9273 = _T_8727 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9274 = _T_9270 | _T_9273; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9275 = _T_9274 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9277 = _T_9275 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9287 = _T_4873 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9290 = _T_8744 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9291 = _T_9287 | _T_9290; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9292 = _T_9291 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9294 = _T_9292 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9304 = _T_4874 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9307 = _T_8761 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9308 = _T_9304 | _T_9307; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9309 = _T_9308 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9311 = _T_9309 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9321 = _T_4875 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9324 = _T_8778 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9325 = _T_9321 | _T_9324; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9326 = _T_9325 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9328 = _T_9326 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9338 = _T_4876 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9341 = _T_8795 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9342 = _T_9338 | _T_9341; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9343 = _T_9342 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9345 = _T_9343 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9355 = _T_4877 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9358 = _T_8812 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9359 = _T_9355 | _T_9358; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9360 = _T_9359 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9362 = _T_9360 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9372 = _T_4878 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9375 = _T_8829 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9376 = _T_9372 | _T_9375; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9377 = _T_9376 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9379 = _T_9377 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9389 = _T_4879 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9392 = _T_8846 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9393 = _T_9389 | _T_9392; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9394 = _T_9393 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9396 = _T_9394 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9406 = _T_4880 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9409 = _T_8863 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9410 = _T_9406 | _T_9409; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9411 = _T_9410 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9413 = _T_9411 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9423 = _T_4881 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9426 = _T_8880 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9427 = _T_9423 | _T_9426; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9428 = _T_9427 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9430 = _T_9428 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9440 = _T_4882 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9443 = _T_8897 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9444 = _T_9440 | _T_9443; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9445 = _T_9444 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9447 = _T_9445 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9457 = _T_4883 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9460 = _T_8914 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9461 = _T_9457 | _T_9460; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9462 = _T_9461 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9464 = _T_9462 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9474 = _T_4884 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9477 = _T_8931 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9478 = _T_9474 | _T_9477; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9479 = _T_9478 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9481 = _T_9479 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9491 = _T_4885 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9494 = _T_8948 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9495 = _T_9491 | _T_9494; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9496 = _T_9495 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9498 = _T_9496 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9508 = _T_4886 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9511 = _T_8965 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9512 = _T_9508 | _T_9511; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9513 = _T_9512 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9515 = _T_9513 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9525 = _T_4887 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9528 = _T_8982 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9529 = _T_9525 | _T_9528; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9530 = _T_9529 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9532 = _T_9530 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9542 = _T_4888 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9545 = _T_8999 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9546 = _T_9542 | _T_9545; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9547 = _T_9546 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9549 = _T_9547 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9559 = _T_4889 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9562 = _T_9016 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9563 = _T_9559 | _T_9562; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9564 = _T_9563 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9566 = _T_9564 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_9576 = _T_4890 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 757:59]
  wire  _T_9579 = _T_9033 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 757:124]
  wire  _T_9580 = _T_9576 | _T_9579; // @[el2_ifu_mem_ctl.scala 757:81]
  wire  _T_9581 = _T_9580 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 757:147]
  wire  _T_9583 = _T_9581 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 757:165]
  wire  _T_10385 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 812:63]
  wire  _T_10386 = _T_10385 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 812:85]
  wire [1:0] _T_10388 = _T_10386 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10395; // @[el2_ifu_mem_ctl.scala 817:57]
  reg  _T_10396; // @[el2_ifu_mem_ctl.scala 818:56]
  reg  _T_10397; // @[el2_ifu_mem_ctl.scala 819:59]
  wire  _T_10398 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 820:80]
  wire  _T_10399 = ifu_bus_arvalid_ff & _T_10398; // @[el2_ifu_mem_ctl.scala 820:78]
  wire  _T_10400 = _T_10399 & miss_pending; // @[el2_ifu_mem_ctl.scala 820:100]
  reg  _T_10401; // @[el2_ifu_mem_ctl.scala 820:58]
  reg  _T_10402; // @[el2_ifu_mem_ctl.scala 821:58]
  wire  _T_10405 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 828:71]
  wire  _T_10407 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 828:124]
  wire  _T_10409 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 829:50]
  wire  _T_10411 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 829:103]
  wire [3:0] _T_10414 = {_T_10405,_T_10407,_T_10409,_T_10411}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 831:53]
  reg  _T_10423; // @[Reg.scala 27:20]
  rvclkhdr rvclkhdr ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_io_l1clk),
    .io_clk(rvclkhdr_io_clk),
    .io_en(rvclkhdr_io_en),
    .io_scan_mode(rvclkhdr_io_scan_mode)
  );
  rvclkhdr rvclkhdr_1 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_1_io_l1clk),
    .io_clk(rvclkhdr_1_io_clk),
    .io_en(rvclkhdr_1_io_en),
    .io_scan_mode(rvclkhdr_1_io_scan_mode)
  );
  rvclkhdr rvclkhdr_2 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_2_io_l1clk),
    .io_clk(rvclkhdr_2_io_clk),
    .io_en(rvclkhdr_2_io_en),
    .io_scan_mode(rvclkhdr_2_io_scan_mode)
  );
  rvclkhdr rvclkhdr_3 ( // @[el2_lib.scala 461:22]
    .io_l1clk(rvclkhdr_3_io_l1clk),
    .io_clk(rvclkhdr_3_io_clk),
    .io_en(rvclkhdr_3_io_en),
    .io_scan_mode(rvclkhdr_3_io_scan_mode)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 329:26]
  assign io_ifu_ic_mb_empty = _T_328 | _T_231; // @[el2_ifu_mem_ctl.scala 328:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 192:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3952; // @[el2_ifu_mem_ctl.scala 700:21]
  assign io_ifu_pmu_ic_miss = _T_10395; // @[el2_ifu_mem_ctl.scala 817:22]
  assign io_ifu_pmu_ic_hit = _T_10396; // @[el2_ifu_mem_ctl.scala 818:21]
  assign io_ifu_pmu_bus_error = _T_10397; // @[el2_ifu_mem_ctl.scala 819:24]
  assign io_ifu_pmu_bus_busy = _T_10401; // @[el2_ifu_mem_ctl.scala 820:23]
  assign io_ifu_pmu_bus_trxn = _T_10402; // @[el2_ifu_mem_ctl.scala 821:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 142:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 141:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 136:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 140:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 138:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 151:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 144:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 135:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 143:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 152:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 561:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2574; // @[el2_ifu_mem_ctl.scala 562:19]
  assign io_ifu_axi_araddr = _T_2576 & _T_2578; // @[el2_ifu_mem_ctl.scala 563:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 566:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 564:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 567:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 565:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 145:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 568:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 659:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 657:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 661:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 652:20]
  assign io_iccm_ready = _T_2672 & _T_2666; // @[el2_ifu_mem_ctl.scala 631:17]
  assign io_ic_rw_addr = _T_340 | _T_341; // @[el2_ifu_mem_ctl.scala 338:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_3938; // @[el2_ifu_mem_ctl.scala 699:15]
  assign io_ic_rd_en = _T_3930 | _T_3935; // @[el2_ifu_mem_ctl.scala 690:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 345:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 345:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 346:23]
  assign io_ifu_ic_debug_rd_data = _T_1211; // @[el2_ifu_mem_ctl.scala 354:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 824:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 826:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 827:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 825:25]
  assign io_ic_debug_way = _T_10414[1:0]; // @[el2_ifu_mem_ctl.scala 828:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10388; // @[el2_ifu_mem_ctl.scala 812:19]
  assign io_iccm_rw_addr = _T_3076 ? io_dma_mem_addr[15:1] : _T_3083; // @[el2_ifu_mem_ctl.scala 663:19]
  assign io_iccm_wren = _T_2676 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 633:16]
  assign io_iccm_rden = _T_2680 | _T_2681; // @[el2_ifu_mem_ctl.scala 634:16]
  assign io_iccm_wr_data = _T_3058 ? _T_3059 : _T_3066; // @[el2_ifu_mem_ctl.scala 640:19]
  assign io_iccm_wr_size = _T_2686 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 636:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 289:15]
  assign io_ic_access_fault_f = _T_2459 & _T_319; // @[el2_ifu_mem_ctl.scala 386:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1273; // @[el2_ifu_mem_ctl.scala 387:29]
  assign io_iccm_rd_ecc_single_err = _T_3875 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 676:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 677:29]
  assign io_ic_error_start = _T_1199 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 348:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 190:24]
  assign io_ic_fetch_val_f = {_T_1281,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 390:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 383:16]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[el2_ifu_mem_ctl.scala 380:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 381:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10423; // @[el2_ifu_mem_ctl.scala 835:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2464; // @[el2_ifu_mem_ctl.scala 480:27]
  assign io_iccm_correction_state = _T_2492 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 515:28 el2_ifu_mem_ctl.scala 528:32 el2_ifu_mem_ctl.scala 535:32 el2_ifu_mem_ctl.scala 542:32]
  assign rvclkhdr_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_io_en = ic_debug_rd_en_ff; // @[el2_lib.scala 463:16]
  assign rvclkhdr_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_1_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_1_io_en = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_lib.scala 463:16]
  assign rvclkhdr_1_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_2_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_2_io_en = _T_2 | scnd_miss_req; // @[el2_lib.scala 463:16]
  assign rvclkhdr_2_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
  assign rvclkhdr_3_io_clk = clock; // @[el2_lib.scala 462:17]
  assign rvclkhdr_3_io_en = _T_309 | io_dec_tlu_force_halt; // @[el2_lib.scala 463:16]
  assign rvclkhdr_3_io_scan_mode = io_scan_mode; // @[el2_lib.scala 464:23]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1211 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_443[6:0];
  _RAND_444 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_446[2:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_449[0:0];
  _RAND_450 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_450[38:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_453[2:0];
  _RAND_454 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_454[0:0];
  _RAND_455 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_455[63:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_456[13:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_458[13:0];
  _RAND_459 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_459[6:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way_status_new_ff = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  ic_valid_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10395 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10396 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10397 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10401 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10402 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_10423 = _RAND_469[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_3986) begin
      way_status_out_0 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_3991) begin
      way_status_out_1 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_3996) begin
      way_status_out_2 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4001) begin
      way_status_out_3 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4006) begin
      way_status_out_4 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4011) begin
      way_status_out_5 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4016) begin
      way_status_out_6 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4021) begin
      way_status_out_7 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4026) begin
      way_status_out_8 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4031) begin
      way_status_out_9 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4036) begin
      way_status_out_10 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4041) begin
      way_status_out_11 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4046) begin
      way_status_out_12 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4051) begin
      way_status_out_13 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4056) begin
      way_status_out_14 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4061) begin
      way_status_out_15 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4066) begin
      way_status_out_16 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4071) begin
      way_status_out_17 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4076) begin
      way_status_out_18 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4081) begin
      way_status_out_19 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4086) begin
      way_status_out_20 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4091) begin
      way_status_out_21 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4096) begin
      way_status_out_22 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4101) begin
      way_status_out_23 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4106) begin
      way_status_out_24 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4111) begin
      way_status_out_25 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4116) begin
      way_status_out_26 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4121) begin
      way_status_out_27 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4126) begin
      way_status_out_28 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4131) begin
      way_status_out_29 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4136) begin
      way_status_out_30 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4141) begin
      way_status_out_31 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4146) begin
      way_status_out_32 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4151) begin
      way_status_out_33 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4156) begin
      way_status_out_34 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4161) begin
      way_status_out_35 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4166) begin
      way_status_out_36 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4171) begin
      way_status_out_37 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4176) begin
      way_status_out_38 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4181) begin
      way_status_out_39 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4186) begin
      way_status_out_40 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4191) begin
      way_status_out_41 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4196) begin
      way_status_out_42 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4201) begin
      way_status_out_43 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4206) begin
      way_status_out_44 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4211) begin
      way_status_out_45 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4216) begin
      way_status_out_46 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4221) begin
      way_status_out_47 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4226) begin
      way_status_out_48 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4231) begin
      way_status_out_49 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4236) begin
      way_status_out_50 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4241) begin
      way_status_out_51 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4246) begin
      way_status_out_52 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4251) begin
      way_status_out_53 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4256) begin
      way_status_out_54 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4261) begin
      way_status_out_55 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4266) begin
      way_status_out_56 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4271) begin
      way_status_out_57 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4276) begin
      way_status_out_58 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4281) begin
      way_status_out_59 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4286) begin
      way_status_out_60 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4291) begin
      way_status_out_61 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4296) begin
      way_status_out_62 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4301) begin
      way_status_out_63 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4306) begin
      way_status_out_64 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4311) begin
      way_status_out_65 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4316) begin
      way_status_out_66 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4321) begin
      way_status_out_67 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4326) begin
      way_status_out_68 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4331) begin
      way_status_out_69 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4336) begin
      way_status_out_70 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4341) begin
      way_status_out_71 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4346) begin
      way_status_out_72 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4351) begin
      way_status_out_73 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4356) begin
      way_status_out_74 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4361) begin
      way_status_out_75 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4366) begin
      way_status_out_76 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4371) begin
      way_status_out_77 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4376) begin
      way_status_out_78 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4381) begin
      way_status_out_79 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4386) begin
      way_status_out_80 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4391) begin
      way_status_out_81 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4396) begin
      way_status_out_82 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4401) begin
      way_status_out_83 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4406) begin
      way_status_out_84 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4411) begin
      way_status_out_85 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4416) begin
      way_status_out_86 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4421) begin
      way_status_out_87 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4426) begin
      way_status_out_88 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4431) begin
      way_status_out_89 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4436) begin
      way_status_out_90 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4441) begin
      way_status_out_91 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4446) begin
      way_status_out_92 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4451) begin
      way_status_out_93 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4456) begin
      way_status_out_94 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4461) begin
      way_status_out_95 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4466) begin
      way_status_out_96 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4471) begin
      way_status_out_97 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4476) begin
      way_status_out_98 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4481) begin
      way_status_out_99 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4486) begin
      way_status_out_100 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4491) begin
      way_status_out_101 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4496) begin
      way_status_out_102 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4501) begin
      way_status_out_103 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4506) begin
      way_status_out_104 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4511) begin
      way_status_out_105 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4516) begin
      way_status_out_106 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4521) begin
      way_status_out_107 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4526) begin
      way_status_out_108 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4531) begin
      way_status_out_109 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4536) begin
      way_status_out_110 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4541) begin
      way_status_out_111 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4546) begin
      way_status_out_112 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4551) begin
      way_status_out_113 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4556) begin
      way_status_out_114 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4561) begin
      way_status_out_115 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4566) begin
      way_status_out_116 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4571) begin
      way_status_out_117 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4576) begin
      way_status_out_118 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4581) begin
      way_status_out_119 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4586) begin
      way_status_out_120 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4591) begin
      way_status_out_121 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4596) begin
      way_status_out_122 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4601) begin
      way_status_out_123 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4606) begin
      way_status_out_124 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4611) begin
      way_status_out_125 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4616) begin
      way_status_out_126 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4621) begin
      way_status_out_127 <= way_status_new_ff;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5792) begin
      ic_tag_valid_out_1_0 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5809) begin
      ic_tag_valid_out_1_1 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5826) begin
      ic_tag_valid_out_1_2 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5843) begin
      ic_tag_valid_out_1_3 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5860) begin
      ic_tag_valid_out_1_4 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5877) begin
      ic_tag_valid_out_1_5 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5894) begin
      ic_tag_valid_out_1_6 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5911) begin
      ic_tag_valid_out_1_7 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5928) begin
      ic_tag_valid_out_1_8 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5945) begin
      ic_tag_valid_out_1_9 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5962) begin
      ic_tag_valid_out_1_10 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5979) begin
      ic_tag_valid_out_1_11 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5996) begin
      ic_tag_valid_out_1_12 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_6013) begin
      ic_tag_valid_out_1_13 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_6030) begin
      ic_tag_valid_out_1_14 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_6047) begin
      ic_tag_valid_out_1_15 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_6064) begin
      ic_tag_valid_out_1_16 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_6081) begin
      ic_tag_valid_out_1_17 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6098) begin
      ic_tag_valid_out_1_18 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6115) begin
      ic_tag_valid_out_1_19 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6132) begin
      ic_tag_valid_out_1_20 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6149) begin
      ic_tag_valid_out_1_21 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6166) begin
      ic_tag_valid_out_1_22 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6183) begin
      ic_tag_valid_out_1_23 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6200) begin
      ic_tag_valid_out_1_24 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6217) begin
      ic_tag_valid_out_1_25 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6234) begin
      ic_tag_valid_out_1_26 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6251) begin
      ic_tag_valid_out_1_27 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6268) begin
      ic_tag_valid_out_1_28 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6285) begin
      ic_tag_valid_out_1_29 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6302) begin
      ic_tag_valid_out_1_30 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6319) begin
      ic_tag_valid_out_1_31 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6880) begin
      ic_tag_valid_out_1_32 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6897) begin
      ic_tag_valid_out_1_33 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6914) begin
      ic_tag_valid_out_1_34 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6931) begin
      ic_tag_valid_out_1_35 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6948) begin
      ic_tag_valid_out_1_36 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6965) begin
      ic_tag_valid_out_1_37 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6982) begin
      ic_tag_valid_out_1_38 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6999) begin
      ic_tag_valid_out_1_39 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_7016) begin
      ic_tag_valid_out_1_40 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_7033) begin
      ic_tag_valid_out_1_41 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_7050) begin
      ic_tag_valid_out_1_42 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_7067) begin
      ic_tag_valid_out_1_43 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_7084) begin
      ic_tag_valid_out_1_44 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_7101) begin
      ic_tag_valid_out_1_45 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_7118) begin
      ic_tag_valid_out_1_46 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_7135) begin
      ic_tag_valid_out_1_47 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7152) begin
      ic_tag_valid_out_1_48 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7169) begin
      ic_tag_valid_out_1_49 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7186) begin
      ic_tag_valid_out_1_50 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7203) begin
      ic_tag_valid_out_1_51 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7220) begin
      ic_tag_valid_out_1_52 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7237) begin
      ic_tag_valid_out_1_53 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7254) begin
      ic_tag_valid_out_1_54 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7271) begin
      ic_tag_valid_out_1_55 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7288) begin
      ic_tag_valid_out_1_56 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7305) begin
      ic_tag_valid_out_1_57 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7322) begin
      ic_tag_valid_out_1_58 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7339) begin
      ic_tag_valid_out_1_59 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7356) begin
      ic_tag_valid_out_1_60 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7373) begin
      ic_tag_valid_out_1_61 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7390) begin
      ic_tag_valid_out_1_62 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7407) begin
      ic_tag_valid_out_1_63 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7968) begin
      ic_tag_valid_out_1_64 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7985) begin
      ic_tag_valid_out_1_65 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_8002) begin
      ic_tag_valid_out_1_66 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_8019) begin
      ic_tag_valid_out_1_67 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_8036) begin
      ic_tag_valid_out_1_68 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_8053) begin
      ic_tag_valid_out_1_69 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_8070) begin
      ic_tag_valid_out_1_70 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_8087) begin
      ic_tag_valid_out_1_71 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_8104) begin
      ic_tag_valid_out_1_72 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_8121) begin
      ic_tag_valid_out_1_73 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_8138) begin
      ic_tag_valid_out_1_74 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_8155) begin
      ic_tag_valid_out_1_75 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_8172) begin
      ic_tag_valid_out_1_76 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_8189) begin
      ic_tag_valid_out_1_77 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_8206) begin
      ic_tag_valid_out_1_78 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8223) begin
      ic_tag_valid_out_1_79 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8240) begin
      ic_tag_valid_out_1_80 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8257) begin
      ic_tag_valid_out_1_81 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8274) begin
      ic_tag_valid_out_1_82 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8291) begin
      ic_tag_valid_out_1_83 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8308) begin
      ic_tag_valid_out_1_84 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8325) begin
      ic_tag_valid_out_1_85 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8342) begin
      ic_tag_valid_out_1_86 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8359) begin
      ic_tag_valid_out_1_87 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8376) begin
      ic_tag_valid_out_1_88 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8393) begin
      ic_tag_valid_out_1_89 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8410) begin
      ic_tag_valid_out_1_90 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8427) begin
      ic_tag_valid_out_1_91 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8444) begin
      ic_tag_valid_out_1_92 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8461) begin
      ic_tag_valid_out_1_93 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8478) begin
      ic_tag_valid_out_1_94 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8495) begin
      ic_tag_valid_out_1_95 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_9056) begin
      ic_tag_valid_out_1_96 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_9073) begin
      ic_tag_valid_out_1_97 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_9090) begin
      ic_tag_valid_out_1_98 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_9107) begin
      ic_tag_valid_out_1_99 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_9124) begin
      ic_tag_valid_out_1_100 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_9141) begin
      ic_tag_valid_out_1_101 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_9158) begin
      ic_tag_valid_out_1_102 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_9175) begin
      ic_tag_valid_out_1_103 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_9192) begin
      ic_tag_valid_out_1_104 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_9209) begin
      ic_tag_valid_out_1_105 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_9226) begin
      ic_tag_valid_out_1_106 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_9243) begin
      ic_tag_valid_out_1_107 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_9260) begin
      ic_tag_valid_out_1_108 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9277) begin
      ic_tag_valid_out_1_109 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9294) begin
      ic_tag_valid_out_1_110 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9311) begin
      ic_tag_valid_out_1_111 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9328) begin
      ic_tag_valid_out_1_112 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9345) begin
      ic_tag_valid_out_1_113 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9362) begin
      ic_tag_valid_out_1_114 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9379) begin
      ic_tag_valid_out_1_115 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9396) begin
      ic_tag_valid_out_1_116 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9413) begin
      ic_tag_valid_out_1_117 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9430) begin
      ic_tag_valid_out_1_118 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9447) begin
      ic_tag_valid_out_1_119 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9464) begin
      ic_tag_valid_out_1_120 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9481) begin
      ic_tag_valid_out_1_121 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9498) begin
      ic_tag_valid_out_1_122 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9515) begin
      ic_tag_valid_out_1_123 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9532) begin
      ic_tag_valid_out_1_124 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9549) begin
      ic_tag_valid_out_1_125 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9566) begin
      ic_tag_valid_out_1_126 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9583) begin
      ic_tag_valid_out_1_127 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5248) begin
      ic_tag_valid_out_0_0 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5265) begin
      ic_tag_valid_out_0_1 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5282) begin
      ic_tag_valid_out_0_2 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5299) begin
      ic_tag_valid_out_0_3 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5316) begin
      ic_tag_valid_out_0_4 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5333) begin
      ic_tag_valid_out_0_5 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5350) begin
      ic_tag_valid_out_0_6 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5367) begin
      ic_tag_valid_out_0_7 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5384) begin
      ic_tag_valid_out_0_8 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5401) begin
      ic_tag_valid_out_0_9 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5418) begin
      ic_tag_valid_out_0_10 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5435) begin
      ic_tag_valid_out_0_11 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5452) begin
      ic_tag_valid_out_0_12 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5469) begin
      ic_tag_valid_out_0_13 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5486) begin
      ic_tag_valid_out_0_14 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5503) begin
      ic_tag_valid_out_0_15 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5520) begin
      ic_tag_valid_out_0_16 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5537) begin
      ic_tag_valid_out_0_17 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5554) begin
      ic_tag_valid_out_0_18 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5571) begin
      ic_tag_valid_out_0_19 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5588) begin
      ic_tag_valid_out_0_20 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5605) begin
      ic_tag_valid_out_0_21 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5622) begin
      ic_tag_valid_out_0_22 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5639) begin
      ic_tag_valid_out_0_23 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5656) begin
      ic_tag_valid_out_0_24 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5673) begin
      ic_tag_valid_out_0_25 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5690) begin
      ic_tag_valid_out_0_26 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5707) begin
      ic_tag_valid_out_0_27 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5724) begin
      ic_tag_valid_out_0_28 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5741) begin
      ic_tag_valid_out_0_29 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5758) begin
      ic_tag_valid_out_0_30 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5775) begin
      ic_tag_valid_out_0_31 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6336) begin
      ic_tag_valid_out_0_32 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6353) begin
      ic_tag_valid_out_0_33 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6370) begin
      ic_tag_valid_out_0_34 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6387) begin
      ic_tag_valid_out_0_35 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6404) begin
      ic_tag_valid_out_0_36 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6421) begin
      ic_tag_valid_out_0_37 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6438) begin
      ic_tag_valid_out_0_38 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6455) begin
      ic_tag_valid_out_0_39 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6472) begin
      ic_tag_valid_out_0_40 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6489) begin
      ic_tag_valid_out_0_41 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6506) begin
      ic_tag_valid_out_0_42 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6523) begin
      ic_tag_valid_out_0_43 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6540) begin
      ic_tag_valid_out_0_44 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6557) begin
      ic_tag_valid_out_0_45 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6574) begin
      ic_tag_valid_out_0_46 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6591) begin
      ic_tag_valid_out_0_47 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6608) begin
      ic_tag_valid_out_0_48 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6625) begin
      ic_tag_valid_out_0_49 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6642) begin
      ic_tag_valid_out_0_50 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6659) begin
      ic_tag_valid_out_0_51 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6676) begin
      ic_tag_valid_out_0_52 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6693) begin
      ic_tag_valid_out_0_53 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6710) begin
      ic_tag_valid_out_0_54 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6727) begin
      ic_tag_valid_out_0_55 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6744) begin
      ic_tag_valid_out_0_56 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6761) begin
      ic_tag_valid_out_0_57 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6778) begin
      ic_tag_valid_out_0_58 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6795) begin
      ic_tag_valid_out_0_59 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6812) begin
      ic_tag_valid_out_0_60 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6829) begin
      ic_tag_valid_out_0_61 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6846) begin
      ic_tag_valid_out_0_62 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6863) begin
      ic_tag_valid_out_0_63 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7424) begin
      ic_tag_valid_out_0_64 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7441) begin
      ic_tag_valid_out_0_65 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7458) begin
      ic_tag_valid_out_0_66 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7475) begin
      ic_tag_valid_out_0_67 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7492) begin
      ic_tag_valid_out_0_68 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7509) begin
      ic_tag_valid_out_0_69 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7526) begin
      ic_tag_valid_out_0_70 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7543) begin
      ic_tag_valid_out_0_71 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7560) begin
      ic_tag_valid_out_0_72 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7577) begin
      ic_tag_valid_out_0_73 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7594) begin
      ic_tag_valid_out_0_74 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7611) begin
      ic_tag_valid_out_0_75 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7628) begin
      ic_tag_valid_out_0_76 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7645) begin
      ic_tag_valid_out_0_77 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7662) begin
      ic_tag_valid_out_0_78 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7679) begin
      ic_tag_valid_out_0_79 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7696) begin
      ic_tag_valid_out_0_80 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7713) begin
      ic_tag_valid_out_0_81 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7730) begin
      ic_tag_valid_out_0_82 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7747) begin
      ic_tag_valid_out_0_83 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7764) begin
      ic_tag_valid_out_0_84 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7781) begin
      ic_tag_valid_out_0_85 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7798) begin
      ic_tag_valid_out_0_86 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7815) begin
      ic_tag_valid_out_0_87 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7832) begin
      ic_tag_valid_out_0_88 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7849) begin
      ic_tag_valid_out_0_89 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7866) begin
      ic_tag_valid_out_0_90 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7883) begin
      ic_tag_valid_out_0_91 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7900) begin
      ic_tag_valid_out_0_92 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7917) begin
      ic_tag_valid_out_0_93 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7934) begin
      ic_tag_valid_out_0_94 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7951) begin
      ic_tag_valid_out_0_95 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8512) begin
      ic_tag_valid_out_0_96 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8529) begin
      ic_tag_valid_out_0_97 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8546) begin
      ic_tag_valid_out_0_98 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8563) begin
      ic_tag_valid_out_0_99 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8580) begin
      ic_tag_valid_out_0_100 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8597) begin
      ic_tag_valid_out_0_101 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8614) begin
      ic_tag_valid_out_0_102 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8631) begin
      ic_tag_valid_out_0_103 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8648) begin
      ic_tag_valid_out_0_104 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8665) begin
      ic_tag_valid_out_0_105 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8682) begin
      ic_tag_valid_out_0_106 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8699) begin
      ic_tag_valid_out_0_107 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8716) begin
      ic_tag_valid_out_0_108 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8733) begin
      ic_tag_valid_out_0_109 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8750) begin
      ic_tag_valid_out_0_110 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8767) begin
      ic_tag_valid_out_0_111 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8784) begin
      ic_tag_valid_out_0_112 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8801) begin
      ic_tag_valid_out_0_113 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8818) begin
      ic_tag_valid_out_0_114 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8835) begin
      ic_tag_valid_out_0_115 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8852) begin
      ic_tag_valid_out_0_116 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8869) begin
      ic_tag_valid_out_0_117 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8886) begin
      ic_tag_valid_out_0_118 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8903) begin
      ic_tag_valid_out_0_119 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8920) begin
      ic_tag_valid_out_0_120 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8937) begin
      ic_tag_valid_out_0_121 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8954) begin
      ic_tag_valid_out_0_122 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8971) begin
      ic_tag_valid_out_0_123 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8988) begin
      ic_tag_valid_out_0_124 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_9005) begin
      ic_tag_valid_out_0_125 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_9022) begin
      ic_tag_valid_out_0_126 <= _T_5238;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_9039) begin
      ic_tag_valid_out_0_127 <= _T_5238;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2566) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2680;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2467) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2469) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2479) begin
        perr_state <= 3'h0;
      end else if (_T_2482) begin
        if (_T_2484) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2488) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2492) begin
        err_stop_state <= 2'h1;
      end else if (_T_2497) begin
        if (_T_2499) begin
          err_stop_state <= 2'h0;
        end else if (_T_2520) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2524) begin
        if (_T_2499) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2541) begin
        if (_T_2545) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1370;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_3961) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1410;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3896;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3070;
    end else begin
      iccm_dma_rdata_temp <= _T_3071;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3892;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3961) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_3964) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_10373) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3964) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10423 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10423 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge rvclkhdr_2_io_l1clk) begin
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10395 <= 1'h0;
    end else begin
      _T_10395 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10396 <= 1'h0;
    end else begin
      _T_10396 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10397 <= 1'h0;
    end else begin
      _T_10397 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10401 <= 1'h0;
    end else begin
      _T_10401 <= _T_10400;
    end
    if (reset) begin
      _T_10402 <= 1'h0;
    end else begin
      _T_10402 <= bus_cmd_sent;
    end
  end
  always @(posedge rvclkhdr_3_io_l1clk) begin
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_231) begin
      bus_rd_addr_count <= imb_ff[4:2];
    end else if (scnd_miss_req_q) begin
      bus_rd_addr_count <= imb_scnd_ff[4:2];
    end else if (bus_cmd_sent) begin
      bus_rd_addr_count <= _T_2613;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (bus_cmd_beat_en) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
  end
  always @(posedge rvclkhdr_1_io_l1clk) begin
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
  end
  always @(posedge rvclkhdr_io_l1clk) begin
    if (reset) begin
      _T_1211 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1211 <= {{5'd0}, _T_1210};
    end else begin
      _T_1211 <= io_ic_debug_rd_data;
    end
  end
endmodule
