typedef struct packed {
	bit [3:0]      BHT_ADDR_HI;
	bit [1:0]      BHT_ADDR_LO;
	bit [10:0]     BHT_ARRAY_DEPTH;
	bit            BHT_GHR_HASH_1;
	bit [3:0]      BHT_GHR_SIZE;
	bit [11:0]     BHT_SIZE;
	bit [4:0]      BTB_ADDR_HI;
	bit [1:0]      BTB_ADDR_LO;
	bit [8:0]      BTB_ARRAY_DEPTH;
	bit            BTB_BTAG_FOLD;
	bit [3:0]      BTB_BTAG_SIZE;
	bit            BTB_FOLD2_INDEX_HASH;
	bit [4:0]      BTB_INDEX1_HI;
	bit [4:0]      BTB_INDEX1_LO;
	bit [4:0]      BTB_INDEX2_HI;
	bit [4:0]      BTB_INDEX2_LO;
	bit [4:0]      BTB_INDEX3_HI;
	bit [4:0]      BTB_INDEX3_LO;
	bit [9:0]      BTB_SIZE;
	bit            BUILD_AHB_LITE;
	bit            BUILD_AXI4;
	bit            BUILD_AXI_NATIVE;
	bit [1:0]      BUS_PRTY_DEFAULT;
	bit [31:0]     DATA_ACCESS_ADDR0;
	bit [31:0]     DATA_ACCESS_ADDR1;
	bit [31:0]     DATA_ACCESS_ADDR2;
	bit [31:0]     DATA_ACCESS_ADDR3;
	bit [31:0]     DATA_ACCESS_ADDR4;
	bit [31:0]     DATA_ACCESS_ADDR5;
	bit [31:0]     DATA_ACCESS_ADDR6;
	bit [31:0]     DATA_ACCESS_ADDR7;
	bit            DATA_ACCESS_ENABLE0;
	bit            DATA_ACCESS_ENABLE1;
	bit            DATA_ACCESS_ENABLE2;
	bit            DATA_ACCESS_ENABLE3;
	bit            DATA_ACCESS_ENABLE4;
	bit            DATA_ACCESS_ENABLE5;
	bit            DATA_ACCESS_ENABLE6;
	bit            DATA_ACCESS_ENABLE7;
	bit [31:0]     DATA_ACCESS_MASK0;
	bit [31:0]     DATA_ACCESS_MASK1;
	bit [31:0]     DATA_ACCESS_MASK2;
	bit [31:0]     DATA_ACCESS_MASK3;
	bit [31:0]     DATA_ACCESS_MASK4;
	bit [31:0]     DATA_ACCESS_MASK5;
	bit [31:0]     DATA_ACCESS_MASK6;
	bit [31:0]     DATA_ACCESS_MASK7;
	bit [2:0]      DCCM_BANK_BITS;
	bit [4:0]      DCCM_BITS;
	bit [2:0]      DCCM_BYTE_WIDTH;
	bit [5:0]      DCCM_DATA_WIDTH;
	bit [2:0]      DCCM_ECC_WIDTH;
	bit            DCCM_ENABLE;
	bit [5:0]      DCCM_FDATA_WIDTH;
	bit [3:0]      DCCM_INDEX_BITS;
	bit [4:0]      DCCM_NUM_BANKS;
	bit [3:0]      DCCM_REGION;
	bit [31:0]     DCCM_SADR;
	bit [9:0]      DCCM_SIZE;
	bit [1:0]      DCCM_WIDTH_BITS;
	bit [2:0]      DMA_BUF_DEPTH;
	bit            DMA_BUS_ID;
	bit [1:0]      DMA_BUS_PRTY;
	bit [3:0]      DMA_BUS_TAG;
	bit            FAST_INTERRUPT_REDIRECT;
	bit            ICACHE_2BANKS;
	bit [2:0]      ICACHE_BANK_BITS;
	bit [2:0]      ICACHE_BANK_HI;
	bit [1:0]      ICACHE_BANK_LO;
	bit [3:0]      ICACHE_BANK_WIDTH;
	bit [2:0]      ICACHE_BANKS_WAY;
	bit [3:0]      ICACHE_BEAT_ADDR_HI;
	bit [3:0]      ICACHE_BEAT_BITS;
	bit [13:0]     ICACHE_DATA_DEPTH;
	bit [2:0]      ICACHE_DATA_INDEX_LO;
	bit [6:0]      ICACHE_DATA_WIDTH;
	bit            ICACHE_ECC;
	bit            ICACHE_ENABLE;
	bit [6:0]      ICACHE_FDATA_WIDTH;
	bit [4:0]      ICACHE_INDEX_HI;
	bit [6:0]      ICACHE_LN_SZ;
	bit [3:0]      ICACHE_NUM_BEATS;
	bit [2:0]      ICACHE_NUM_WAYS;
	bit            ICACHE_ONLY;
	bit [3:0]      ICACHE_SCND_LAST;
	bit [8:0]      ICACHE_SIZE;
	bit [2:0]      ICACHE_STATUS_BITS;
	bit [12:0]     ICACHE_TAG_DEPTH;
	bit [2:0]      ICACHE_TAG_INDEX_LO;
	bit [4:0]      ICACHE_TAG_LO;
	bit            ICACHE_WAYPACK;
	bit [2:0]      ICCM_BANK_BITS;
	bit [4:0]      ICCM_BANK_HI;
	bit [4:0]      ICCM_BANK_INDEX_LO;
	bit [4:0]      ICCM_BITS;
	bit            ICCM_ENABLE;
	bit            ICCM_ICACHE;
	bit [3:0]      ICCM_INDEX_BITS;
	bit [4:0]      ICCM_NUM_BANKS;
	bit            ICCM_ONLY;
	bit [3:0]      ICCM_REGION;
	bit [31:0]     ICCM_SADR;
	bit [9:0]      ICCM_SIZE;
	bit            IFU_BUS_ID;
	bit [1:0]      IFU_BUS_PRTY;
	bit [3:0]      IFU_BUS_TAG;
	bit [31:0]     INST_ACCESS_ADDR0;
	bit [31:0]     INST_ACCESS_ADDR1;
	bit [31:0]     INST_ACCESS_ADDR2;
	bit [31:0]     INST_ACCESS_ADDR3;
	bit [31:0]     INST_ACCESS_ADDR4;
	bit [31:0]     INST_ACCESS_ADDR5;
	bit [31:0]     INST_ACCESS_ADDR6;
	bit [31:0]     INST_ACCESS_ADDR7;
	bit            INST_ACCESS_ENABLE0;
	bit            INST_ACCESS_ENABLE1;
	bit            INST_ACCESS_ENABLE2;
	bit            INST_ACCESS_ENABLE3;
	bit            INST_ACCESS_ENABLE4;
	bit            INST_ACCESS_ENABLE5;
	bit            INST_ACCESS_ENABLE6;
	bit            INST_ACCESS_ENABLE7;
	bit [31:0]     INST_ACCESS_MASK0;
	bit [31:0]     INST_ACCESS_MASK1;
	bit [31:0]     INST_ACCESS_MASK2;
	bit [31:0]     INST_ACCESS_MASK3;
	bit [31:0]     INST_ACCESS_MASK4;
	bit [31:0]     INST_ACCESS_MASK5;
	bit [31:0]     INST_ACCESS_MASK6;
	bit [31:0]     INST_ACCESS_MASK7;
	bit            LOAD_TO_USE_PLUS1;
	bit            LSU2DMA;
	bit            LSU_BUS_ID;
	bit [1:0]      LSU_BUS_PRTY;
	bit [3:0]      LSU_BUS_TAG;
	bit [4:0]      LSU_NUM_NBLOAD;
	bit [2:0]      LSU_NUM_NBLOAD_WIDTH;
	bit [4:0]      LSU_SB_BITS;
	bit [3:0]      LSU_STBUF_DEPTH;
	bit            NO_ICCM_NO_ICACHE;
	bit            PIC_2CYCLE;
	bit [31:0]     PIC_BASE_ADDR;
	bit [4:0]      PIC_BITS;
	bit [3:0]      PIC_INT_WORDS;
	bit [3:0]      PIC_REGION;
	bit [8:0]      PIC_SIZE;
	bit [7:0]      PIC_TOTAL_INT;
	bit [8:0]      PIC_TOTAL_INT_PLUS1;
	bit [3:0]      RET_STACK_SIZE;
	bit            SB_BUS_ID;
	bit [1:0]      SB_BUS_PRTY;
	bit [3:0]      SB_BUS_TAG;
	bit            TIMER_LEGAL_EN;
} param_t;

