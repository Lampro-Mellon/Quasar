module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  input         io_ifu_axi_arready,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  input         io_ifu_axi_rvalid,
  output        io_ifu_axi_rready,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [63:0] _RAND_159;
  reg [63:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [63:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [63:0] _RAND_165;
  reg [63:0] _RAND_166;
  reg [63:0] _RAND_167;
  reg [63:0] _RAND_168;
  reg [63:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [63:0] _RAND_172;
  reg [63:0] _RAND_173;
  reg [63:0] _RAND_174;
  reg [63:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [95:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [63:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 178:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 311:36]
  wire  _T_308 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 312:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_308; // @[el2_ifu_mem_ctl.scala 312:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 244:30]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 180:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 299:34]
  wire [4:0] _GEN_463 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 652:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_463 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 652:53]
  wire [1:0] _GEN_464 = {{1'd0}, _T_308}; // @[el2_ifu_mem_ctl.scala 655:91]
  wire [1:0] _T_3063 = ic_fetch_val_shift_right[3:2] & _GEN_464; // @[el2_ifu_mem_ctl.scala 655:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 313:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 266:46]
  wire [1:0] _GEN_465 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 655:113]
  wire [1:0] _T_3064 = _T_3063 & _GEN_465; // @[el2_ifu_mem_ctl.scala 655:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 641:59]
  wire [1:0] _GEN_466 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 655:130]
  wire [1:0] _T_3065 = _T_3064 | _GEN_466; // @[el2_ifu_mem_ctl.scala 655:130]
  wire  _T_3066 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 655:154]
  wire [1:0] _GEN_467 = {{1'd0}, _T_3066}; // @[el2_ifu_mem_ctl.scala 655:152]
  wire [1:0] _T_3067 = _T_3065 & _GEN_467; // @[el2_ifu_mem_ctl.scala 655:152]
  wire [1:0] _T_3056 = ic_fetch_val_shift_right[1:0] & _GEN_464; // @[el2_ifu_mem_ctl.scala 655:91]
  wire [1:0] _T_3057 = _T_3056 & _GEN_465; // @[el2_ifu_mem_ctl.scala 655:113]
  wire [1:0] _T_3058 = _T_3057 | _GEN_466; // @[el2_ifu_mem_ctl.scala 655:130]
  wire [1:0] _T_3060 = _T_3058 & _GEN_467; // @[el2_ifu_mem_ctl.scala 655:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3067,_T_3060}; // @[Cat.scala 29:58]
  wire  _T_3167 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_3168 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_3169 = _T_3167 ^ _T_3168; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3177 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_3178 = ^_T_3177; // @[el2_lib.scala 301:83]
  wire  _T_3179 = io_iccm_rd_data_ecc[37] ^ _T_3178; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3186 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3194 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3186}; // @[el2_lib.scala 301:103]
  wire  _T_3195 = ^_T_3194; // @[el2_lib.scala 301:110]
  wire  _T_3196 = io_iccm_rd_data_ecc[36] ^ _T_3195; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3203 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3211 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3203}; // @[el2_lib.scala 301:130]
  wire  _T_3212 = ^_T_3211; // @[el2_lib.scala 301:137]
  wire  _T_3213 = io_iccm_rd_data_ecc[35] ^ _T_3212; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3222 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3231 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3222}; // @[el2_lib.scala 301:157]
  wire  _T_3232 = ^_T_3231; // @[el2_lib.scala 301:164]
  wire  _T_3233 = io_iccm_rd_data_ecc[34] ^ _T_3232; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3242 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3251 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3242}; // @[el2_lib.scala 301:184]
  wire  _T_3252 = ^_T_3251; // @[el2_lib.scala 301:191]
  wire  _T_3253 = io_iccm_rd_data_ecc[33] ^ _T_3252; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3262 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3271 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3262}; // @[el2_lib.scala 301:211]
  wire  _T_3272 = ^_T_3271; // @[el2_lib.scala 301:218]
  wire  _T_3273 = io_iccm_rd_data_ecc[32] ^ _T_3272; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3279 = {_T_3169,_T_3179,_T_3196,_T_3213,_T_3233,_T_3253,_T_3273}; // @[Cat.scala 29:58]
  wire  _T_3280 = _T_3279 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3281 = iccm_ecc_word_enable[0] & _T_3280; // @[el2_lib.scala 302:32]
  wire  _T_3283 = _T_3281 & _T_3279[6]; // @[el2_lib.scala 302:53]
  wire  _T_3552 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_3553 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_3554 = _T_3552 ^ _T_3553; // @[el2_lib.scala 301:35]
  wire [5:0] _T_3562 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_3563 = ^_T_3562; // @[el2_lib.scala 301:83]
  wire  _T_3564 = io_iccm_rd_data_ecc[76] ^ _T_3563; // @[el2_lib.scala 301:71]
  wire [6:0] _T_3571 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_3579 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3571}; // @[el2_lib.scala 301:103]
  wire  _T_3580 = ^_T_3579; // @[el2_lib.scala 301:110]
  wire  _T_3581 = io_iccm_rd_data_ecc[75] ^ _T_3580; // @[el2_lib.scala 301:98]
  wire [6:0] _T_3588 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_3596 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3588}; // @[el2_lib.scala 301:130]
  wire  _T_3597 = ^_T_3596; // @[el2_lib.scala 301:137]
  wire  _T_3598 = io_iccm_rd_data_ecc[74] ^ _T_3597; // @[el2_lib.scala 301:125]
  wire [8:0] _T_3607 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_3616 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3607}; // @[el2_lib.scala 301:157]
  wire  _T_3617 = ^_T_3616; // @[el2_lib.scala 301:164]
  wire  _T_3618 = io_iccm_rd_data_ecc[73] ^ _T_3617; // @[el2_lib.scala 301:152]
  wire [8:0] _T_3627 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_3636 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3627}; // @[el2_lib.scala 301:184]
  wire  _T_3637 = ^_T_3636; // @[el2_lib.scala 301:191]
  wire  _T_3638 = io_iccm_rd_data_ecc[72] ^ _T_3637; // @[el2_lib.scala 301:179]
  wire [8:0] _T_3647 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_3656 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3647}; // @[el2_lib.scala 301:211]
  wire  _T_3657 = ^_T_3656; // @[el2_lib.scala 301:218]
  wire  _T_3658 = io_iccm_rd_data_ecc[71] ^ _T_3657; // @[el2_lib.scala 301:206]
  wire [6:0] _T_3664 = {_T_3554,_T_3564,_T_3581,_T_3598,_T_3618,_T_3638,_T_3658}; // @[Cat.scala 29:58]
  wire  _T_3665 = _T_3664 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_3666 = iccm_ecc_word_enable[1] & _T_3665; // @[el2_lib.scala 302:32]
  wire  _T_3668 = _T_3666 & _T_3664[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_3283,_T_3668}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 183:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 619:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 184:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 185:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 465:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 185:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 185:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 185:72]
  wire  _T_2434 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2439 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2459 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 515:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 381:42]
  wire  _T_2461 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 515:79]
  wire  _T_2462 = _T_2459 | _T_2461; // @[el2_ifu_mem_ctl.scala 515:56]
  wire  _T_2463 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 515:122]
  wire  _T_2464 = ~_T_2463; // @[el2_ifu_mem_ctl.scala 515:101]
  wire  _T_2465 = _T_2462 & _T_2464; // @[el2_ifu_mem_ctl.scala 515:99]
  wire  _T_2466 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2480 = io_ifu_fetch_val[0] & _T_308; // @[el2_ifu_mem_ctl.scala 522:45]
  wire  _T_2481 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 522:69]
  wire  _T_2482 = _T_2480 & _T_2481; // @[el2_ifu_mem_ctl.scala 522:67]
  wire  _T_2483 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = _T_2466 ? _T_2482 : _T_2483; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2439 ? _T_2465 : _GEN_54; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2434 ? 1'h0 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 185:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 186:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 186:65]
  wire  _T_218 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 274:37]
  wire  _T_219 = ~_T_218; // @[el2_ifu_mem_ctl.scala 274:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 687:53]
  wire  _T_220 = _T_219 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 274:41]
  wire  _T_198 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 265:48]
  wire  _T_199 = ifc_fetch_req_f & _T_198; // @[el2_ifu_mem_ctl.scala 265:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 315:42]
  wire  _T_200 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 265:69]
  wire  fetch_req_icache_f = _T_199 & _T_200; // @[el2_ifu_mem_ctl.scala 265:67]
  wire  _T_221 = _T_220 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 274:59]
  wire  _T_222 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 274:82]
  wire  _T_223 = _T_221 & _T_222; // @[el2_ifu_mem_ctl.scala 274:80]
  wire  ic_act_miss_f = _T_223 & _T_200; // @[el2_ifu_mem_ctl.scala 274:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 535:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 576:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 603:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 301:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 584:56]
  wire  _T_2583 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 601:69]
  wire  _T_2584 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 601:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2583 : _T_2584; // @[el2_ifu_mem_ctl.scala 601:28]
  wire  _T_2530 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 580:68]
  wire  _T_2531 = ic_act_miss_f | _T_2530; // @[el2_ifu_mem_ctl.scala 580:48]
  wire  bus_reset_data_beat_cnt = _T_2531 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 580:91]
  wire  _T_2527 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 579:50]
  wire  _T_2528 = bus_ifu_wr_en_ff & _T_2527; // @[el2_ifu_mem_ctl.scala 579:48]
  wire  _T_2529 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 579:72]
  wire  bus_inc_data_beat_cnt = _T_2528 & _T_2529; // @[el2_ifu_mem_ctl.scala 579:70]
  wire [2:0] _T_2535 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 583:115]
  wire [2:0] _T_2537 = bus_inc_data_beat_cnt ? _T_2535 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2532 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 581:32]
  wire  _T_2533 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 581:57]
  wire  bus_hold_data_beat_cnt = _T_2532 & _T_2533; // @[el2_ifu_mem_ctl.scala 581:55]
  wire [2:0] _T_2538 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2537 | _T_2538; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 186:111]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 186:85]
  wire  _T_17 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 187:39]
  wire  _T_25 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_27 = ic_act_miss_f & _T_308; // @[el2_ifu_mem_ctl.scala 193:43]
  wire [2:0] _T_29 = _T_27 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 193:27]
  wire  _T_32 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 417:45]
  wire  _T_2099 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 438:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 394:60]
  wire  _T_2130 = _T_2099 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2103 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2131 = _T_2103 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2138 = _T_2130 | _T_2131; // @[Mux.scala 27:72]
  wire  _T_2107 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2132 = _T_2107 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2139 = _T_2138 | _T_2132; // @[Mux.scala 27:72]
  wire  _T_2111 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2133 = _T_2111 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2140 = _T_2139 | _T_2133; // @[Mux.scala 27:72]
  wire  _T_2115 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2134 = _T_2115 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2141 = _T_2140 | _T_2134; // @[Mux.scala 27:72]
  wire  _T_2119 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2135 = _T_2119 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2142 = _T_2141 | _T_2135; // @[Mux.scala 27:72]
  wire  _T_2123 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2136 = _T_2123 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2143 = _T_2142 | _T_2136; // @[Mux.scala 27:72]
  wire  _T_2127 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 438:127]
  wire  _T_2137 = _T_2127 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2143 | _T_2137; // @[Mux.scala 27:72]
  wire  _T_2185 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 440:69]
  wire  _T_2186 = ic_miss_buff_data_valid_bypass_index & _T_2185; // @[el2_ifu_mem_ctl.scala 440:67]
  wire  _T_2188 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 440:91]
  wire  _T_2189 = _T_2186 & _T_2188; // @[el2_ifu_mem_ctl.scala 440:89]
  wire  _T_2194 = _T_2186 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 441:65]
  wire  _T_2195 = _T_2189 | _T_2194; // @[el2_ifu_mem_ctl.scala 440:112]
  wire  _T_2197 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 442:43]
  wire  _T_2200 = _T_2197 & _T_2188; // @[el2_ifu_mem_ctl.scala 442:65]
  wire  _T_2201 = _T_2195 | _T_2200; // @[el2_ifu_mem_ctl.scala 441:88]
  wire  _T_2205 = _T_2197 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 443:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 420:75]
  wire  _T_2145 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2169 = _T_2145 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2148 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2170 = _T_2148 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2177 = _T_2169 | _T_2170; // @[Mux.scala 27:72]
  wire  _T_2151 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2171 = _T_2151 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2178 = _T_2177 | _T_2171; // @[Mux.scala 27:72]
  wire  _T_2154 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2172 = _T_2154 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2179 = _T_2178 | _T_2172; // @[Mux.scala 27:72]
  wire  _T_2157 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2173 = _T_2157 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2180 = _T_2179 | _T_2173; // @[Mux.scala 27:72]
  wire  _T_2160 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2174 = _T_2160 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2181 = _T_2180 | _T_2174; // @[Mux.scala 27:72]
  wire  _T_2163 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2175 = _T_2163 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2182 = _T_2181 | _T_2175; // @[Mux.scala 27:72]
  wire  _T_2166 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 439:110]
  wire  _T_2176 = _T_2166 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2182 | _T_2176; // @[Mux.scala 27:72]
  wire  _T_2206 = _T_2205 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 443:87]
  wire  _T_2207 = _T_2201 | _T_2206; // @[el2_ifu_mem_ctl.scala 442:88]
  wire  _T_2217 = _T_2189 & _T_2127; // @[el2_ifu_mem_ctl.scala 444:87]
  wire  miss_buff_hit_unq_f = _T_2207 | _T_2217; // @[el2_ifu_mem_ctl.scala 443:131]
  wire  _T_2232 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 449:55]
  wire  _T_2233 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 449:87]
  wire  _T_2234 = _T_2232 | _T_2233; // @[el2_ifu_mem_ctl.scala 449:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2234; // @[el2_ifu_mem_ctl.scala 449:41]
  wire  _T_2218 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 446:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 302:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 437:51]
  wire  _T_2219 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 446:68]
  wire  _T_2220 = miss_buff_hit_unq_f & _T_2219; // @[el2_ifu_mem_ctl.scala 446:66]
  wire  stream_hit_f = _T_2218 & _T_2220; // @[el2_ifu_mem_ctl.scala 446:43]
  wire  _T_206 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 269:35]
  wire  _T_207 = _T_206 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 269:52]
  wire  ic_byp_hit_f = _T_207 & miss_pending; // @[el2_ifu_mem_ctl.scala 269:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 586:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 613:35]
  wire  _T_33 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 196:112]
  wire  _T_34 = last_data_recieved_ff | _T_33; // @[el2_ifu_mem_ctl.scala 196:92]
  wire  _T_35 = ic_byp_hit_f & _T_34; // @[el2_ifu_mem_ctl.scala 196:66]
  wire  _T_36 = _T_35 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 196:126]
  wire  _T_37 = io_dec_tlu_force_halt | _T_36; // @[el2_ifu_mem_ctl.scala 196:51]
  wire  _T_39 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 197:30]
  wire  _T_40 = ic_byp_hit_f & _T_39; // @[el2_ifu_mem_ctl.scala 197:27]
  wire  _T_41 = _T_40 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 197:53]
  wire  _T_43 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 198:16]
  wire  _T_45 = _T_43 & _T_308; // @[el2_ifu_mem_ctl.scala 198:30]
  wire  _T_47 = _T_45 & _T_33; // @[el2_ifu_mem_ctl.scala 198:52]
  wire  _T_48 = _T_47 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 198:85]
  wire  _T_51 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 199:51]
  wire  _T_52 = _T_33 & _T_51; // @[el2_ifu_mem_ctl.scala 199:49]
  wire  _T_54 = ic_byp_hit_f | bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 200:34]
  wire  _T_56 = _T_54 & _T_308; // @[el2_ifu_mem_ctl.scala 200:54]
  wire  _T_58 = ~_T_33; // @[el2_ifu_mem_ctl.scala 200:78]
  wire  _T_59 = _T_56 & _T_58; // @[el2_ifu_mem_ctl.scala 200:76]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 189:52]
  wire  _T_60 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 200:112]
  wire  _T_61 = _T_59 & _T_60; // @[el2_ifu_mem_ctl.scala 200:110]
  wire  _T_63 = _T_61 & _T_51; // @[el2_ifu_mem_ctl.scala 200:134]
  wire  _T_71 = _T_47 & _T_51; // @[el2_ifu_mem_ctl.scala 201:100]
  wire  _T_73 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 202:44]
  wire  _T_76 = _T_73 & _T_58; // @[el2_ifu_mem_ctl.scala 202:68]
  wire [2:0] _T_78 = _T_76 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 202:22]
  wire [2:0] _T_79 = _T_71 ? 3'h0 : _T_78; // @[el2_ifu_mem_ctl.scala 201:20]
  wire [2:0] _T_80 = _T_63 ? 3'h6 : _T_79; // @[el2_ifu_mem_ctl.scala 200:18]
  wire [2:0] _T_81 = _T_52 ? 3'h0 : _T_80; // @[el2_ifu_mem_ctl.scala 199:16]
  wire [2:0] _T_82 = _T_48 ? 3'h1 : _T_81; // @[el2_ifu_mem_ctl.scala 198:14]
  wire [2:0] _T_83 = _T_41 ? 3'h3 : _T_82; // @[el2_ifu_mem_ctl.scala 197:12]
  wire [2:0] _T_84 = _T_37 ? 3'h0 : _T_83; // @[el2_ifu_mem_ctl.scala 196:27]
  wire  _T_93 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_97 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2229 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 448:60]
  wire  _T_2230 = _T_2229 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 448:92]
  wire  stream_eol_f = _T_2230 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_99 = _T_73 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 210:72]
  wire  _T_102 = _T_99 & _T_58; // @[el2_ifu_mem_ctl.scala 210:87]
  wire  _T_104 = _T_102 & _T_2529; // @[el2_ifu_mem_ctl.scala 210:122]
  wire [2:0] _T_106 = _T_104 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 210:27]
  wire  _T_112 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_115 = io_exu_flush_final & _T_58; // @[el2_ifu_mem_ctl.scala 214:48]
  wire  _T_117 = _T_115 & _T_2529; // @[el2_ifu_mem_ctl.scala 214:82]
  wire [2:0] _T_119 = _T_117 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 214:27]
  wire  _T_123 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_227 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 275:28]
  wire  _T_228 = _T_227 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 275:42]
  wire  _T_229 = _T_228 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 275:60]
  wire  _T_230 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 275:94]
  wire  _T_231 = _T_229 & _T_230; // @[el2_ifu_mem_ctl.scala 275:81]
  wire  _T_234 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 276:39]
  wire  _T_235 = _T_231 & _T_234; // @[el2_ifu_mem_ctl.scala 275:111]
  wire  _T_237 = _T_235 & _T_51; // @[el2_ifu_mem_ctl.scala 276:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 329:51]
  wire  _T_238 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 276:116]
  wire  _T_239 = _T_237 & _T_238; // @[el2_ifu_mem_ctl.scala 276:114]
  wire  ic_miss_under_miss_f = _T_239 & _T_200; // @[el2_ifu_mem_ctl.scala 276:132]
  wire  _T_126 = ic_miss_under_miss_f & _T_58; // @[el2_ifu_mem_ctl.scala 218:50]
  wire  _T_128 = _T_126 & _T_2529; // @[el2_ifu_mem_ctl.scala 218:84]
  wire  _T_247 = _T_221 & _T_230; // @[el2_ifu_mem_ctl.scala 277:85]
  wire  _T_250 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 278:39]
  wire  _T_251 = _T_250 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 278:91]
  wire  ic_ignore_2nd_miss_f = _T_247 & _T_251; // @[el2_ifu_mem_ctl.scala 277:117]
  wire  _T_132 = ic_ignore_2nd_miss_f & _T_58; // @[el2_ifu_mem_ctl.scala 219:35]
  wire  _T_134 = _T_132 & _T_2529; // @[el2_ifu_mem_ctl.scala 219:69]
  wire [2:0] _T_136 = _T_134 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 219:12]
  wire [2:0] _T_137 = _T_128 ? 3'h5 : _T_136; // @[el2_ifu_mem_ctl.scala 218:27]
  wire  _T_142 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_145 = _T_33 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 224:12]
  wire [2:0] _T_146 = io_exu_flush_final ? _T_145 : 3'h1; // @[el2_ifu_mem_ctl.scala 223:62]
  wire [2:0] _T_147 = io_dec_tlu_force_halt ? 3'h0 : _T_146; // @[el2_ifu_mem_ctl.scala 223:27]
  wire  _T_151 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_145 : 3'h0; // @[el2_ifu_mem_ctl.scala 228:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 228:27]
  wire [2:0] _GEN_0 = _T_151 ? _T_156 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_142 ? _T_147 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_123 ? _T_137 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_112 ? _T_119 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_97 ? _T_106 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_93 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_32 ? _T_84 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_25 ? _T_29 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_18 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 187:71]
  wire  _T_19 = _T_17 | _T_18; // @[el2_ifu_mem_ctl.scala 187:55]
  wire  _T_20 = uncacheable_miss_ff >> _T_19; // @[el2_ifu_mem_ctl.scala 187:26]
  wire  _T_22 = ~_T_20; // @[el2_ifu_mem_ctl.scala 187:5]
  wire  _T_23 = _T_16 & _T_22; // @[el2_ifu_mem_ctl.scala 186:116]
  wire  scnd_miss_req_in = _T_23 & _T_308; // @[el2_ifu_mem_ctl.scala 187:89]
  wire  _T_31 = ic_act_miss_f & _T_2529; // @[el2_ifu_mem_ctl.scala 194:38]
  wire  _T_85 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 203:46]
  wire  _T_86 = _T_85 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 203:67]
  wire  _T_87 = _T_86 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 203:82]
  wire  _T_89 = _T_87 | _T_33; // @[el2_ifu_mem_ctl.scala 203:105]
  wire  _T_91 = bus_ifu_wr_en_ff & _T_51; // @[el2_ifu_mem_ctl.scala 203:158]
  wire  _T_92 = _T_89 | _T_91; // @[el2_ifu_mem_ctl.scala 203:138]
  wire  _T_94 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 207:43]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:59]
  wire  _T_96 = _T_95 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 207:74]
  wire  _T_110 = _T_99 | _T_33; // @[el2_ifu_mem_ctl.scala 211:84]
  wire  _T_111 = _T_110 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 211:118]
  wire  _T_121 = io_exu_flush_final | _T_33; // @[el2_ifu_mem_ctl.scala 215:43]
  wire  _T_122 = _T_121 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 215:76]
  wire  _T_139 = _T_33 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 220:55]
  wire  _T_140 = _T_139 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 220:78]
  wire  _T_141 = _T_140 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 220:101]
  wire  _T_149 = _T_33 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 225:55]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _GEN_1 = _T_151 & _T_150; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_142 ? _T_150 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_123 ? _T_141 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_112 ? _T_122 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_97 ? _T_111 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_93 ? _T_96 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_32 ? _T_92 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_25 ? _T_31 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_165 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 245:95]
  wire  _T_166 = _T_2232 & _T_165; // @[el2_ifu_mem_ctl.scala 245:93]
  wire  crit_wd_byp_ok_ff = _T_2233 | _T_166; // @[el2_ifu_mem_ctl.scala 245:58]
  wire  _T_169 = miss_pending & _T_58; // @[el2_ifu_mem_ctl.scala 246:36]
  wire  _T_171 = _T_2232 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 246:106]
  wire  _T_172 = ~_T_171; // @[el2_ifu_mem_ctl.scala 246:72]
  wire  _T_173 = _T_169 & _T_172; // @[el2_ifu_mem_ctl.scala 246:70]
  wire  _T_175 = _T_2232 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 247:57]
  wire  _T_176 = ~_T_175; // @[el2_ifu_mem_ctl.scala 247:23]
  wire  _T_177 = _T_173 & _T_176; // @[el2_ifu_mem_ctl.scala 246:128]
  wire  _T_178 = _T_177 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 247:77]
  wire  _T_179 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 248:36]
  wire  _T_180 = miss_pending & _T_179; // @[el2_ifu_mem_ctl.scala 248:19]
  wire  sel_hold_imb = _T_178 | _T_180; // @[el2_ifu_mem_ctl.scala 247:93]
  wire  _T_182 = _T_17 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 250:57]
  wire  sel_hold_imb_scnd = _T_182 & _T_165; // @[el2_ifu_mem_ctl.scala 250:81]
  reg [6:0] _T_5108; // @[el2_ifu_mem_ctl.scala 715:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_5108[5:0]; // @[el2_ifu_mem_ctl.scala 714:27]
  wire [6:0] _GEN_472 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 711:121]
  wire  _T_4973 = _GEN_472 == 7'h7f; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4975 = _T_4973 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4464; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_4464[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_473 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4976 = _T_4975 & _GEN_473; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4969 = _GEN_472 == 7'h7e; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4971 = _T_4969 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4460; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_4460[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_475 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4972 = _T_4971 & _GEN_475; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4965 = _GEN_472 == 7'h7d; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4967 = _T_4965 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4456; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_4456[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_477 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4968 = _T_4967 & _GEN_477; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4961 = _GEN_472 == 7'h7c; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4963 = _T_4961 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4452; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_4452[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_479 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4964 = _T_4963 & _GEN_479; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4957 = _GEN_472 == 7'h7b; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4959 = _T_4957 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4448; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_4448[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_481 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4960 = _T_4959 & _GEN_481; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4953 = _GEN_472 == 7'h7a; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4955 = _T_4953 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4444; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_4444[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_483 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4956 = _T_4955 & _GEN_483; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4949 = _GEN_472 == 7'h79; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4951 = _T_4949 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4440; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_4440[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_485 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4952 = _T_4951 & _GEN_485; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4945 = _GEN_472 == 7'h78; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4947 = _T_4945 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4436; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_4436[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_487 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4948 = _T_4947 & _GEN_487; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4941 = _GEN_472 == 7'h77; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4943 = _T_4941 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4432; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_4432[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_489 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4944 = _T_4943 & _GEN_489; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4937 = _GEN_472 == 7'h76; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4939 = _T_4937 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4428; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_4428[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_491 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4940 = _T_4939 & _GEN_491; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [59:0] _T_4985 = {_T_4976,_T_4972,_T_4968,_T_4964,_T_4960,_T_4956,_T_4952,_T_4948,_T_4944,_T_4940}; // @[Cat.scala 29:58]
  wire  _T_4933 = _GEN_472 == 7'h75; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4935 = _T_4933 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4424; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_4424[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_493 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4936 = _T_4935 & _GEN_493; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4929 = _GEN_472 == 7'h74; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4931 = _T_4929 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4420; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_4420[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_495 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4932 = _T_4931 & _GEN_495; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4925 = _GEN_472 == 7'h73; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4927 = _T_4925 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4416; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_4416[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_497 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4928 = _T_4927 & _GEN_497; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4921 = _GEN_472 == 7'h72; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4923 = _T_4921 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4412; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_4412[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_499 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4924 = _T_4923 & _GEN_499; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4917 = _GEN_472 == 7'h71; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4919 = _T_4917 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4408; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_4408[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_501 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4920 = _T_4919 & _GEN_501; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4913 = _GEN_472 == 7'h70; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4915 = _T_4913 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4404; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_4404[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_503 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4916 = _T_4915 & _GEN_503; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4909 = _GEN_472 == 7'h6f; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4911 = _T_4909 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4400; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_4400[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_505 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4912 = _T_4911 & _GEN_505; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4905 = _GEN_472 == 7'h6e; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4907 = _T_4905 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4396; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_4396[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_507 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4908 = _T_4907 & _GEN_507; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4901 = _GEN_472 == 7'h6d; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4903 = _T_4901 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4392; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_4392[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_509 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4904 = _T_4903 & _GEN_509; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [113:0] _T_4994 = {_T_4985,_T_4936,_T_4932,_T_4928,_T_4924,_T_4920,_T_4916,_T_4912,_T_4908,_T_4904}; // @[Cat.scala 29:58]
  wire  _T_4897 = _GEN_472 == 7'h6c; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4899 = _T_4897 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4388; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_4388[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_511 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4900 = _T_4899 & _GEN_511; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4893 = _GEN_472 == 7'h6b; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4895 = _T_4893 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4384; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_4384[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_513 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4896 = _T_4895 & _GEN_513; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4889 = _GEN_472 == 7'h6a; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4891 = _T_4889 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4380; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_4380[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_515 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4892 = _T_4891 & _GEN_515; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4885 = _GEN_472 == 7'h69; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4887 = _T_4885 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4376; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_4376[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_517 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4888 = _T_4887 & _GEN_517; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4881 = _GEN_472 == 7'h68; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4883 = _T_4881 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4372; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_4372[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_519 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4884 = _T_4883 & _GEN_519; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4877 = _GEN_472 == 7'h67; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4879 = _T_4877 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4368; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_4368[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_521 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4880 = _T_4879 & _GEN_521; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4873 = _GEN_472 == 7'h66; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4875 = _T_4873 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4364; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_4364[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_523 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4876 = _T_4875 & _GEN_523; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4869 = _GEN_472 == 7'h65; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4871 = _T_4869 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4360; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_4360[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_525 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4872 = _T_4871 & _GEN_525; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4865 = _GEN_472 == 7'h64; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4867 = _T_4865 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4356; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_4356[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_527 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4868 = _T_4867 & _GEN_527; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [167:0] _T_5003 = {_T_4994,_T_4900,_T_4896,_T_4892,_T_4888,_T_4884,_T_4880,_T_4876,_T_4872,_T_4868}; // @[Cat.scala 29:58]
  wire  _T_4861 = _GEN_472 == 7'h63; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4863 = _T_4861 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4352; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_4352[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_529 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4864 = _T_4863 & _GEN_529; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4857 = _GEN_472 == 7'h62; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4859 = _T_4857 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4348; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_4348[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_531 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4860 = _T_4859 & _GEN_531; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4853 = _GEN_472 == 7'h61; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4855 = _T_4853 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4344; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_4344[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_533 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4856 = _T_4855 & _GEN_533; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4849 = _GEN_472 == 7'h60; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4851 = _T_4849 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4340; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_4340[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_535 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4852 = _T_4851 & _GEN_535; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4845 = _GEN_472 == 7'h5f; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4847 = _T_4845 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4336; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_4336[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_537 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4848 = _T_4847 & _GEN_537; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4841 = _GEN_472 == 7'h5e; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4843 = _T_4841 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4332; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_4332[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_539 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4844 = _T_4843 & _GEN_539; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4837 = _GEN_472 == 7'h5d; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4839 = _T_4837 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4328; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_4328[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_541 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4840 = _T_4839 & _GEN_541; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4833 = _GEN_472 == 7'h5c; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4835 = _T_4833 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4324; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_4324[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_543 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4836 = _T_4835 & _GEN_543; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4829 = _GEN_472 == 7'h5b; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4831 = _T_4829 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4320; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_4320[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_545 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4832 = _T_4831 & _GEN_545; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [221:0] _T_5012 = {_T_5003,_T_4864,_T_4860,_T_4856,_T_4852,_T_4848,_T_4844,_T_4840,_T_4836,_T_4832}; // @[Cat.scala 29:58]
  wire  _T_4825 = _GEN_472 == 7'h5a; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4827 = _T_4825 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4316; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_4316[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_547 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4828 = _T_4827 & _GEN_547; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4821 = _GEN_472 == 7'h59; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4823 = _T_4821 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4312; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_4312[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_549 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4824 = _T_4823 & _GEN_549; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4817 = _GEN_472 == 7'h58; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4819 = _T_4817 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4308; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_4308[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_551 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4820 = _T_4819 & _GEN_551; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4813 = _GEN_472 == 7'h57; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4815 = _T_4813 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4304; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_4304[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_553 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4816 = _T_4815 & _GEN_553; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4809 = _GEN_472 == 7'h56; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4811 = _T_4809 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4300; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_4300[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_555 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4812 = _T_4811 & _GEN_555; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4805 = _GEN_472 == 7'h55; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4807 = _T_4805 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4296; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_4296[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_557 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4808 = _T_4807 & _GEN_557; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4801 = _GEN_472 == 7'h54; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4803 = _T_4801 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4292; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_4292[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_559 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4804 = _T_4803 & _GEN_559; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4797 = _GEN_472 == 7'h53; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4799 = _T_4797 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4288; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_4288[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_561 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4800 = _T_4799 & _GEN_561; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4793 = _GEN_472 == 7'h52; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4795 = _T_4793 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4284; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_4284[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_563 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4796 = _T_4795 & _GEN_563; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [275:0] _T_5021 = {_T_5012,_T_4828,_T_4824,_T_4820,_T_4816,_T_4812,_T_4808,_T_4804,_T_4800,_T_4796}; // @[Cat.scala 29:58]
  wire  _T_4789 = _GEN_472 == 7'h51; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4791 = _T_4789 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4280; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_4280[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_565 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4792 = _T_4791 & _GEN_565; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4785 = _GEN_472 == 7'h50; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4787 = _T_4785 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4276; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_4276[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_567 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4788 = _T_4787 & _GEN_567; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4781 = _GEN_472 == 7'h4f; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4783 = _T_4781 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4272; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_4272[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_569 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4784 = _T_4783 & _GEN_569; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4777 = _GEN_472 == 7'h4e; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4779 = _T_4777 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4268; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_4268[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_571 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4780 = _T_4779 & _GEN_571; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4773 = _GEN_472 == 7'h4d; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4775 = _T_4773 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4264; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_4264[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_573 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4776 = _T_4775 & _GEN_573; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4769 = _GEN_472 == 7'h4c; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4771 = _T_4769 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4260; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_4260[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_575 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4772 = _T_4771 & _GEN_575; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4765 = _GEN_472 == 7'h4b; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4767 = _T_4765 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4256; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_4256[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_577 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4768 = _T_4767 & _GEN_577; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4761 = _GEN_472 == 7'h4a; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4763 = _T_4761 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4252; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_4252[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_579 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4764 = _T_4763 & _GEN_579; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4757 = _GEN_472 == 7'h49; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4759 = _T_4757 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4248; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_4248[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_581 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4760 = _T_4759 & _GEN_581; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [329:0] _T_5030 = {_T_5021,_T_4792,_T_4788,_T_4784,_T_4780,_T_4776,_T_4772,_T_4768,_T_4764,_T_4760}; // @[Cat.scala 29:58]
  wire  _T_4753 = _GEN_472 == 7'h48; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4755 = _T_4753 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4244; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_4244[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_583 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4756 = _T_4755 & _GEN_583; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4749 = _GEN_472 == 7'h47; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4751 = _T_4749 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4240; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_4240[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_585 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4752 = _T_4751 & _GEN_585; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4745 = _GEN_472 == 7'h46; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4747 = _T_4745 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4236; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_4236[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_587 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4748 = _T_4747 & _GEN_587; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4741 = _GEN_472 == 7'h45; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4743 = _T_4741 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4232; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_4232[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_589 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4744 = _T_4743 & _GEN_589; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4737 = _GEN_472 == 7'h44; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4739 = _T_4737 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4228; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_4228[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_591 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4740 = _T_4739 & _GEN_591; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4733 = _GEN_472 == 7'h43; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4735 = _T_4733 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4224; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_4224[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_593 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4736 = _T_4735 & _GEN_593; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4729 = _GEN_472 == 7'h42; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4731 = _T_4729 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4220; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_4220[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_595 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4732 = _T_4731 & _GEN_595; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4725 = _GEN_472 == 7'h41; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4727 = _T_4725 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4216; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_4216[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_597 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4728 = _T_4727 & _GEN_597; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4721 = _GEN_472 == 7'h40; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4723 = _T_4721 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4212; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_4212[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_599 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4724 = _T_4723 & _GEN_599; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [383:0] _T_5039 = {_T_5030,_T_4756,_T_4752,_T_4748,_T_4744,_T_4740,_T_4736,_T_4732,_T_4728,_T_4724}; // @[Cat.scala 29:58]
  wire  _T_4717 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4719 = _T_4717 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4208; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_4208[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4720 = _T_4719 & _GEN_600; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4713 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4715 = _T_4713 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4204; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_4204[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4716 = _T_4715 & _GEN_601; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4709 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4711 = _T_4709 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4200; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_4200[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4712 = _T_4711 & _GEN_602; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4705 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4707 = _T_4705 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4196; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_4196[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4708 = _T_4707 & _GEN_603; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4701 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4703 = _T_4701 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4192; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_4192[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4704 = _T_4703 & _GEN_604; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4697 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4699 = _T_4697 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4188; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_4188[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4700 = _T_4699 & _GEN_605; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4693 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4695 = _T_4693 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4184; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_4184[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4696 = _T_4695 & _GEN_606; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4689 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4691 = _T_4689 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4180; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_4180[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4692 = _T_4691 & _GEN_607; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4685 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4687 = _T_4685 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4176; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_4176[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4688 = _T_4687 & _GEN_608; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [437:0] _T_5048 = {_T_5039,_T_4720,_T_4716,_T_4712,_T_4708,_T_4704,_T_4700,_T_4696,_T_4692,_T_4688}; // @[Cat.scala 29:58]
  wire  _T_4681 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4683 = _T_4681 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4172; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_4172[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4684 = _T_4683 & _GEN_609; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4677 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4679 = _T_4677 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4168; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_4168[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4680 = _T_4679 & _GEN_610; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4673 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4675 = _T_4673 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4164; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_4164[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4676 = _T_4675 & _GEN_611; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4669 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4671 = _T_4669 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4160; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_4160[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4672 = _T_4671 & _GEN_612; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4665 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4667 = _T_4665 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4156; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_4156[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4668 = _T_4667 & _GEN_613; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4661 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4663 = _T_4661 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4152; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_4152[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4664 = _T_4663 & _GEN_614; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4657 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4659 = _T_4657 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4148; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_4148[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4660 = _T_4659 & _GEN_615; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4653 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4655 = _T_4653 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4144; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_4144[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4656 = _T_4655 & _GEN_616; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4649 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4651 = _T_4649 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4140; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_4140[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4652 = _T_4651 & _GEN_617; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [491:0] _T_5057 = {_T_5048,_T_4684,_T_4680,_T_4676,_T_4672,_T_4668,_T_4664,_T_4660,_T_4656,_T_4652}; // @[Cat.scala 29:58]
  wire  _T_4645 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4647 = _T_4645 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4136; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_4136[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4648 = _T_4647 & _GEN_618; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4641 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4643 = _T_4641 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4132; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_4132[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4644 = _T_4643 & _GEN_619; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4637 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4639 = _T_4637 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4128; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_4128[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4640 = _T_4639 & _GEN_620; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4633 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4635 = _T_4633 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4124; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_4124[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4636 = _T_4635 & _GEN_621; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4629 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4631 = _T_4629 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4120; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_4120[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4632 = _T_4631 & _GEN_622; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4625 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4627 = _T_4625 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4116; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_4116[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4628 = _T_4627 & _GEN_623; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4621 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4623 = _T_4621 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4112; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_4112[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4624 = _T_4623 & _GEN_624; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4617 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4619 = _T_4617 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4108; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_4108[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4620 = _T_4619 & _GEN_625; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4613 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4615 = _T_4613 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4104; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_4104[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4616 = _T_4615 & _GEN_626; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [545:0] _T_5066 = {_T_5057,_T_4648,_T_4644,_T_4640,_T_4636,_T_4632,_T_4628,_T_4624,_T_4620,_T_4616}; // @[Cat.scala 29:58]
  wire  _T_4609 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4611 = _T_4609 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4100; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_4100[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4612 = _T_4611 & _GEN_627; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4605 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4607 = _T_4605 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4096; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_4096[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4608 = _T_4607 & _GEN_628; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4601 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4603 = _T_4601 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4092; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_4092[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4604 = _T_4603 & _GEN_629; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4597 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4599 = _T_4597 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4088; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_4088[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4600 = _T_4599 & _GEN_630; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4593 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4595 = _T_4593 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4084; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_4084[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4596 = _T_4595 & _GEN_631; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4589 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4591 = _T_4589 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4080; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_4080[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4592 = _T_4591 & _GEN_632; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4585 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4587 = _T_4585 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4076; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_4076[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4588 = _T_4587 & _GEN_633; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4581 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4583 = _T_4581 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4072; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_4072[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4584 = _T_4583 & _GEN_634; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4577 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4579 = _T_4577 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4068; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_4068[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4580 = _T_4579 & _GEN_635; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [599:0] _T_5075 = {_T_5066,_T_4612,_T_4608,_T_4604,_T_4600,_T_4596,_T_4592,_T_4588,_T_4584,_T_4580}; // @[Cat.scala 29:58]
  wire  _T_4573 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4575 = _T_4573 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4064; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_4064[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4576 = _T_4575 & _GEN_636; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4569 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4571 = _T_4569 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4060; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_4060[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4572 = _T_4571 & _GEN_637; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4565 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4567 = _T_4565 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4056; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_4056[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4568 = _T_4567 & _GEN_638; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4561 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4563 = _T_4561 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4052; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_4052[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4564 = _T_4563 & _GEN_639; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4557 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4559 = _T_4557 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4048; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_4048[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4560 = _T_4559 & _GEN_640; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4553 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4555 = _T_4553 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4044; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_4044[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4556 = _T_4555 & _GEN_641; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4549 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4551 = _T_4549 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4040; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_4040[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4552 = _T_4551 & _GEN_642; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4545 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4547 = _T_4545 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4036; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_4036[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4548 = _T_4547 & _GEN_643; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4541 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4543 = _T_4541 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4032; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_4032[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4544 = _T_4543 & _GEN_644; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [653:0] _T_5084 = {_T_5075,_T_4576,_T_4572,_T_4568,_T_4564,_T_4560,_T_4556,_T_4552,_T_4548,_T_4544}; // @[Cat.scala 29:58]
  wire  _T_4537 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4539 = _T_4537 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4028; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_4028[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4540 = _T_4539 & _GEN_645; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4533 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4535 = _T_4533 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4024; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_4024[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4536 = _T_4535 & _GEN_646; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4529 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4531 = _T_4529 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4020; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_4020[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4532 = _T_4531 & _GEN_647; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4525 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4527 = _T_4525 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4016; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_4016[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4528 = _T_4527 & _GEN_648; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4521 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4523 = _T_4521 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4012; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_4012[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4524 = _T_4523 & _GEN_649; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4517 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4519 = _T_4517 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4008; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_4008[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4520 = _T_4519 & _GEN_650; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4513 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4515 = _T_4513 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4004; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_4004[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4516 = _T_4515 & _GEN_651; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4509 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4511 = _T_4509 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_4000; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_4000[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4512 = _T_4511 & _GEN_652; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4505 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4507 = _T_4505 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3996; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_3996[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4508 = _T_4507 & _GEN_653; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [707:0] _T_5093 = {_T_5084,_T_4540,_T_4536,_T_4532,_T_4528,_T_4524,_T_4520,_T_4516,_T_4512,_T_4508}; // @[Cat.scala 29:58]
  wire  _T_4501 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4503 = _T_4501 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3992; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3992[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4504 = _T_4503 & _GEN_654; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4497 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4499 = _T_4497 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3988; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3988[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4500 = _T_4499 & _GEN_655; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4493 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4495 = _T_4493 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3984; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3984[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4496 = _T_4495 & _GEN_656; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4489 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4491 = _T_4489 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3980; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3980[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4492 = _T_4491 & _GEN_657; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4485 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4487 = _T_4485 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3976; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3976[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4488 = _T_4487 & _GEN_658; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4481 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4483 = _T_4481 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3972; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3972[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4484 = _T_4483 & _GEN_659; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4477 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4479 = _T_4477 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3968; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3968[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4480 = _T_4479 & _GEN_660; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4473 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4475 = _T_4473 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3964; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3964[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4476 = _T_4475 & _GEN_661; // @[el2_ifu_mem_ctl.scala 711:130]
  wire  _T_4469 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4471 = _T_4469 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3960; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3960[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4472 = _T_4471 & _GEN_662; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [761:0] _T_5102 = {_T_5093,_T_4504,_T_4500,_T_4496,_T_4492,_T_4488,_T_4484,_T_4480,_T_4476,_T_4472}; // @[Cat.scala 29:58]
  wire  _T_4465 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 711:121]
  wire [5:0] _T_4467 = _T_4465 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3956; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3956[0]; // @[el2_ifu_mem_ctl.scala 708:30 el2_ifu_mem_ctl.scala 710:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [5:0] _T_4468 = _T_4467 & _GEN_663; // @[el2_ifu_mem_ctl.scala 711:130]
  wire [767:0] _T_5103 = {_T_5102,_T_4468}; // @[Cat.scala 29:58]
  wire  way_status = _T_5103[0]; // @[el2_ifu_mem_ctl.scala 711:16]
  wire  _T_186 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 253:96]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 257:25]
  wire [2:0] _T_197 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_197; // @[el2_ifu_mem_ctl.scala 262:45]
  wire  _T_203 = _T_222 | _T_230; // @[el2_ifu_mem_ctl.scala 267:59]
  wire  _T_205 = _T_203 | _T_2218; // @[el2_ifu_mem_ctl.scala 267:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_205; // @[el2_ifu_mem_ctl.scala 267:41]
  wire  _T_210 = _T_218 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 273:39]
  wire  _T_212 = _T_210 & _T_186; // @[el2_ifu_mem_ctl.scala 273:60]
  wire  _T_216 = _T_212 & _T_203; // @[el2_ifu_mem_ctl.scala 273:78]
  wire  ic_act_hit_f = _T_216 & _T_238; // @[el2_ifu_mem_ctl.scala 273:126]
  wire  _T_253 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 280:31]
  wire  _T_254 = _T_253 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 280:46]
  wire  _T_255 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 280:94]
  wire  uncacheable_miss_in = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 281:84]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2604 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 609:48]
  wire  _T_2605 = _T_2604 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 609:52]
  wire  bus_ifu_wr_data_error_ff = _T_2605 & miss_pending; // @[el2_ifu_mem_ctl.scala 609:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 356:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 355:55]
  wire  _T_267 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 284:145]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 536:52]
  wire  _T_288 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 296:36]
  wire  _T_289 = miss_pending & _T_288; // @[el2_ifu_mem_ctl.scala 296:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 297:25]
  wire  _T_290 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 296:72]
  wire  reset_ic_in = _T_289 & _T_290; // @[el2_ifu_mem_ctl.scala 296:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 298:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 306:23]
  wire  _T_304 = _T_2232 & flush_final_f; // @[el2_ifu_mem_ctl.scala 310:87]
  wire  _T_305 = ~_T_304; // @[el2_ifu_mem_ctl.scala 310:55]
  wire  _T_306 = io_ifc_fetch_req_bf & _T_305; // @[el2_ifu_mem_ctl.scala 310:53]
  wire  stream_miss_f = stream_hit_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 447:83]
  wire  _T_307 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 310:106]
  wire  ifc_fetch_req_qual_bf = _T_306 & _T_307; // @[el2_ifu_mem_ctl.scala 310:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 316:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_314 = _T_230 | _T_2218; // @[el2_ifu_mem_ctl.scala 318:55]
  wire  _T_317 = _T_314 & _T_58; // @[el2_ifu_mem_ctl.scala 318:82]
  wire  _T_2238 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 452:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2238}; // @[Cat.scala 29:58]
  wire  _T_2239 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2263 = _T_2239 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2242 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2264 = _T_2242 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2271 = _T_2263 | _T_2264; // @[Mux.scala 27:72]
  wire  _T_2245 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2265 = _T_2245 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2272 = _T_2271 | _T_2265; // @[Mux.scala 27:72]
  wire  _T_2248 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2266 = _T_2248 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2273 = _T_2272 | _T_2266; // @[Mux.scala 27:72]
  wire  _T_2251 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2267 = _T_2251 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2274 = _T_2273 | _T_2267; // @[Mux.scala 27:72]
  wire  _T_2254 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2268 = _T_2254 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2275 = _T_2274 | _T_2268; // @[Mux.scala 27:72]
  wire  _T_2257 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2269 = _T_2257 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2276 = _T_2275 | _T_2269; // @[Mux.scala 27:72]
  wire  _T_2260 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 453:81]
  wire  _T_2270 = _T_2260 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2276 | _T_2270; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 454:46]
  wire  _T_321 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 322:35]
  wire  _T_323 = _T_321 & _T_51; // @[el2_ifu_mem_ctl.scala 322:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 606:61]
  wire  _T_2598 = ic_act_miss_f_delayed & _T_2233; // @[el2_ifu_mem_ctl.scala 607:53]
  wire  reset_tag_valid_for_miss = _T_2598 & _T_51; // @[el2_ifu_mem_ctl.scala 607:84]
  wire  sel_mb_addr = _T_323 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 322:79]
  wire [30:0] _T_328 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_330 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 324:37]
  wire [30:0] _T_331 = sel_mb_addr ? _T_328 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_332 = _T_330 ? ifu_fetch_addr_int_f : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_331 | _T_332; // @[Mux.scala 27:72]
  wire  _T_337 = _T_323 & last_beat; // @[el2_ifu_mem_ctl.scala 326:84]
  wire  _T_2592 = ~_T_2604; // @[el2_ifu_mem_ctl.scala 604:84]
  wire  _T_2593 = _T_91 & _T_2592; // @[el2_ifu_mem_ctl.scala 604:82]
  wire  bus_ifu_wr_en_ff_q = _T_2593 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 604:108]
  wire  sel_mb_status_addr = _T_337 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 326:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_328 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 327:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [7:0] _T_561 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_570 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_561}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_578 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_587 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_578}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_588 = {_T_587,_T_570}; // @[el2_lib.scala 348:27]
  wire  _T_589 = ^_T_588; // @[el2_lib.scala 348:34]
  wire [7:0] _T_596 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_605 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_596}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_613 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_622 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_613}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_623 = {_T_622,_T_605}; // @[el2_lib.scala 348:44]
  wire  _T_624 = ^_T_623; // @[el2_lib.scala 348:51]
  wire [7:0] _T_631 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_640 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_631}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_648 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_657 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_648}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_658 = {_T_657,_T_640}; // @[el2_lib.scala 348:61]
  wire  _T_659 = ^_T_658; // @[el2_lib.scala 348:68]
  wire [6:0] _T_665 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_673 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_665}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_680 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_689 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_680,_T_673}; // @[el2_lib.scala 348:78]
  wire  _T_690 = ^_T_689; // @[el2_lib.scala 348:85]
  wire [6:0] _T_696 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_704 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_696}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_711 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_720 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_711,_T_704}; // @[el2_lib.scala 348:95]
  wire  _T_721 = ^_T_720; // @[el2_lib.scala 348:102]
  wire [6:0] _T_727 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_735 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_727}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_751 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_711,_T_735}; // @[el2_lib.scala 348:112]
  wire  _T_752 = ^_T_751; // @[el2_lib.scala 348:119]
  wire [6:0] _T_758 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 348:129]
  wire  _T_759 = ^_T_758; // @[el2_lib.scala 348:136]
  wire [3:0] _T_2279 = {ifu_bus_rid_ff[2:1],_T_2238,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2280 = _T_2279 == 4'h0; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1286; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_0 = _T_1286[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2327 = _T_2280 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2283 = _T_2279 == 4'h1; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1288; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_1 = _T_1288[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2328 = _T_2283 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2343 = _T_2327 | _T_2328; // @[Mux.scala 27:72]
  wire  _T_2286 = _T_2279 == 4'h2; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1290; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_2 = _T_1290[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2329 = _T_2286 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2344 = _T_2343 | _T_2329; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2279 == 4'h3; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1292; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_3 = _T_1292[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2330 = _T_2289 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2345 = _T_2344 | _T_2330; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2279 == 4'h4; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1294; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_4 = _T_1294[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2331 = _T_2292 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2346 = _T_2345 | _T_2331; // @[Mux.scala 27:72]
  wire  _T_2295 = _T_2279 == 4'h5; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1296; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_5 = _T_1296[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2332 = _T_2295 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2347 = _T_2346 | _T_2332; // @[Mux.scala 27:72]
  wire  _T_2298 = _T_2279 == 4'h6; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1298; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_6 = _T_1298[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2333 = _T_2298 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2348 = _T_2347 | _T_2333; // @[Mux.scala 27:72]
  wire  _T_2301 = _T_2279 == 4'h7; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1300; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_7 = _T_1300[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2334 = _T_2301 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2349 = _T_2348 | _T_2334; // @[Mux.scala 27:72]
  wire  _T_2304 = _T_2279 == 4'h8; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1302; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_8 = _T_1302[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2335 = _T_2304 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2350 = _T_2349 | _T_2335; // @[Mux.scala 27:72]
  wire  _T_2307 = _T_2279 == 4'h9; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1304; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_9 = _T_1304[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2336 = _T_2307 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2351 = _T_2350 | _T_2336; // @[Mux.scala 27:72]
  wire  _T_2310 = _T_2279 == 4'ha; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1306; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_10 = _T_1306[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2337 = _T_2310 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2352 = _T_2351 | _T_2337; // @[Mux.scala 27:72]
  wire  _T_2313 = _T_2279 == 4'hb; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1308; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_11 = _T_1308[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2338 = _T_2313 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2353 = _T_2352 | _T_2338; // @[Mux.scala 27:72]
  wire  _T_2316 = _T_2279 == 4'hc; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1310; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_12 = _T_1310[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2339 = _T_2316 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2354 = _T_2353 | _T_2339; // @[Mux.scala 27:72]
  wire  _T_2319 = _T_2279 == 4'hd; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1312; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_13 = _T_1312[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2340 = _T_2319 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2355 = _T_2354 | _T_2340; // @[Mux.scala 27:72]
  wire  _T_2322 = _T_2279 == 4'he; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1314; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_14 = _T_1314[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 390:26]
  wire [31:0] _T_2341 = _T_2322 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2356 = _T_2355 | _T_2341; // @[Mux.scala 27:72]
  wire  _T_2325 = _T_2279 == 4'hf; // @[el2_ifu_mem_ctl.scala 455:89]
  reg [63:0] _T_1316; // @[Reg.scala 27:20]
  wire [31:0] ic_miss_buff_data_15 = _T_1316[31:0]; // @[el2_ifu_mem_ctl.scala 388:31 el2_ifu_mem_ctl.scala 391:28]
  wire [31:0] _T_2342 = _T_2325 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2357 = _T_2356 | _T_2342; // @[Mux.scala 27:72]
  wire [3:0] _T_2359 = {ifu_bus_rid_ff[2:1],_T_2238,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2360 = _T_2359 == 4'h0; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2383 = _T_2360 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2363 = _T_2359 == 4'h1; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2384 = _T_2363 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2391 = _T_2383 | _T_2384; // @[Mux.scala 27:72]
  wire  _T_2366 = _T_2359 == 4'h2; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2385 = _T_2366 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2392 = _T_2391 | _T_2385; // @[Mux.scala 27:72]
  wire  _T_2369 = _T_2359 == 4'h3; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2386 = _T_2369 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2393 = _T_2392 | _T_2386; // @[Mux.scala 27:72]
  wire  _T_2372 = _T_2359 == 4'h4; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2387 = _T_2372 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2394 = _T_2393 | _T_2387; // @[Mux.scala 27:72]
  wire  _T_2375 = _T_2359 == 4'h5; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2388 = _T_2375 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2395 = _T_2394 | _T_2388; // @[Mux.scala 27:72]
  wire  _T_2378 = _T_2359 == 4'h6; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2389 = _T_2378 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2396 = _T_2395 | _T_2389; // @[Mux.scala 27:72]
  wire  _T_2381 = _T_2359 == 4'h7; // @[el2_ifu_mem_ctl.scala 456:64]
  wire [31:0] _T_2390 = _T_2381 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2397 = _T_2396 | _T_2390; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2357,_T_2397}; // @[Cat.scala 29:58]
  wire [7:0] _T_983 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:27]
  wire [16:0] _T_992 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_983}; // @[el2_lib.scala 348:27]
  wire [8:0] _T_1000 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 348:27]
  wire [17:0] _T_1009 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1000}; // @[el2_lib.scala 348:27]
  wire [34:0] _T_1010 = {_T_1009,_T_992}; // @[el2_lib.scala 348:27]
  wire  _T_1011 = ^_T_1010; // @[el2_lib.scala 348:34]
  wire [7:0] _T_1018 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 348:44]
  wire [16:0] _T_1027 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1018}; // @[el2_lib.scala 348:44]
  wire [8:0] _T_1035 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:44]
  wire [17:0] _T_1044 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1035}; // @[el2_lib.scala 348:44]
  wire [34:0] _T_1045 = {_T_1044,_T_1027}; // @[el2_lib.scala 348:44]
  wire  _T_1046 = ^_T_1045; // @[el2_lib.scala 348:51]
  wire [7:0] _T_1053 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 348:61]
  wire [16:0] _T_1062 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1053}; // @[el2_lib.scala 348:61]
  wire [8:0] _T_1070 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 348:61]
  wire [17:0] _T_1079 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1070}; // @[el2_lib.scala 348:61]
  wire [34:0] _T_1080 = {_T_1079,_T_1062}; // @[el2_lib.scala 348:61]
  wire  _T_1081 = ^_T_1080; // @[el2_lib.scala 348:68]
  wire [6:0] _T_1087 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 348:78]
  wire [14:0] _T_1095 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1087}; // @[el2_lib.scala 348:78]
  wire [7:0] _T_1102 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 348:78]
  wire [30:0] _T_1111 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1102,_T_1095}; // @[el2_lib.scala 348:78]
  wire  _T_1112 = ^_T_1111; // @[el2_lib.scala 348:85]
  wire [6:0] _T_1118 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 348:95]
  wire [14:0] _T_1126 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1118}; // @[el2_lib.scala 348:95]
  wire [7:0] _T_1133 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 348:95]
  wire [30:0] _T_1142 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1133,_T_1126}; // @[el2_lib.scala 348:95]
  wire  _T_1143 = ^_T_1142; // @[el2_lib.scala 348:102]
  wire [6:0] _T_1149 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 348:112]
  wire [14:0] _T_1157 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_1149}; // @[el2_lib.scala 348:112]
  wire [30:0] _T_1173 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1133,_T_1157}; // @[el2_lib.scala 348:112]
  wire  _T_1174 = ^_T_1173; // @[el2_lib.scala 348:119]
  wire [6:0] _T_1180 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 348:129]
  wire  _T_1181 = ^_T_1180; // @[el2_lib.scala 348:136]
  wire [70:0] _T_1228 = {_T_589,_T_624,_T_659,_T_690,_T_721,_T_752,_T_759,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1227 = {_T_1011,_T_1046,_T_1081,_T_1112,_T_1143,_T_1174,_T_1181,_T_2357,_T_2397}; // @[Cat.scala 29:58]
  wire [141:0] _T_1229 = {_T_589,_T_624,_T_659,_T_690,_T_721,_T_752,_T_759,ifu_bus_rdata_ff,_T_1227}; // @[Cat.scala 29:58]
  wire [141:0] _T_1232 = {_T_1011,_T_1046,_T_1081,_T_1112,_T_1143,_T_1174,_T_1181,_T_2357,_T_2397,_T_1228}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1229 : _T_1232; // @[el2_ifu_mem_ctl.scala 348:28]
  wire  _T_1189 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 338:56]
  wire  _T_1190 = _T_1189 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 338:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 402:28]
  wire  _T_1392 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 602:35]
  wire  _T_1277 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1277; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1318 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 393:118]
  wire  _T_1319 = ic_miss_buff_data_valid[0] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1319; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1415 = _T_1392 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1395 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1278 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1278; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1322 = ic_miss_buff_data_valid[1] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1322; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1416 = _T_1395 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1423 = _T_1415 | _T_1416; // @[Mux.scala 27:72]
  wire  _T_1398 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1279 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1279; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1325 = ic_miss_buff_data_valid[2] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1325; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1417 = _T_1398 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1424 = _T_1423 | _T_1417; // @[Mux.scala 27:72]
  wire  _T_1401 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1280 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1280; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1328 = ic_miss_buff_data_valid[3] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1328; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1418 = _T_1401 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1425 = _T_1424 | _T_1418; // @[Mux.scala 27:72]
  wire  _T_1404 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1281 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1281; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1331 = ic_miss_buff_data_valid[4] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1331; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1419 = _T_1404 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1426 = _T_1425 | _T_1419; // @[Mux.scala 27:72]
  wire  _T_1407 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1282 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1334 = ic_miss_buff_data_valid[5] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1334; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1420 = _T_1407 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1427 = _T_1426 | _T_1420; // @[Mux.scala 27:72]
  wire  _T_1410 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1337 = ic_miss_buff_data_valid[6] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1337; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1421 = _T_1410 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1428 = _T_1427 | _T_1421; // @[Mux.scala 27:72]
  wire  _T_1413 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 404:114]
  wire  _T_1284 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 387:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 387:73]
  wire  _T_1340 = ic_miss_buff_data_valid[7] & _T_1318; // @[el2_ifu_mem_ctl.scala 393:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1340; // @[el2_ifu_mem_ctl.scala 393:88]
  wire  _T_1422 = _T_1413 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1428 | _T_1422; // @[Mux.scala 27:72]
  wire  _T_1431 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 405:58]
  wire  _T_1432 = bypass_valid_value_check & _T_1431; // @[el2_ifu_mem_ctl.scala 405:56]
  wire  _T_1434 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 405:77]
  wire  _T_1435 = _T_1432 & _T_1434; // @[el2_ifu_mem_ctl.scala 405:75]
  wire  _T_1440 = _T_1432 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 406:75]
  wire  _T_1441 = _T_1435 | _T_1440; // @[el2_ifu_mem_ctl.scala 405:95]
  wire  _T_1443 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 407:56]
  wire  _T_1446 = _T_1443 & _T_1434; // @[el2_ifu_mem_ctl.scala 407:74]
  wire  _T_1447 = _T_1441 | _T_1446; // @[el2_ifu_mem_ctl.scala 406:94]
  wire  _T_1451 = _T_1443 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 408:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 403:70]
  wire  _T_1452 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1468 = _T_1452 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1454 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1469 = _T_1454 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1476 = _T_1468 | _T_1469; // @[Mux.scala 27:72]
  wire  _T_1456 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1470 = _T_1456 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1477 = _T_1476 | _T_1470; // @[Mux.scala 27:72]
  wire  _T_1458 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1471 = _T_1458 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1478 = _T_1477 | _T_1471; // @[Mux.scala 27:72]
  wire  _T_1460 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1472 = _T_1460 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1479 = _T_1478 | _T_1472; // @[Mux.scala 27:72]
  wire  _T_1462 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1473 = _T_1462 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1480 = _T_1479 | _T_1473; // @[Mux.scala 27:72]
  wire  _T_1464 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1474 = _T_1464 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1481 = _T_1480 | _T_1474; // @[Mux.scala 27:72]
  wire  _T_1466 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 408:132]
  wire  _T_1475 = _T_1466 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1482 = _T_1481 | _T_1475; // @[Mux.scala 27:72]
  wire  _T_1484 = _T_1451 & _T_1482; // @[el2_ifu_mem_ctl.scala 408:69]
  wire  _T_1485 = _T_1447 | _T_1484; // @[el2_ifu_mem_ctl.scala 407:94]
  wire [4:0] _GEN_664 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 409:95]
  wire  _T_1488 = _GEN_664 == 5'h1f; // @[el2_ifu_mem_ctl.scala 409:95]
  wire  _T_1489 = bypass_valid_value_check & _T_1488; // @[el2_ifu_mem_ctl.scala 409:56]
  wire  bypass_data_ready_in = _T_1485 | _T_1489; // @[el2_ifu_mem_ctl.scala 408:181]
  wire  _T_1490 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 413:53]
  wire  _T_1491 = _T_1490 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 413:73]
  wire  _T_1493 = _T_1491 & _T_308; // @[el2_ifu_mem_ctl.scala 413:96]
  wire  _T_1495 = _T_1493 & _T_60; // @[el2_ifu_mem_ctl.scala 413:118]
  wire  _T_1497 = crit_wd_byp_ok_ff & _T_51; // @[el2_ifu_mem_ctl.scala 414:73]
  wire  _T_1499 = _T_1497 & _T_308; // @[el2_ifu_mem_ctl.scala 414:96]
  wire  _T_1501 = _T_1499 & _T_60; // @[el2_ifu_mem_ctl.scala 414:118]
  wire  _T_1502 = _T_1495 | _T_1501; // @[el2_ifu_mem_ctl.scala 413:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 416:58]
  wire  _T_1503 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 415:54]
  wire  _T_1504 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 415:76]
  wire  _T_1505 = _T_1503 & _T_1504; // @[el2_ifu_mem_ctl.scala 415:74]
  wire  _T_1507 = _T_1505 & _T_308; // @[el2_ifu_mem_ctl.scala 415:96]
  wire  ic_crit_wd_rdy_new_in = _T_1502 | _T_1507; // @[el2_ifu_mem_ctl.scala 414:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 612:43]
  wire  _T_1244 = ic_crit_wd_rdy | _T_2218; // @[el2_ifu_mem_ctl.scala 360:38]
  wire  _T_1246 = _T_1244 | _T_2233; // @[el2_ifu_mem_ctl.scala 360:64]
  wire  _T_1247 = ~_T_1246; // @[el2_ifu_mem_ctl.scala 360:21]
  wire  _T_1248 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 360:98]
  wire  sel_ic_data = _T_1247 & _T_1248; // @[el2_ifu_mem_ctl.scala 360:96]
  wire  _T_2400 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 458:44]
  wire  _T_1601 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 427:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 399:60]
  wire  _T_1545 = _T_1392 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1546 = _T_1395 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1553 = _T_1545 | _T_1546; // @[Mux.scala 27:72]
  wire  _T_1547 = _T_1398 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1554 = _T_1553 | _T_1547; // @[Mux.scala 27:72]
  wire  _T_1548 = _T_1401 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1555 = _T_1554 | _T_1548; // @[Mux.scala 27:72]
  wire  _T_1549 = _T_1404 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1556 = _T_1555 | _T_1549; // @[Mux.scala 27:72]
  wire  _T_1550 = _T_1407 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1556 | _T_1550; // @[Mux.scala 27:72]
  wire  _T_1551 = _T_1410 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1558 = _T_1557 | _T_1551; // @[Mux.scala 27:72]
  wire  _T_1552 = _T_1413 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1558 | _T_1552; // @[Mux.scala 27:72]
  wire  _T_1584 = _T_2145 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1585 = _T_2148 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1592 = _T_1584 | _T_1585; // @[Mux.scala 27:72]
  wire  _T_1586 = _T_2151 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1593 = _T_1592 | _T_1586; // @[Mux.scala 27:72]
  wire  _T_1587 = _T_2154 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1594 = _T_1593 | _T_1587; // @[Mux.scala 27:72]
  wire  _T_1588 = _T_2157 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1595 = _T_1594 | _T_1588; // @[Mux.scala 27:72]
  wire  _T_1589 = _T_2160 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1596 = _T_1595 | _T_1589; // @[Mux.scala 27:72]
  wire  _T_1590 = _T_2163 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1597 = _T_1596 | _T_1590; // @[Mux.scala 27:72]
  wire  _T_1591 = _T_2166 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1597 | _T_1591; // @[Mux.scala 27:72]
  wire  _T_1602 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 429:70]
  wire  ifu_byp_data_err_new = _T_1601 ? ic_miss_buff_data_error_bypass : _T_1602; // @[el2_ifu_mem_ctl.scala 427:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 371:42]
  wire  _T_2401 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 458:91]
  wire  _T_2402 = ~_T_2401; // @[el2_ifu_mem_ctl.scala 458:60]
  wire  ic_rd_parity_final_err = _T_2400 & _T_2402; // @[el2_ifu_mem_ctl.scala 458:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_9671 = _T_4465 ? 1'h0 : ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 739:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_9673 = _T_4469 ? 1'h0 : ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9926 = _T_9671 | _T_9673; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_9675 = _T_4473 ? 1'h0 : ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9927 = _T_9926 | _T_9675; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_9677 = _T_4477 ? 1'h0 : ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9928 = _T_9927 | _T_9677; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_9679 = _T_4481 ? 1'h0 : ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9929 = _T_9928 | _T_9679; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_9681 = _T_4485 ? 1'h0 : ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9930 = _T_9929 | _T_9681; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_9683 = _T_4489 ? 1'h0 : ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9931 = _T_9930 | _T_9683; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_9685 = _T_4493 ? 1'h0 : ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9932 = _T_9931 | _T_9685; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_9687 = _T_4497 ? 1'h0 : ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9933 = _T_9932 | _T_9687; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_9689 = _T_4501 ? 1'h0 : ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9934 = _T_9933 | _T_9689; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_9691 = _T_4505 ? 1'h0 : ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9935 = _T_9934 | _T_9691; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_9693 = _T_4509 ? 1'h0 : ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9936 = _T_9935 | _T_9693; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_9695 = _T_4513 ? 1'h0 : ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9937 = _T_9936 | _T_9695; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_9697 = _T_4517 ? 1'h0 : ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9938 = _T_9937 | _T_9697; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_9699 = _T_4521 ? 1'h0 : ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9939 = _T_9938 | _T_9699; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_9701 = _T_4525 ? 1'h0 : ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9940 = _T_9939 | _T_9701; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_9703 = _T_4529 ? 1'h0 : ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9941 = _T_9940 | _T_9703; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_9705 = _T_4533 ? 1'h0 : ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9942 = _T_9941 | _T_9705; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_9707 = _T_4537 ? 1'h0 : ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9943 = _T_9942 | _T_9707; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_9709 = _T_4541 ? 1'h0 : ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9944 = _T_9943 | _T_9709; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_9711 = _T_4545 ? 1'h0 : ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9945 = _T_9944 | _T_9711; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_9713 = _T_4549 ? 1'h0 : ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9946 = _T_9945 | _T_9713; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_9715 = _T_4553 ? 1'h0 : ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9947 = _T_9946 | _T_9715; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_9717 = _T_4557 ? 1'h0 : ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9948 = _T_9947 | _T_9717; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_9719 = _T_4561 ? 1'h0 : ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9949 = _T_9948 | _T_9719; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_9721 = _T_4565 ? 1'h0 : ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9950 = _T_9949 | _T_9721; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_9723 = _T_4569 ? 1'h0 : ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9951 = _T_9950 | _T_9723; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_9725 = _T_4573 ? 1'h0 : ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9952 = _T_9951 | _T_9725; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_9727 = _T_4577 ? 1'h0 : ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9953 = _T_9952 | _T_9727; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_9729 = _T_4581 ? 1'h0 : ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9954 = _T_9953 | _T_9729; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_9731 = _T_4585 ? 1'h0 : ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9955 = _T_9954 | _T_9731; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_9733 = _T_4589 ? 1'h0 : ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9956 = _T_9955 | _T_9733; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_9735 = _T_4593 ? 1'h0 : ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9957 = _T_9956 | _T_9735; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_9737 = _T_4597 ? 1'h0 : ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9958 = _T_9957 | _T_9737; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_9739 = _T_4601 ? 1'h0 : ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9959 = _T_9958 | _T_9739; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_9741 = _T_4605 ? 1'h0 : ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9960 = _T_9959 | _T_9741; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_9743 = _T_4609 ? 1'h0 : ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9961 = _T_9960 | _T_9743; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_9745 = _T_4613 ? 1'h0 : ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9962 = _T_9961 | _T_9745; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_9747 = _T_4617 ? 1'h0 : ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9963 = _T_9962 | _T_9747; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_9749 = _T_4621 ? 1'h0 : ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9964 = _T_9963 | _T_9749; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_9751 = _T_4625 ? 1'h0 : ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9965 = _T_9964 | _T_9751; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_9753 = _T_4629 ? 1'h0 : ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9966 = _T_9965 | _T_9753; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_9755 = _T_4633 ? 1'h0 : ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9967 = _T_9966 | _T_9755; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_9757 = _T_4637 ? 1'h0 : ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9968 = _T_9967 | _T_9757; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_9759 = _T_4641 ? 1'h0 : ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9969 = _T_9968 | _T_9759; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_9761 = _T_4645 ? 1'h0 : ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9970 = _T_9969 | _T_9761; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_9763 = _T_4649 ? 1'h0 : ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9971 = _T_9970 | _T_9763; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_9765 = _T_4653 ? 1'h0 : ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9972 = _T_9971 | _T_9765; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_9767 = _T_4657 ? 1'h0 : ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9973 = _T_9972 | _T_9767; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_9769 = _T_4661 ? 1'h0 : ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9974 = _T_9973 | _T_9769; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_9771 = _T_4665 ? 1'h0 : ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9975 = _T_9974 | _T_9771; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_9773 = _T_4669 ? 1'h0 : ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9976 = _T_9975 | _T_9773; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_9775 = _T_4673 ? 1'h0 : ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9977 = _T_9976 | _T_9775; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_9777 = _T_4677 ? 1'h0 : ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9978 = _T_9977 | _T_9777; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_9779 = _T_4681 ? 1'h0 : ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9979 = _T_9978 | _T_9779; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_9781 = _T_4685 ? 1'h0 : ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9980 = _T_9979 | _T_9781; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_9783 = _T_4689 ? 1'h0 : ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9981 = _T_9980 | _T_9783; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9785 = _T_4693 ? 1'h0 : ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9982 = _T_9981 | _T_9785; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9787 = _T_4697 ? 1'h0 : ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9983 = _T_9982 | _T_9787; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9789 = _T_4701 ? 1'h0 : ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9984 = _T_9983 | _T_9789; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9791 = _T_4705 ? 1'h0 : ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9985 = _T_9984 | _T_9791; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9793 = _T_4709 ? 1'h0 : ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9986 = _T_9985 | _T_9793; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9795 = _T_4713 ? 1'h0 : ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9987 = _T_9986 | _T_9795; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9797 = _T_4717 ? 1'h0 : ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9988 = _T_9987 | _T_9797; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9799 = _T_4721 ? 1'h0 : ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9989 = _T_9988 | _T_9799; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9801 = _T_4725 ? 1'h0 : ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9990 = _T_9989 | _T_9801; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9803 = _T_4729 ? 1'h0 : ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9991 = _T_9990 | _T_9803; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9805 = _T_4733 ? 1'h0 : ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9992 = _T_9991 | _T_9805; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9807 = _T_4737 ? 1'h0 : ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9993 = _T_9992 | _T_9807; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9809 = _T_4741 ? 1'h0 : ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9994 = _T_9993 | _T_9809; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9811 = _T_4745 ? 1'h0 : ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9995 = _T_9994 | _T_9811; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9813 = _T_4749 ? 1'h0 : ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9996 = _T_9995 | _T_9813; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9815 = _T_4753 ? 1'h0 : ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9997 = _T_9996 | _T_9815; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9817 = _T_4757 ? 1'h0 : ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9998 = _T_9997 | _T_9817; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9819 = _T_4761 ? 1'h0 : ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9999 = _T_9998 | _T_9819; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9821 = _T_4765 ? 1'h0 : ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10000 = _T_9999 | _T_9821; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9823 = _T_4769 ? 1'h0 : ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10001 = _T_10000 | _T_9823; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9825 = _T_4773 ? 1'h0 : ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10002 = _T_10001 | _T_9825; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9827 = _T_4777 ? 1'h0 : ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10003 = _T_10002 | _T_9827; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9829 = _T_4781 ? 1'h0 : ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10004 = _T_10003 | _T_9829; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9831 = _T_4785 ? 1'h0 : ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10005 = _T_10004 | _T_9831; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9833 = _T_4789 ? 1'h0 : ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10006 = _T_10005 | _T_9833; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9835 = _T_4793 ? 1'h0 : ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10007 = _T_10006 | _T_9835; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9837 = _T_4797 ? 1'h0 : ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10008 = _T_10007 | _T_9837; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9839 = _T_4801 ? 1'h0 : ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10009 = _T_10008 | _T_9839; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9841 = _T_4805 ? 1'h0 : ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10010 = _T_10009 | _T_9841; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9843 = _T_4809 ? 1'h0 : ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10011 = _T_10010 | _T_9843; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9845 = _T_4813 ? 1'h0 : ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10012 = _T_10011 | _T_9845; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9847 = _T_4817 ? 1'h0 : ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10013 = _T_10012 | _T_9847; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9849 = _T_4821 ? 1'h0 : ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10014 = _T_10013 | _T_9849; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9851 = _T_4825 ? 1'h0 : ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10015 = _T_10014 | _T_9851; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9853 = _T_4829 ? 1'h0 : ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10016 = _T_10015 | _T_9853; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9855 = _T_4833 ? 1'h0 : ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10017 = _T_10016 | _T_9855; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9857 = _T_4837 ? 1'h0 : ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10018 = _T_10017 | _T_9857; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9859 = _T_4841 ? 1'h0 : ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10019 = _T_10018 | _T_9859; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9861 = _T_4845 ? 1'h0 : ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10020 = _T_10019 | _T_9861; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9863 = _T_4849 ? 1'h0 : ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10021 = _T_10020 | _T_9863; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9865 = _T_4853 ? 1'h0 : ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10022 = _T_10021 | _T_9865; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9867 = _T_4857 ? 1'h0 : ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10023 = _T_10022 | _T_9867; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9869 = _T_4861 ? 1'h0 : ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10024 = _T_10023 | _T_9869; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9871 = _T_4865 ? 1'h0 : ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10025 = _T_10024 | _T_9871; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9873 = _T_4869 ? 1'h0 : ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10026 = _T_10025 | _T_9873; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9875 = _T_4873 ? 1'h0 : ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10027 = _T_10026 | _T_9875; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9877 = _T_4877 ? 1'h0 : ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10028 = _T_10027 | _T_9877; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9879 = _T_4881 ? 1'h0 : ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10029 = _T_10028 | _T_9879; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9881 = _T_4885 ? 1'h0 : ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10030 = _T_10029 | _T_9881; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9883 = _T_4889 ? 1'h0 : ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10031 = _T_10030 | _T_9883; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9885 = _T_4893 ? 1'h0 : ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10032 = _T_10031 | _T_9885; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9887 = _T_4897 ? 1'h0 : ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10033 = _T_10032 | _T_9887; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9889 = _T_4901 ? 1'h0 : ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10034 = _T_10033 | _T_9889; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9891 = _T_4905 ? 1'h0 : ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10035 = _T_10034 | _T_9891; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9893 = _T_4909 ? 1'h0 : ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10036 = _T_10035 | _T_9893; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9895 = _T_4913 ? 1'h0 : ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10037 = _T_10036 | _T_9895; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9897 = _T_4917 ? 1'h0 : ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10038 = _T_10037 | _T_9897; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9899 = _T_4921 ? 1'h0 : ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10039 = _T_10038 | _T_9899; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9901 = _T_4925 ? 1'h0 : ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10040 = _T_10039 | _T_9901; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9903 = _T_4929 ? 1'h0 : ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10041 = _T_10040 | _T_9903; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9905 = _T_4933 ? 1'h0 : ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10042 = _T_10041 | _T_9905; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9907 = _T_4937 ? 1'h0 : ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10043 = _T_10042 | _T_9907; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9909 = _T_4941 ? 1'h0 : ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10044 = _T_10043 | _T_9909; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9911 = _T_4945 ? 1'h0 : ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10045 = _T_10044 | _T_9911; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9913 = _T_4949 ? 1'h0 : ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10046 = _T_10045 | _T_9913; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9915 = _T_4953 ? 1'h0 : ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10047 = _T_10046 | _T_9915; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9917 = _T_4957 ? 1'h0 : ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10048 = _T_10047 | _T_9917; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9919 = _T_4961 ? 1'h0 : ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10049 = _T_10048 | _T_9919; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9921 = _T_4965 ? 1'h0 : ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10050 = _T_10049 | _T_9921; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9923 = _T_4969 ? 1'h0 : ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10051 = _T_10050 | _T_9923; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9925 = _T_4973 ? 1'h0 : ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_10052 = _T_10051 | _T_9925; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9288 = _T_4465 ? 1'h0 : ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 739:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9290 = _T_4469 ? 1'h0 : ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9543 = _T_9288 | _T_9290; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9292 = _T_4473 ? 1'h0 : ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9544 = _T_9543 | _T_9292; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9294 = _T_4477 ? 1'h0 : ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9545 = _T_9544 | _T_9294; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9296 = _T_4481 ? 1'h0 : ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9546 = _T_9545 | _T_9296; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9298 = _T_4485 ? 1'h0 : ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9547 = _T_9546 | _T_9298; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9300 = _T_4489 ? 1'h0 : ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9548 = _T_9547 | _T_9300; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9302 = _T_4493 ? 1'h0 : ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9549 = _T_9548 | _T_9302; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9304 = _T_4497 ? 1'h0 : ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9550 = _T_9549 | _T_9304; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9306 = _T_4501 ? 1'h0 : ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9551 = _T_9550 | _T_9306; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9308 = _T_4505 ? 1'h0 : ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9552 = _T_9551 | _T_9308; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9310 = _T_4509 ? 1'h0 : ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9553 = _T_9552 | _T_9310; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9312 = _T_4513 ? 1'h0 : ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9554 = _T_9553 | _T_9312; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9314 = _T_4517 ? 1'h0 : ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9555 = _T_9554 | _T_9314; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9316 = _T_4521 ? 1'h0 : ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9556 = _T_9555 | _T_9316; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9318 = _T_4525 ? 1'h0 : ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9557 = _T_9556 | _T_9318; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9320 = _T_4529 ? 1'h0 : ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9558 = _T_9557 | _T_9320; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9322 = _T_4533 ? 1'h0 : ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9559 = _T_9558 | _T_9322; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9324 = _T_4537 ? 1'h0 : ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9560 = _T_9559 | _T_9324; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9326 = _T_4541 ? 1'h0 : ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9561 = _T_9560 | _T_9326; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9328 = _T_4545 ? 1'h0 : ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9562 = _T_9561 | _T_9328; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9330 = _T_4549 ? 1'h0 : ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9563 = _T_9562 | _T_9330; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9332 = _T_4553 ? 1'h0 : ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9564 = _T_9563 | _T_9332; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9334 = _T_4557 ? 1'h0 : ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9565 = _T_9564 | _T_9334; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9336 = _T_4561 ? 1'h0 : ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9566 = _T_9565 | _T_9336; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9338 = _T_4565 ? 1'h0 : ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9567 = _T_9566 | _T_9338; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9340 = _T_4569 ? 1'h0 : ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9568 = _T_9567 | _T_9340; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9342 = _T_4573 ? 1'h0 : ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9569 = _T_9568 | _T_9342; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9344 = _T_4577 ? 1'h0 : ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9570 = _T_9569 | _T_9344; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9346 = _T_4581 ? 1'h0 : ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9571 = _T_9570 | _T_9346; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9348 = _T_4585 ? 1'h0 : ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9572 = _T_9571 | _T_9348; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9350 = _T_4589 ? 1'h0 : ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9573 = _T_9572 | _T_9350; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9352 = _T_4593 ? 1'h0 : ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9574 = _T_9573 | _T_9352; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9354 = _T_4597 ? 1'h0 : ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9575 = _T_9574 | _T_9354; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9356 = _T_4601 ? 1'h0 : ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9576 = _T_9575 | _T_9356; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9358 = _T_4605 ? 1'h0 : ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9577 = _T_9576 | _T_9358; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9360 = _T_4609 ? 1'h0 : ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9578 = _T_9577 | _T_9360; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9362 = _T_4613 ? 1'h0 : ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9579 = _T_9578 | _T_9362; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9364 = _T_4617 ? 1'h0 : ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9580 = _T_9579 | _T_9364; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9366 = _T_4621 ? 1'h0 : ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9581 = _T_9580 | _T_9366; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9368 = _T_4625 ? 1'h0 : ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9582 = _T_9581 | _T_9368; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9370 = _T_4629 ? 1'h0 : ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9583 = _T_9582 | _T_9370; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9372 = _T_4633 ? 1'h0 : ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9584 = _T_9583 | _T_9372; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9374 = _T_4637 ? 1'h0 : ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9585 = _T_9584 | _T_9374; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9376 = _T_4641 ? 1'h0 : ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9586 = _T_9585 | _T_9376; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9378 = _T_4645 ? 1'h0 : ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9587 = _T_9586 | _T_9378; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9380 = _T_4649 ? 1'h0 : ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9588 = _T_9587 | _T_9380; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9382 = _T_4653 ? 1'h0 : ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9589 = _T_9588 | _T_9382; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9384 = _T_4657 ? 1'h0 : ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9590 = _T_9589 | _T_9384; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9386 = _T_4661 ? 1'h0 : ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9591 = _T_9590 | _T_9386; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9388 = _T_4665 ? 1'h0 : ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9592 = _T_9591 | _T_9388; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9390 = _T_4669 ? 1'h0 : ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9593 = _T_9592 | _T_9390; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9392 = _T_4673 ? 1'h0 : ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9594 = _T_9593 | _T_9392; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9394 = _T_4677 ? 1'h0 : ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9595 = _T_9594 | _T_9394; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9396 = _T_4681 ? 1'h0 : ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9596 = _T_9595 | _T_9396; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9398 = _T_4685 ? 1'h0 : ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9597 = _T_9596 | _T_9398; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9400 = _T_4689 ? 1'h0 : ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9598 = _T_9597 | _T_9400; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9402 = _T_4693 ? 1'h0 : ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9599 = _T_9598 | _T_9402; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9404 = _T_4697 ? 1'h0 : ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9600 = _T_9599 | _T_9404; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9406 = _T_4701 ? 1'h0 : ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9601 = _T_9600 | _T_9406; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9408 = _T_4705 ? 1'h0 : ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9602 = _T_9601 | _T_9408; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9410 = _T_4709 ? 1'h0 : ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9603 = _T_9602 | _T_9410; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9412 = _T_4713 ? 1'h0 : ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9604 = _T_9603 | _T_9412; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9414 = _T_4717 ? 1'h0 : ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9605 = _T_9604 | _T_9414; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9416 = _T_4721 ? 1'h0 : ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9606 = _T_9605 | _T_9416; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9418 = _T_4725 ? 1'h0 : ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9607 = _T_9606 | _T_9418; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9420 = _T_4729 ? 1'h0 : ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9608 = _T_9607 | _T_9420; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9422 = _T_4733 ? 1'h0 : ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9609 = _T_9608 | _T_9422; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9424 = _T_4737 ? 1'h0 : ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9610 = _T_9609 | _T_9424; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9426 = _T_4741 ? 1'h0 : ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9611 = _T_9610 | _T_9426; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9428 = _T_4745 ? 1'h0 : ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9612 = _T_9611 | _T_9428; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9430 = _T_4749 ? 1'h0 : ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9613 = _T_9612 | _T_9430; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9432 = _T_4753 ? 1'h0 : ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9614 = _T_9613 | _T_9432; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9434 = _T_4757 ? 1'h0 : ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9615 = _T_9614 | _T_9434; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9436 = _T_4761 ? 1'h0 : ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9616 = _T_9615 | _T_9436; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9438 = _T_4765 ? 1'h0 : ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9617 = _T_9616 | _T_9438; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9440 = _T_4769 ? 1'h0 : ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9618 = _T_9617 | _T_9440; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9442 = _T_4773 ? 1'h0 : ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9619 = _T_9618 | _T_9442; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9444 = _T_4777 ? 1'h0 : ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9620 = _T_9619 | _T_9444; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9446 = _T_4781 ? 1'h0 : ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9621 = _T_9620 | _T_9446; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9448 = _T_4785 ? 1'h0 : ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9622 = _T_9621 | _T_9448; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9450 = _T_4789 ? 1'h0 : ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9623 = _T_9622 | _T_9450; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9452 = _T_4793 ? 1'h0 : ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9624 = _T_9623 | _T_9452; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9454 = _T_4797 ? 1'h0 : ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9625 = _T_9624 | _T_9454; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9456 = _T_4801 ? 1'h0 : ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9626 = _T_9625 | _T_9456; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9458 = _T_4805 ? 1'h0 : ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9627 = _T_9626 | _T_9458; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9460 = _T_4809 ? 1'h0 : ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9628 = _T_9627 | _T_9460; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9462 = _T_4813 ? 1'h0 : ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9629 = _T_9628 | _T_9462; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9464 = _T_4817 ? 1'h0 : ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9630 = _T_9629 | _T_9464; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9466 = _T_4821 ? 1'h0 : ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9631 = _T_9630 | _T_9466; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9468 = _T_4825 ? 1'h0 : ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9632 = _T_9631 | _T_9468; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9470 = _T_4829 ? 1'h0 : ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9633 = _T_9632 | _T_9470; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9472 = _T_4833 ? 1'h0 : ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9634 = _T_9633 | _T_9472; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9474 = _T_4837 ? 1'h0 : ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9635 = _T_9634 | _T_9474; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9476 = _T_4841 ? 1'h0 : ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9636 = _T_9635 | _T_9476; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9478 = _T_4845 ? 1'h0 : ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9637 = _T_9636 | _T_9478; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9480 = _T_4849 ? 1'h0 : ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9638 = _T_9637 | _T_9480; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9482 = _T_4853 ? 1'h0 : ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9639 = _T_9638 | _T_9482; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9484 = _T_4857 ? 1'h0 : ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9640 = _T_9639 | _T_9484; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9486 = _T_4861 ? 1'h0 : ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9641 = _T_9640 | _T_9486; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9488 = _T_4865 ? 1'h0 : ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9642 = _T_9641 | _T_9488; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9490 = _T_4869 ? 1'h0 : ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9643 = _T_9642 | _T_9490; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9492 = _T_4873 ? 1'h0 : ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9644 = _T_9643 | _T_9492; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9494 = _T_4877 ? 1'h0 : ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9645 = _T_9644 | _T_9494; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9496 = _T_4881 ? 1'h0 : ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9646 = _T_9645 | _T_9496; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9498 = _T_4885 ? 1'h0 : ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9647 = _T_9646 | _T_9498; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9500 = _T_4889 ? 1'h0 : ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9648 = _T_9647 | _T_9500; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9502 = _T_4893 ? 1'h0 : ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9649 = _T_9648 | _T_9502; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9504 = _T_4897 ? 1'h0 : ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9650 = _T_9649 | _T_9504; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9506 = _T_4901 ? 1'h0 : ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9651 = _T_9650 | _T_9506; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9508 = _T_4905 ? 1'h0 : ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9652 = _T_9651 | _T_9508; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9510 = _T_4909 ? 1'h0 : ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9653 = _T_9652 | _T_9510; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9512 = _T_4913 ? 1'h0 : ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9654 = _T_9653 | _T_9512; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9514 = _T_4917 ? 1'h0 : ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9655 = _T_9654 | _T_9514; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_9516 = _T_4921 ? 1'h0 : ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9656 = _T_9655 | _T_9516; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_9518 = _T_4925 ? 1'h0 : ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9657 = _T_9656 | _T_9518; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_9520 = _T_4929 ? 1'h0 : ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9658 = _T_9657 | _T_9520; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_9522 = _T_4933 ? 1'h0 : ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9659 = _T_9658 | _T_9522; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_9524 = _T_4937 ? 1'h0 : ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9660 = _T_9659 | _T_9524; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_9526 = _T_4941 ? 1'h0 : ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9661 = _T_9660 | _T_9526; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_9528 = _T_4945 ? 1'h0 : ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9662 = _T_9661 | _T_9528; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_9530 = _T_4949 ? 1'h0 : ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9663 = _T_9662 | _T_9530; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_9532 = _T_4953 ? 1'h0 : ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9664 = _T_9663 | _T_9532; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_9534 = _T_4957 ? 1'h0 : ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9665 = _T_9664 | _T_9534; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_9536 = _T_4961 ? 1'h0 : ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9666 = _T_9665 | _T_9536; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_9538 = _T_4965 ? 1'h0 : ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9667 = _T_9666 | _T_9538; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_9540 = _T_4969 ? 1'h0 : ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9668 = _T_9667 | _T_9540; // @[el2_ifu_mem_ctl.scala 739:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_9542 = _T_4973 ? 1'h0 : ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 739:10]
  wire  _T_9669 = _T_9668 | _T_9542; // @[el2_ifu_mem_ctl.scala 739:91]
  wire [1:0] ic_tag_valid_unq = {_T_10052,_T_9669}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 810:54]
  wire [1:0] _T_10091 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10092 = ic_debug_way_ff & _T_10091; // @[el2_ifu_mem_ctl.scala 793:67]
  wire [1:0] _T_10093 = ic_tag_valid_unq & _T_10092; // @[el2_ifu_mem_ctl.scala 793:48]
  wire  ic_debug_tag_val_rd_out = |_T_10093; // @[el2_ifu_mem_ctl.scala 793:115]
  wire [65:0] _T_1201 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1202; // @[el2_ifu_mem_ctl.scala 344:37]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2533; // @[el2_ifu_mem_ctl.scala 354:80]
  wire  _T_1242 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 359:98]
  wire  sel_byp_data = _T_1246 & _T_1242; // @[el2_ifu_mem_ctl.scala 359:96]
  wire [63:0] _T_1253 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1254 = _T_1253 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 366:64]
  wire [63:0] _T_1256 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2092 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 435:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1606 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1654 = _T_1606 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1609 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1655 = _T_1609 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1670 = _T_1654 | _T_1655; // @[Mux.scala 27:72]
  wire  _T_1612 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1656 = _T_1612 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1671 = _T_1670 | _T_1656; // @[Mux.scala 27:72]
  wire  _T_1615 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1657 = _T_1615 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1672 = _T_1671 | _T_1657; // @[Mux.scala 27:72]
  wire  _T_1618 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1658 = _T_1618 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1673 = _T_1672 | _T_1658; // @[Mux.scala 27:72]
  wire  _T_1621 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1659 = _T_1621 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1674 = _T_1673 | _T_1659; // @[Mux.scala 27:72]
  wire  _T_1624 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1660 = _T_1624 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1675 = _T_1674 | _T_1660; // @[Mux.scala 27:72]
  wire  _T_1627 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1661 = _T_1627 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1676 = _T_1675 | _T_1661; // @[Mux.scala 27:72]
  wire  _T_1630 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1662 = _T_1630 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1677 = _T_1676 | _T_1662; // @[Mux.scala 27:72]
  wire  _T_1633 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1663 = _T_1633 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1678 = _T_1677 | _T_1663; // @[Mux.scala 27:72]
  wire  _T_1636 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1664 = _T_1636 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1679 = _T_1678 | _T_1664; // @[Mux.scala 27:72]
  wire  _T_1639 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1665 = _T_1639 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1680 = _T_1679 | _T_1665; // @[Mux.scala 27:72]
  wire  _T_1642 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1666 = _T_1642 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1681 = _T_1680 | _T_1666; // @[Mux.scala 27:72]
  wire  _T_1645 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1667 = _T_1645 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1682 = _T_1681 | _T_1667; // @[Mux.scala 27:72]
  wire  _T_1648 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1668 = _T_1648 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1683 = _T_1682 | _T_1668; // @[Mux.scala 27:72]
  wire  _T_1651 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 432:73]
  wire [15:0] _T_1669 = _T_1651 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1684 = _T_1683 | _T_1669; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1686 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1734 = _T_1686 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1689 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1735 = _T_1689 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1750 = _T_1734 | _T_1735; // @[Mux.scala 27:72]
  wire  _T_1692 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1736 = _T_1692 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1751 = _T_1750 | _T_1736; // @[Mux.scala 27:72]
  wire  _T_1695 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1737 = _T_1695 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1752 = _T_1751 | _T_1737; // @[Mux.scala 27:72]
  wire  _T_1698 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1738 = _T_1698 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1753 = _T_1752 | _T_1738; // @[Mux.scala 27:72]
  wire  _T_1701 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1739 = _T_1701 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1754 = _T_1753 | _T_1739; // @[Mux.scala 27:72]
  wire  _T_1704 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1740 = _T_1704 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1755 = _T_1754 | _T_1740; // @[Mux.scala 27:72]
  wire  _T_1707 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1741 = _T_1707 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1756 = _T_1755 | _T_1741; // @[Mux.scala 27:72]
  wire  _T_1710 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1742 = _T_1710 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1757 = _T_1756 | _T_1742; // @[Mux.scala 27:72]
  wire  _T_1713 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1743 = _T_1713 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1758 = _T_1757 | _T_1743; // @[Mux.scala 27:72]
  wire  _T_1716 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1744 = _T_1716 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1759 = _T_1758 | _T_1744; // @[Mux.scala 27:72]
  wire  _T_1719 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1745 = _T_1719 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1760 = _T_1759 | _T_1745; // @[Mux.scala 27:72]
  wire  _T_1722 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1746 = _T_1722 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1761 = _T_1760 | _T_1746; // @[Mux.scala 27:72]
  wire  _T_1725 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1747 = _T_1725 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1762 = _T_1761 | _T_1747; // @[Mux.scala 27:72]
  wire  _T_1728 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1748 = _T_1728 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1763 = _T_1762 | _T_1748; // @[Mux.scala 27:72]
  wire  _T_1731 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 432:179]
  wire [31:0] _T_1749 = _T_1731 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1764 = _T_1763 | _T_1749; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1766 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1814 = _T_1766 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1769 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1815 = _T_1769 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1830 = _T_1814 | _T_1815; // @[Mux.scala 27:72]
  wire  _T_1772 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1816 = _T_1772 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1831 = _T_1830 | _T_1816; // @[Mux.scala 27:72]
  wire  _T_1775 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1817 = _T_1775 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1832 = _T_1831 | _T_1817; // @[Mux.scala 27:72]
  wire  _T_1778 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1818 = _T_1778 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1833 = _T_1832 | _T_1818; // @[Mux.scala 27:72]
  wire  _T_1781 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1819 = _T_1781 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1834 = _T_1833 | _T_1819; // @[Mux.scala 27:72]
  wire  _T_1784 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1820 = _T_1784 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1835 = _T_1834 | _T_1820; // @[Mux.scala 27:72]
  wire  _T_1787 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1821 = _T_1787 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1836 = _T_1835 | _T_1821; // @[Mux.scala 27:72]
  wire  _T_1790 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1822 = _T_1790 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1837 = _T_1836 | _T_1822; // @[Mux.scala 27:72]
  wire  _T_1793 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1823 = _T_1793 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1838 = _T_1837 | _T_1823; // @[Mux.scala 27:72]
  wire  _T_1796 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1824 = _T_1796 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1839 = _T_1838 | _T_1824; // @[Mux.scala 27:72]
  wire  _T_1799 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1825 = _T_1799 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1840 = _T_1839 | _T_1825; // @[Mux.scala 27:72]
  wire  _T_1802 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1826 = _T_1802 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1841 = _T_1840 | _T_1826; // @[Mux.scala 27:72]
  wire  _T_1805 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1827 = _T_1805 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1842 = _T_1841 | _T_1827; // @[Mux.scala 27:72]
  wire  _T_1808 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1828 = _T_1808 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1843 = _T_1842 | _T_1828; // @[Mux.scala 27:72]
  wire  _T_1811 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 432:285]
  wire [31:0] _T_1829 = _T_1811 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1844 = _T_1843 | _T_1829; // @[Mux.scala 27:72]
  wire [79:0] _T_1847 = {_T_1684,_T_1764,_T_1844}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1848 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1896 = _T_1848 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1851 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1897 = _T_1851 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1912 = _T_1896 | _T_1897; // @[Mux.scala 27:72]
  wire  _T_1854 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1898 = _T_1854 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1913 = _T_1912 | _T_1898; // @[Mux.scala 27:72]
  wire  _T_1857 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1899 = _T_1857 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1914 = _T_1913 | _T_1899; // @[Mux.scala 27:72]
  wire  _T_1860 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1900 = _T_1860 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1915 = _T_1914 | _T_1900; // @[Mux.scala 27:72]
  wire  _T_1863 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1901 = _T_1863 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1916 = _T_1915 | _T_1901; // @[Mux.scala 27:72]
  wire  _T_1866 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1902 = _T_1866 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1917 = _T_1916 | _T_1902; // @[Mux.scala 27:72]
  wire  _T_1869 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1903 = _T_1869 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1918 = _T_1917 | _T_1903; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1904 = _T_1872 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1919 = _T_1918 | _T_1904; // @[Mux.scala 27:72]
  wire  _T_1875 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1905 = _T_1875 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1920 = _T_1919 | _T_1905; // @[Mux.scala 27:72]
  wire  _T_1878 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1906 = _T_1878 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1921 = _T_1920 | _T_1906; // @[Mux.scala 27:72]
  wire  _T_1881 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1907 = _T_1881 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1922 = _T_1921 | _T_1907; // @[Mux.scala 27:72]
  wire  _T_1884 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1908 = _T_1884 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1923 = _T_1922 | _T_1908; // @[Mux.scala 27:72]
  wire  _T_1887 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1909 = _T_1887 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1924 = _T_1923 | _T_1909; // @[Mux.scala 27:72]
  wire  _T_1890 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1910 = _T_1890 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1925 = _T_1924 | _T_1910; // @[Mux.scala 27:72]
  wire  _T_1893 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 433:73]
  wire [15:0] _T_1911 = _T_1893 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1926 = _T_1925 | _T_1911; // @[Mux.scala 27:72]
  wire [31:0] _T_1976 = _T_1606 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1977 = _T_1609 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1992 = _T_1976 | _T_1977; // @[Mux.scala 27:72]
  wire [31:0] _T_1978 = _T_1612 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1993 = _T_1992 | _T_1978; // @[Mux.scala 27:72]
  wire [31:0] _T_1979 = _T_1615 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1994 = _T_1993 | _T_1979; // @[Mux.scala 27:72]
  wire [31:0] _T_1980 = _T_1618 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1995 = _T_1994 | _T_1980; // @[Mux.scala 27:72]
  wire [31:0] _T_1981 = _T_1621 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1996 = _T_1995 | _T_1981; // @[Mux.scala 27:72]
  wire [31:0] _T_1982 = _T_1624 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1996 | _T_1982; // @[Mux.scala 27:72]
  wire [31:0] _T_1983 = _T_1627 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1997 | _T_1983; // @[Mux.scala 27:72]
  wire [31:0] _T_1984 = _T_1630 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1998 | _T_1984; // @[Mux.scala 27:72]
  wire [31:0] _T_1985 = _T_1633 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1999 | _T_1985; // @[Mux.scala 27:72]
  wire [31:0] _T_1986 = _T_1636 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_2000 | _T_1986; // @[Mux.scala 27:72]
  wire [31:0] _T_1987 = _T_1639 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_2001 | _T_1987; // @[Mux.scala 27:72]
  wire [31:0] _T_1988 = _T_1642 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_2002 | _T_1988; // @[Mux.scala 27:72]
  wire [31:0] _T_1989 = _T_1645 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_2003 | _T_1989; // @[Mux.scala 27:72]
  wire [31:0] _T_1990 = _T_1648 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_2004 | _T_1990; // @[Mux.scala 27:72]
  wire [31:0] _T_1991 = _T_1651 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_2005 | _T_1991; // @[Mux.scala 27:72]
  wire [79:0] _T_2089 = {_T_1926,_T_2006,_T_1764}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_2092 ? _T_1847 : _T_2089; // @[el2_ifu_mem_ctl.scala 431:37]
  wire [79:0] _T_2094 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2092 ? ic_byp_data_only_pre_new : _T_2094; // @[el2_ifu_mem_ctl.scala 435:30]
  wire [79:0] _GEN_793 = {{16'd0}, _T_1256}; // @[el2_ifu_mem_ctl.scala 366:109]
  wire [79:0] _T_1257 = _GEN_793 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 366:109]
  wire [79:0] _GEN_794 = {{16'd0}, _T_1254}; // @[el2_ifu_mem_ctl.scala 366:83]
  wire [79:0] ic_premux_data = _GEN_794 | _T_1257; // @[el2_ifu_mem_ctl.scala 366:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_308; // @[el2_ifu_mem_ctl.scala 373:38]
  wire [1:0] _T_1266 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 377:8]
  wire [7:0] _T_1347 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1352 = ic_miss_buff_data_error[0] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  _T_2601 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 608:47]
  wire  _T_2602 = _T_2601 & _T_13; // @[el2_ifu_mem_ctl.scala 608:50]
  wire  bus_ifu_wr_data_error = _T_2602 & miss_pending; // @[el2_ifu_mem_ctl.scala 608:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1352; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1356 = ic_miss_buff_data_error[1] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1356; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1360 = ic_miss_buff_data_error[2] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1360; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1364 = ic_miss_buff_data_error[3] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1364; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1368 = ic_miss_buff_data_error[4] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1368; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1372 = ic_miss_buff_data_error[5] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1372; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1376 = ic_miss_buff_data_error[6] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1376; // @[el2_ifu_mem_ctl.scala 397:72]
  wire  _T_1380 = ic_miss_buff_data_error[7] & _T_1318; // @[el2_ifu_mem_ctl.scala 398:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1380; // @[el2_ifu_mem_ctl.scala 397:72]
  wire [7:0] _T_1387 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2409 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2417 = _T_6 & _T_308; // @[el2_ifu_mem_ctl.scala 478:65]
  wire  _T_2418 = _T_2417 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 478:88]
  wire  _T_2420 = _T_2418 & _T_2529; // @[el2_ifu_mem_ctl.scala 478:112]
  wire  _T_2421 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2422 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 483:50]
  wire  _T_2424 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2430 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2432 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_38 = _T_2430 | _T_2432; // @[Conditional.scala 39:67]
  wire  _GEN_40 = _T_2424 ? _T_2422 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_2421 ? _T_2422 : _GEN_40; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2409 ? _T_2420 : _GEN_42; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2409 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2423 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 484:56]
  wire  _GEN_43 = _T_2421 & _T_2423; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2409 ? 1'h0 : _GEN_43; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 469:58]
  wire  _T_2406 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 468:49]
  wire  _T_2411 = io_ic_error_start & _T_308; // @[el2_ifu_mem_ctl.scala 477:87]
  wire  _T_2425 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 487:54]
  wire  _T_2426 = _T_2425 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 487:84]
  wire  _T_2435 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 508:66]
  wire  _T_2436 = io_dec_tlu_flush_err_wb & _T_2435; // @[el2_ifu_mem_ctl.scala 508:52]
  wire  _T_2438 = _T_2436 & _T_2529; // @[el2_ifu_mem_ctl.scala 508:81]
  wire  _T_2440 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 511:59]
  wire  _T_2441 = _T_2440 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 511:86]
  wire  _T_2455 = _T_2440 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 514:81]
  wire  _T_2456 = _T_2455 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 514:103]
  wire  _T_2457 = _T_2456 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 514:126]
  wire  _T_2477 = _T_2455 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 521:103]
  wire  _T_2484 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 526:62]
  wire  _T_2485 = io_dec_tlu_flush_lower_wb & _T_2484; // @[el2_ifu_mem_ctl.scala 526:60]
  wire  _T_2486 = _T_2485 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 526:88]
  wire  _T_2487 = _T_2486 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 526:115]
  wire  _GEN_50 = _T_2483 & _T_2441; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_2466 ? _T_2477 : _GEN_50; // @[Conditional.scala 39:67]
  wire  _GEN_55 = _T_2466 | _T_2483; // @[Conditional.scala 39:67]
  wire  _GEN_57 = _T_2439 ? _T_2457 : _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2439 | _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2434 ? _T_2438 : _GEN_57; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2497 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 542:64]
  wire  _T_2499 = _T_2497 & _T_2529; // @[el2_ifu_mem_ctl.scala 542:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2501 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 542:133]
  wire  _T_2502 = _T_2501 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 542:164]
  wire  _T_2503 = _T_2502 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 542:184]
  wire  _T_2504 = _T_2503 & miss_pending; // @[el2_ifu_mem_ctl.scala 542:204]
  wire  _T_2505 = ~_T_2504; // @[el2_ifu_mem_ctl.scala 542:112]
  wire  ifc_bus_ic_req_ff_in = _T_2499 & _T_2505; // @[el2_ifu_mem_ctl.scala 542:110]
  wire  _T_2506 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 543:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 574:45]
  wire  _T_2523 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 577:35]
  wire  _T_2524 = _T_2523 & miss_pending; // @[el2_ifu_mem_ctl.scala 577:53]
  wire  bus_cmd_sent = _T_2524 & _T_2529; // @[el2_ifu_mem_ctl.scala 577:68]
  wire [2:0] _T_2514 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2516 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2518 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 575:51]
  wire  _T_2547 = last_data_recieved_ff & _T_1318; // @[el2_ifu_mem_ctl.scala 585:114]
  wire  last_data_recieved_in = _T_2530 | _T_2547; // @[el2_ifu_mem_ctl.scala 585:89]
  wire [2:0] _T_2553 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 590:45]
  wire  _T_2556 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 591:81]
  wire  _T_2557 = _T_2556 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 591:97]
  wire  _T_2559 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 593:48]
  wire  _T_2560 = _T_2559 & miss_pending; // @[el2_ifu_mem_ctl.scala 593:68]
  wire  bus_inc_cmd_beat_cnt = _T_2560 & _T_2529; // @[el2_ifu_mem_ctl.scala 593:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 595:57]
  wire  _T_2564 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 596:31]
  wire  _T_2566 = ic_act_miss_f | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 596:87]
  wire  _T_2567 = ~_T_2566; // @[el2_ifu_mem_ctl.scala 596:55]
  wire  bus_hold_cmd_beat_cnt = _T_2564 & _T_2567; // @[el2_ifu_mem_ctl.scala 596:53]
  wire  _T_2568 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 597:46]
  wire  bus_cmd_beat_en = _T_2568 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 597:62]
  wire [2:0] _T_2571 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 599:46]
  wire [2:0] _T_2573 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2574 = bus_inc_cmd_beat_cnt ? _T_2571 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2575 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2577 = _T_2573 | _T_2574; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2577 | _T_2575; // @[Mux.scala 27:72]
  wire  _T_2581 = _T_2557 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 600:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 611:62]
  wire  _T_2609 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 616:50]
  wire  _T_2610 = io_ifc_dma_access_ok & _T_2609; // @[el2_ifu_mem_ctl.scala 616:47]
  wire  _T_2611 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 616:70]
  wire  ifc_dma_access_ok_d = _T_2610 & _T_2611; // @[el2_ifu_mem_ctl.scala 616:68]
  wire  _T_2615 = _T_2610 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 617:72]
  wire  _T_2616 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 617:111]
  wire  _T_2617 = _T_2615 & _T_2616; // @[el2_ifu_mem_ctl.scala 617:97]
  wire  ifc_dma_access_q_ok = _T_2617 & _T_2611; // @[el2_ifu_mem_ctl.scala 617:127]
  wire  _T_2620 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 620:40]
  wire  _T_2621 = _T_2620 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 620:58]
  wire  _T_2624 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 621:60]
  wire  _T_2625 = _T_2620 & _T_2624; // @[el2_ifu_mem_ctl.scala 621:58]
  wire  _T_2626 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 621:104]
  wire [2:0] _T_2631 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_2737 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2746 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_2737}; // @[el2_lib.scala 268:22]
  wire  _T_2747 = ^_T_2746; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2755 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2764 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_2755}; // @[el2_lib.scala 268:39]
  wire  _T_2765 = ^_T_2764; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2773 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2782 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_2773}; // @[el2_lib.scala 268:56]
  wire  _T_2783 = ^_T_2782; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2789 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2797 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2789}; // @[el2_lib.scala 268:73]
  wire  _T_2798 = ^_T_2797; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2812 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2789}; // @[el2_lib.scala 268:90]
  wire  _T_2813 = ^_T_2812; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2818 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2819 = ^_T_2818; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2824 = {_T_2747,_T_2765,_T_2783,_T_2798,_T_2813,_T_2819}; // @[Cat.scala 29:58]
  wire  _T_2825 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2826 = ^_T_2824; // @[el2_lib.scala 269:23]
  wire  _T_2827 = _T_2825 ^ _T_2826; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2933 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2942 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2933}; // @[el2_lib.scala 268:22]
  wire  _T_2943 = ^_T_2942; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2951 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2960 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2951}; // @[el2_lib.scala 268:39]
  wire  _T_2961 = ^_T_2960; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2969 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2978 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2969}; // @[el2_lib.scala 268:56]
  wire  _T_2979 = ^_T_2978; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2985 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2993 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2985}; // @[el2_lib.scala 268:73]
  wire  _T_2994 = ^_T_2993; // @[el2_lib.scala 268:80]
  wire [14:0] _T_3008 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2985}; // @[el2_lib.scala 268:90]
  wire  _T_3009 = ^_T_3008; // @[el2_lib.scala 268:97]
  wire [5:0] _T_3014 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_3015 = ^_T_3014; // @[el2_lib.scala 268:114]
  wire [5:0] _T_3020 = {_T_2943,_T_2961,_T_2979,_T_2994,_T_3009,_T_3015}; // @[Cat.scala 29:58]
  wire  _T_3021 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_3022 = ^_T_3020; // @[el2_lib.scala 269:23]
  wire  _T_3023 = _T_3021 ^ _T_3022; // @[el2_lib.scala 269:18]
  wire [6:0] _T_3024 = {_T_3023,_T_2943,_T_2961,_T_2979,_T_2994,_T_3009,_T_3015}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2827,_T_2747,_T_2765,_T_2783,_T_2798,_T_2813,_T_2819,_T_3024}; // @[Cat.scala 29:58]
  wire  _T_3026 = ~_T_2620; // @[el2_ifu_mem_ctl.scala 626:45]
  wire  _T_3027 = iccm_correct_ecc & _T_3026; // @[el2_ifu_mem_ctl.scala 626:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3028 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3035 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 640:53]
  wire  _T_3367 = _T_3279[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3365 = _T_3279[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3363 = _T_3279[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3361 = _T_3279[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3359 = _T_3279[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3357 = _T_3279[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3355 = _T_3279[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3353 = _T_3279[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3351 = _T_3279[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3349 = _T_3279[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3425 = {_T_3367,_T_3365,_T_3363,_T_3361,_T_3359,_T_3357,_T_3355,_T_3353,_T_3351,_T_3349}; // @[el2_lib.scala 310:69]
  wire  _T_3347 = _T_3279[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3345 = _T_3279[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3343 = _T_3279[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3341 = _T_3279[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3339 = _T_3279[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3337 = _T_3279[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3335 = _T_3279[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3333 = _T_3279[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3331 = _T_3279[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3329 = _T_3279[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3416 = {_T_3347,_T_3345,_T_3343,_T_3341,_T_3339,_T_3337,_T_3335,_T_3333,_T_3331,_T_3329}; // @[el2_lib.scala 310:69]
  wire  _T_3327 = _T_3279[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3325 = _T_3279[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3323 = _T_3279[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3321 = _T_3279[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3319 = _T_3279[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3317 = _T_3279[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3315 = _T_3279[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3313 = _T_3279[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3311 = _T_3279[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3309 = _T_3279[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3406 = {_T_3327,_T_3325,_T_3323,_T_3321,_T_3319,_T_3317,_T_3315,_T_3313,_T_3311,_T_3309}; // @[el2_lib.scala 310:69]
  wire  _T_3307 = _T_3279[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3305 = _T_3279[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3303 = _T_3279[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3301 = _T_3279[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3299 = _T_3279[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3297 = _T_3279[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3295 = _T_3279[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3293 = _T_3279[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3291 = _T_3279[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3407 = {_T_3406,_T_3307,_T_3305,_T_3303,_T_3301,_T_3299,_T_3297,_T_3295,_T_3293,_T_3291}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3427 = {_T_3425,_T_3416,_T_3407}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3382 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3388 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3382}; // @[Cat.scala 29:58]
  wire [38:0] _T_3428 = _T_3427 ^ _T_3388; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3429 = _T_3283 ? _T_3428 : _T_3388; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3429[37:32],_T_3429[30:16],_T_3429[14:8],_T_3429[6:4],_T_3429[2]}; // @[Cat.scala 29:58]
  wire  _T_3752 = _T_3664[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_3750 = _T_3664[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_3748 = _T_3664[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_3746 = _T_3664[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_3744 = _T_3664[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_3742 = _T_3664[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_3740 = _T_3664[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_3738 = _T_3664[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_3736 = _T_3664[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_3734 = _T_3664[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3810 = {_T_3752,_T_3750,_T_3748,_T_3746,_T_3744,_T_3742,_T_3740,_T_3738,_T_3736,_T_3734}; // @[el2_lib.scala 310:69]
  wire  _T_3732 = _T_3664[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_3730 = _T_3664[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_3728 = _T_3664[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_3726 = _T_3664[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_3724 = _T_3664[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_3722 = _T_3664[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_3720 = _T_3664[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_3718 = _T_3664[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_3716 = _T_3664[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_3714 = _T_3664[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3801 = {_T_3732,_T_3730,_T_3728,_T_3726,_T_3724,_T_3722,_T_3720,_T_3718,_T_3716,_T_3714}; // @[el2_lib.scala 310:69]
  wire  _T_3712 = _T_3664[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_3710 = _T_3664[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_3708 = _T_3664[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_3706 = _T_3664[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_3704 = _T_3664[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_3702 = _T_3664[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_3700 = _T_3664[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_3698 = _T_3664[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_3696 = _T_3664[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_3694 = _T_3664[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3791 = {_T_3712,_T_3710,_T_3708,_T_3706,_T_3704,_T_3702,_T_3700,_T_3698,_T_3696,_T_3694}; // @[el2_lib.scala 310:69]
  wire  _T_3692 = _T_3664[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_3690 = _T_3664[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_3688 = _T_3664[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_3686 = _T_3664[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_3684 = _T_3664[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_3682 = _T_3664[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_3680 = _T_3664[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_3678 = _T_3664[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_3676 = _T_3664[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3792 = {_T_3791,_T_3692,_T_3690,_T_3688,_T_3686,_T_3684,_T_3682,_T_3680,_T_3678,_T_3676}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3812 = {_T_3810,_T_3801,_T_3792}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_3767 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3773 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3767}; // @[Cat.scala 29:58]
  wire [38:0] _T_3813 = _T_3812 ^ _T_3773; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3814 = _T_3668 ? _T_3813 : _T_3773; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3814[37:32],_T_3814[30:16],_T_3814[14:8],_T_3814[6:4],_T_3814[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 632:35]
  wire  _T_3287 = ~_T_3279[6]; // @[el2_lib.scala 303:55]
  wire  _T_3288 = _T_3281 & _T_3287; // @[el2_lib.scala 303:53]
  wire  _T_3672 = ~_T_3664[6]; // @[el2_lib.scala 303:55]
  wire  _T_3673 = _T_3666 & _T_3672; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_3288,_T_3673}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 634:53]
  wire [63:0] _T_3039 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3040 = {iccm_dma_rdata_1_muxed,_T_3429[37:32],_T_3429[30:16],_T_3429[14:8],_T_3429[6:4],_T_3429[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 636:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 637:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 642:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 646:70]
  wire  _T_3045 = _T_2620 & _T_2609; // @[el2_ifu_mem_ctl.scala 649:65]
  wire  _T_3048 = _T_3026 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 650:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3049 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3051 = _T_3048 ? {{1'd0}, _T_3049} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 650:8]
  wire [31:0] _T_3052 = _T_3045 ? io_dma_mem_addr : {{16'd0}, _T_3051}; // @[el2_ifu_mem_ctl.scala 649:25]
  wire  _T_3441 = _T_3279 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3442 = _T_3429[38] ^ _T_3441; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3442,_T_3429[31],_T_3429[15],_T_3429[7],_T_3429[3],_T_3429[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3826 = _T_3664 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3827 = _T_3814[38] ^ _T_3826; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3827,_T_3814[31],_T_3814[15],_T_3814[7],_T_3814[3],_T_3814[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3843 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 662:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 664:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 665:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 673:62]
  wire  _T_3851 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 667:76]
  wire  _T_3852 = io_iccm_rd_ecc_single_err & _T_3851; // @[el2_ifu_mem_ctl.scala 667:74]
  wire  _T_3854 = _T_3852 & _T_308; // @[el2_ifu_mem_ctl.scala 667:104]
  wire  iccm_ecc_write_status = _T_3854 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 667:127]
  wire  _T_3855 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 668:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3855 & _T_308; // @[el2_ifu_mem_ctl.scala 668:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 672:51]
  wire [13:0] _T_3860 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 671:102]
  wire [38:0] _T_3864 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3869 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 676:41]
  wire  _T_3870 = io_ifc_fetch_req_bf & _T_3869; // @[el2_ifu_mem_ctl.scala 676:39]
  wire  _T_3871 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 676:72]
  wire  _T_3872 = _T_3870 & _T_3871; // @[el2_ifu_mem_ctl.scala 676:70]
  wire  _T_3874 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 677:34]
  wire  _T_3875 = _T_2218 & _T_3874; // @[el2_ifu_mem_ctl.scala 677:32]
  wire  _T_3878 = _T_2233 & _T_3874; // @[el2_ifu_mem_ctl.scala 678:37]
  wire  _T_3879 = _T_3875 | _T_3878; // @[el2_ifu_mem_ctl.scala 677:88]
  wire  _T_3880 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 679:19]
  wire  _T_3882 = _T_3880 & _T_3874; // @[el2_ifu_mem_ctl.scala 679:41]
  wire  _T_3883 = _T_3879 | _T_3882; // @[el2_ifu_mem_ctl.scala 678:88]
  wire  _T_3884 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 680:19]
  wire  _T_3886 = _T_3884 & _T_3874; // @[el2_ifu_mem_ctl.scala 680:35]
  wire  _T_3887 = _T_3883 | _T_3886; // @[el2_ifu_mem_ctl.scala 679:88]
  wire  _T_3890 = _T_2232 & _T_3874; // @[el2_ifu_mem_ctl.scala 681:38]
  wire  _T_3891 = _T_3887 | _T_3890; // @[el2_ifu_mem_ctl.scala 680:88]
  wire  _T_3893 = _T_2233 & miss_state_en; // @[el2_ifu_mem_ctl.scala 682:37]
  wire  _T_3894 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 682:71]
  wire  _T_3895 = _T_3893 & _T_3894; // @[el2_ifu_mem_ctl.scala 682:54]
  wire  _T_3896 = _T_3891 | _T_3895; // @[el2_ifu_mem_ctl.scala 681:57]
  wire  _T_3897 = ~_T_3896; // @[el2_ifu_mem_ctl.scala 677:5]
  wire  _T_3898 = _T_3872 & _T_3897; // @[el2_ifu_mem_ctl.scala 676:96]
  wire  _T_3899 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 683:28]
  wire  _T_3901 = _T_3899 & _T_3869; // @[el2_ifu_mem_ctl.scala 683:50]
  wire  _T_3903 = _T_3901 & _T_3871; // @[el2_ifu_mem_ctl.scala 683:81]
  wire  _T_3912 = ~_T_99; // @[el2_ifu_mem_ctl.scala 686:106]
  wire  _T_3913 = _T_2218 & _T_3912; // @[el2_ifu_mem_ctl.scala 686:104]
  wire  _T_3914 = _T_2233 | _T_3913; // @[el2_ifu_mem_ctl.scala 686:77]
  wire  _T_3918 = ~_T_52; // @[el2_ifu_mem_ctl.scala 686:172]
  wire  _T_3919 = _T_3914 & _T_3918; // @[el2_ifu_mem_ctl.scala 686:170]
  wire  _T_3920 = ~_T_3919; // @[el2_ifu_mem_ctl.scala 686:44]
  wire  _T_3924 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 689:64]
  wire  _T_3925 = ~_T_3924; // @[el2_ifu_mem_ctl.scala 689:50]
  wire  _T_3926 = _T_267 & _T_3925; // @[el2_ifu_mem_ctl.scala 689:48]
  wire  _T_3927 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 689:81]
  wire  ic_valid = _T_3926 & _T_3927; // @[el2_ifu_mem_ctl.scala 689:79]
  wire  _T_3929 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 690:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 693:14]
  wire  _T_3932 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 696:74]
  wire  _T_10074 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 770:45]
  wire  way_status_wr_en = _T_10074 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 770:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3932; // @[el2_ifu_mem_ctl.scala 696:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 698:14]
  wire [2:0] _T_3936 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 702:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 766:41]
  wire  way_status_new = _T_10074 | way_status_hit_new; // @[el2_ifu_mem_ctl.scala 769:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 704:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 706:132]
  wire  _T_3953 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3954 = _T_3953 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3955 = _T_3954 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3957 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3958 = _T_3957 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3959 = _T_3958 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3961 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3962 = _T_3961 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3963 = _T_3962 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3965 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3966 = _T_3965 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3967 = _T_3966 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3969 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3970 = _T_3969 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3971 = _T_3970 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3973 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3974 = _T_3973 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3975 = _T_3974 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3977 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3978 = _T_3977 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3979 = _T_3978 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3981 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 710:93]
  wire  _T_3982 = _T_3981 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 710:102]
  wire  _T_3983 = _T_3982 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3987 = _T_3954 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3991 = _T_3958 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3995 = _T_3962 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_3999 = _T_3966 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4003 = _T_3970 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4007 = _T_3974 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4011 = _T_3978 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4015 = _T_3982 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4019 = _T_3954 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4023 = _T_3958 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4027 = _T_3962 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4031 = _T_3966 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4035 = _T_3970 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4039 = _T_3974 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4043 = _T_3978 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4047 = _T_3982 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4051 = _T_3954 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4055 = _T_3958 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4059 = _T_3962 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4063 = _T_3966 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4067 = _T_3970 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4071 = _T_3974 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4075 = _T_3978 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4079 = _T_3982 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4083 = _T_3954 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4087 = _T_3958 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4091 = _T_3962 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4095 = _T_3966 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4099 = _T_3970 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4103 = _T_3974 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4107 = _T_3978 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4111 = _T_3982 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4115 = _T_3954 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4119 = _T_3958 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4123 = _T_3962 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4127 = _T_3966 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4131 = _T_3970 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4135 = _T_3974 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4139 = _T_3978 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4143 = _T_3982 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4147 = _T_3954 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4151 = _T_3958 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4155 = _T_3962 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4159 = _T_3966 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4163 = _T_3970 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4167 = _T_3974 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4171 = _T_3978 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4175 = _T_3982 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4179 = _T_3954 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4183 = _T_3958 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4187 = _T_3962 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4191 = _T_3966 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4195 = _T_3970 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4199 = _T_3974 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4203 = _T_3978 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4207 = _T_3982 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4211 = _T_3954 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4215 = _T_3958 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4219 = _T_3962 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4223 = _T_3966 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4227 = _T_3970 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4231 = _T_3974 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4235 = _T_3978 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4239 = _T_3982 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4243 = _T_3954 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4247 = _T_3958 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4251 = _T_3962 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4255 = _T_3966 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4259 = _T_3970 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4263 = _T_3974 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4267 = _T_3978 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4271 = _T_3982 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4275 = _T_3954 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4279 = _T_3958 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4283 = _T_3962 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4287 = _T_3966 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4291 = _T_3970 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4295 = _T_3974 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4299 = _T_3978 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4303 = _T_3982 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4307 = _T_3954 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4311 = _T_3958 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4315 = _T_3962 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4319 = _T_3966 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4323 = _T_3970 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4327 = _T_3974 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4331 = _T_3978 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4335 = _T_3982 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4339 = _T_3954 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4343 = _T_3958 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4347 = _T_3962 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4351 = _T_3966 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4355 = _T_3970 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4359 = _T_3974 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4363 = _T_3978 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4367 = _T_3982 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4371 = _T_3954 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4375 = _T_3958 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4379 = _T_3962 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4383 = _T_3966 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4387 = _T_3970 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4391 = _T_3974 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4395 = _T_3978 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4399 = _T_3982 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4403 = _T_3954 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4407 = _T_3958 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4411 = _T_3962 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4415 = _T_3966 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4419 = _T_3970 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4423 = _T_3974 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4427 = _T_3978 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4431 = _T_3982 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4435 = _T_3954 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4439 = _T_3958 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4443 = _T_3962 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4447 = _T_3966 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4451 = _T_3970 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4455 = _T_3974 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4459 = _T_3978 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_4463 = _T_3982 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 710:124]
  wire  _T_10079 = _T_91 & miss_pending; // @[el2_ifu_mem_ctl.scala 773:108]
  wire  bus_wren_last_0 = _T_10079 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 773:123]
  wire  _T_10082 = bus_wren_last_0 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 775:73]
  wire [1:0] ifu_tag_wren = {1'h0,_T_10082}; // @[Cat.scala 29:58]
  wire [1:0] _T_10117 = _T_3932 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10117 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 806:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 719:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 721:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 725:14]
  wire  _T_5112 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 729:82]
  wire  _T_5114 = _T_5112 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5116 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 730:74]
  wire  _T_5118 = _T_5116 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5119 = _T_5114 | _T_5118; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5120 = _T_5119 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire  _T_5124 = _T_5112 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5128 = _T_5116 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5129 = _T_5124 | _T_5128; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5130 = _T_5129 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire [1:0] tag_valid_clken_0 = {_T_5120,_T_5130}; // @[Cat.scala 29:58]
  wire  _T_5132 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 729:82]
  wire  _T_5134 = _T_5132 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5136 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 730:74]
  wire  _T_5138 = _T_5136 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5139 = _T_5134 | _T_5138; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5140 = _T_5139 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire  _T_5144 = _T_5132 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5148 = _T_5136 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5149 = _T_5144 | _T_5148; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5150 = _T_5149 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire [1:0] tag_valid_clken_1 = {_T_5140,_T_5150}; // @[Cat.scala 29:58]
  wire  _T_5152 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 729:82]
  wire  _T_5154 = _T_5152 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5156 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 730:74]
  wire  _T_5158 = _T_5156 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5159 = _T_5154 | _T_5158; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5160 = _T_5159 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire  _T_5164 = _T_5152 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5168 = _T_5156 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5169 = _T_5164 | _T_5168; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5170 = _T_5169 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire [1:0] tag_valid_clken_2 = {_T_5160,_T_5170}; // @[Cat.scala 29:58]
  wire  _T_5172 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 729:82]
  wire  _T_5174 = _T_5172 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5176 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 730:74]
  wire  _T_5178 = _T_5176 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5179 = _T_5174 | _T_5178; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5180 = _T_5179 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire  _T_5184 = _T_5172 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 729:91]
  wire  _T_5188 = _T_5176 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 730:83]
  wire  _T_5189 = _T_5184 | _T_5188; // @[el2_ifu_mem_ctl.scala 729:113]
  wire  _T_5190 = _T_5189 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 730:106]
  wire [1:0] tag_valid_clken_3 = {_T_5180,_T_5190}; // @[Cat.scala 29:58]
  wire  _T_5193 = ic_valid_ff & _T_186; // @[el2_ifu_mem_ctl.scala 735:64]
  wire  _T_5194 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 735:91]
  wire  _T_5195 = _T_5193 & _T_5194; // @[el2_ifu_mem_ctl.scala 735:89]
  wire  _T_5198 = _T_4465 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5199 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5201 = _T_5199 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5203 = _T_5201 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5204 = _T_5198 | _T_5203; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5214 = _T_4469 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5215 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5217 = _T_5215 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5219 = _T_5217 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5220 = _T_5214 | _T_5219; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5230 = _T_4473 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5231 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5233 = _T_5231 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5235 = _T_5233 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5236 = _T_5230 | _T_5235; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5246 = _T_4477 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5247 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5249 = _T_5247 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5251 = _T_5249 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5252 = _T_5246 | _T_5251; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5262 = _T_4481 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5263 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5265 = _T_5263 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5267 = _T_5265 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5268 = _T_5262 | _T_5267; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5278 = _T_4485 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5279 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5281 = _T_5279 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5283 = _T_5281 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5284 = _T_5278 | _T_5283; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5294 = _T_4489 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5295 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5297 = _T_5295 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5299 = _T_5297 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5300 = _T_5294 | _T_5299; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5310 = _T_4493 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5311 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5313 = _T_5311 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5315 = _T_5313 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5316 = _T_5310 | _T_5315; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5326 = _T_4497 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5327 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5329 = _T_5327 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5331 = _T_5329 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5332 = _T_5326 | _T_5331; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5342 = _T_4501 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5343 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5345 = _T_5343 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5347 = _T_5345 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5348 = _T_5342 | _T_5347; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5358 = _T_4505 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5359 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5361 = _T_5359 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5363 = _T_5361 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5364 = _T_5358 | _T_5363; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5374 = _T_4509 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5375 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5377 = _T_5375 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5379 = _T_5377 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5380 = _T_5374 | _T_5379; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5390 = _T_4513 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5391 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5393 = _T_5391 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5395 = _T_5393 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5396 = _T_5390 | _T_5395; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5406 = _T_4517 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5407 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5409 = _T_5407 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5411 = _T_5409 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5412 = _T_5406 | _T_5411; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5422 = _T_4521 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5423 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5425 = _T_5423 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5427 = _T_5425 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5428 = _T_5422 | _T_5427; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5438 = _T_4525 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5439 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5441 = _T_5439 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5443 = _T_5441 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5444 = _T_5438 | _T_5443; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5454 = _T_4529 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5455 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5457 = _T_5455 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5459 = _T_5457 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5460 = _T_5454 | _T_5459; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5470 = _T_4533 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5471 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5473 = _T_5471 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5475 = _T_5473 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5476 = _T_5470 | _T_5475; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5486 = _T_4537 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5487 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5489 = _T_5487 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5491 = _T_5489 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5492 = _T_5486 | _T_5491; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5502 = _T_4541 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5503 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5505 = _T_5503 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5507 = _T_5505 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5508 = _T_5502 | _T_5507; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5518 = _T_4545 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5519 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5521 = _T_5519 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5523 = _T_5521 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5524 = _T_5518 | _T_5523; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5534 = _T_4549 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5535 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5537 = _T_5535 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5539 = _T_5537 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5540 = _T_5534 | _T_5539; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5550 = _T_4553 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5551 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5553 = _T_5551 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5555 = _T_5553 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5556 = _T_5550 | _T_5555; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5566 = _T_4557 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5567 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5569 = _T_5567 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5571 = _T_5569 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5572 = _T_5566 | _T_5571; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5582 = _T_4561 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5583 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5585 = _T_5583 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5587 = _T_5585 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5588 = _T_5582 | _T_5587; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5598 = _T_4565 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5599 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5601 = _T_5599 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5603 = _T_5601 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5604 = _T_5598 | _T_5603; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5614 = _T_4569 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5615 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5617 = _T_5615 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5619 = _T_5617 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5620 = _T_5614 | _T_5619; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5630 = _T_4573 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5631 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5633 = _T_5631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5635 = _T_5633 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5636 = _T_5630 | _T_5635; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5646 = _T_4577 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5647 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5649 = _T_5647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5651 = _T_5649 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5652 = _T_5646 | _T_5651; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5662 = _T_4581 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5663 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5665 = _T_5663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5667 = _T_5665 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5668 = _T_5662 | _T_5667; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5678 = _T_4585 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5679 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5681 = _T_5679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5683 = _T_5681 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5684 = _T_5678 | _T_5683; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5694 = _T_4589 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5695 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_5697 = _T_5695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5699 = _T_5697 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5700 = _T_5694 | _T_5699; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5710 = _T_4465 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5713 = _T_5199 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5715 = _T_5713 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5716 = _T_5710 | _T_5715; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5726 = _T_4469 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5729 = _T_5215 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5731 = _T_5729 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5732 = _T_5726 | _T_5731; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5742 = _T_4473 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5745 = _T_5231 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5747 = _T_5745 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5748 = _T_5742 | _T_5747; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5758 = _T_4477 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5761 = _T_5247 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5763 = _T_5761 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5764 = _T_5758 | _T_5763; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5774 = _T_4481 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5777 = _T_5263 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5779 = _T_5777 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5780 = _T_5774 | _T_5779; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5790 = _T_4485 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5793 = _T_5279 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5795 = _T_5793 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5796 = _T_5790 | _T_5795; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5806 = _T_4489 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5809 = _T_5295 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5811 = _T_5809 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5812 = _T_5806 | _T_5811; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5822 = _T_4493 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5825 = _T_5311 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5827 = _T_5825 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5828 = _T_5822 | _T_5827; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5838 = _T_4497 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5841 = _T_5327 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5843 = _T_5841 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5844 = _T_5838 | _T_5843; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5854 = _T_4501 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5857 = _T_5343 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5859 = _T_5857 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5860 = _T_5854 | _T_5859; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5870 = _T_4505 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5873 = _T_5359 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5875 = _T_5873 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5876 = _T_5870 | _T_5875; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5886 = _T_4509 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5889 = _T_5375 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5891 = _T_5889 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5892 = _T_5886 | _T_5891; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5902 = _T_4513 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5905 = _T_5391 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5907 = _T_5905 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5908 = _T_5902 | _T_5907; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5918 = _T_4517 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5921 = _T_5407 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5923 = _T_5921 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5924 = _T_5918 | _T_5923; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5934 = _T_4521 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5937 = _T_5423 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5939 = _T_5937 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5940 = _T_5934 | _T_5939; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5950 = _T_4525 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5953 = _T_5439 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5955 = _T_5953 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5956 = _T_5950 | _T_5955; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5966 = _T_4529 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5969 = _T_5455 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5971 = _T_5969 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5972 = _T_5966 | _T_5971; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5982 = _T_4533 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_5985 = _T_5471 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_5987 = _T_5985 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_5988 = _T_5982 | _T_5987; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_5998 = _T_4537 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6001 = _T_5487 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6003 = _T_6001 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6004 = _T_5998 | _T_6003; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6014 = _T_4541 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6017 = _T_5503 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6019 = _T_6017 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6020 = _T_6014 | _T_6019; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6030 = _T_4545 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6033 = _T_5519 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6035 = _T_6033 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6036 = _T_6030 | _T_6035; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6046 = _T_4549 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6049 = _T_5535 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6051 = _T_6049 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6052 = _T_6046 | _T_6051; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6062 = _T_4553 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6065 = _T_5551 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6067 = _T_6065 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6068 = _T_6062 | _T_6067; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6078 = _T_4557 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6081 = _T_5567 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6083 = _T_6081 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6084 = _T_6078 | _T_6083; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6094 = _T_4561 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6097 = _T_5583 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6099 = _T_6097 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6100 = _T_6094 | _T_6099; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6110 = _T_4565 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6113 = _T_5599 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6115 = _T_6113 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6116 = _T_6110 | _T_6115; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6126 = _T_4569 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6129 = _T_5615 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6131 = _T_6129 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6132 = _T_6126 | _T_6131; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6142 = _T_4573 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6145 = _T_5631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6147 = _T_6145 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6148 = _T_6142 | _T_6147; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6158 = _T_4577 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6161 = _T_5647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6163 = _T_6161 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6164 = _T_6158 | _T_6163; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6174 = _T_4581 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6177 = _T_5663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6179 = _T_6177 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6180 = _T_6174 | _T_6179; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6190 = _T_4585 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6193 = _T_5679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6195 = _T_6193 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6196 = _T_6190 | _T_6195; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6206 = _T_4589 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6209 = _T_5695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6211 = _T_6209 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6212 = _T_6206 | _T_6211; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6222 = _T_4593 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6223 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6225 = _T_6223 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6227 = _T_6225 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6228 = _T_6222 | _T_6227; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6238 = _T_4597 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6239 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6241 = _T_6239 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6243 = _T_6241 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6244 = _T_6238 | _T_6243; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6254 = _T_4601 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6255 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6257 = _T_6255 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6259 = _T_6257 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6260 = _T_6254 | _T_6259; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6270 = _T_4605 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6271 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6273 = _T_6271 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6275 = _T_6273 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6276 = _T_6270 | _T_6275; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6286 = _T_4609 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6287 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6289 = _T_6287 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6291 = _T_6289 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6292 = _T_6286 | _T_6291; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6302 = _T_4613 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6303 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6305 = _T_6303 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6307 = _T_6305 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6308 = _T_6302 | _T_6307; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6318 = _T_4617 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6319 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6321 = _T_6319 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6323 = _T_6321 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6324 = _T_6318 | _T_6323; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6334 = _T_4621 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6335 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6337 = _T_6335 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6339 = _T_6337 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6340 = _T_6334 | _T_6339; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6350 = _T_4625 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6351 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6353 = _T_6351 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6355 = _T_6353 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6356 = _T_6350 | _T_6355; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6366 = _T_4629 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6367 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6369 = _T_6367 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6371 = _T_6369 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6372 = _T_6366 | _T_6371; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6382 = _T_4633 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6383 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6385 = _T_6383 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6387 = _T_6385 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6388 = _T_6382 | _T_6387; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6398 = _T_4637 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6399 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6401 = _T_6399 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6403 = _T_6401 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6404 = _T_6398 | _T_6403; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6414 = _T_4641 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6415 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6417 = _T_6415 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6419 = _T_6417 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6420 = _T_6414 | _T_6419; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6430 = _T_4645 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6431 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6433 = _T_6431 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6435 = _T_6433 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6436 = _T_6430 | _T_6435; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6446 = _T_4649 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6447 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6449 = _T_6447 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6451 = _T_6449 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6452 = _T_6446 | _T_6451; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6462 = _T_4653 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6463 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6465 = _T_6463 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6467 = _T_6465 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6468 = _T_6462 | _T_6467; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6478 = _T_4657 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6479 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6481 = _T_6479 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6483 = _T_6481 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6484 = _T_6478 | _T_6483; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6494 = _T_4661 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6495 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6497 = _T_6495 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6499 = _T_6497 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6500 = _T_6494 | _T_6499; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6510 = _T_4665 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6511 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6513 = _T_6511 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6515 = _T_6513 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6516 = _T_6510 | _T_6515; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6526 = _T_4669 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6527 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6529 = _T_6527 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6531 = _T_6529 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6532 = _T_6526 | _T_6531; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6542 = _T_4673 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6543 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6545 = _T_6543 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6547 = _T_6545 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6548 = _T_6542 | _T_6547; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6558 = _T_4677 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6559 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6561 = _T_6559 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6563 = _T_6561 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6564 = _T_6558 | _T_6563; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6574 = _T_4681 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6575 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6577 = _T_6575 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6579 = _T_6577 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6580 = _T_6574 | _T_6579; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6590 = _T_4685 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6591 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6593 = _T_6591 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6595 = _T_6593 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6596 = _T_6590 | _T_6595; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6606 = _T_4689 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6607 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6609 = _T_6607 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6611 = _T_6609 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6612 = _T_6606 | _T_6611; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6622 = _T_4693 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6623 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6625 = _T_6623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6627 = _T_6625 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6628 = _T_6622 | _T_6627; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6638 = _T_4697 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6639 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6641 = _T_6639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6643 = _T_6641 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6644 = _T_6638 | _T_6643; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6654 = _T_4701 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6655 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6657 = _T_6655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6659 = _T_6657 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6660 = _T_6654 | _T_6659; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6670 = _T_4705 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6671 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6673 = _T_6671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6675 = _T_6673 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6676 = _T_6670 | _T_6675; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6686 = _T_4709 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6687 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6689 = _T_6687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6691 = _T_6689 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6692 = _T_6686 | _T_6691; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6702 = _T_4713 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6703 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6705 = _T_6703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6707 = _T_6705 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6708 = _T_6702 | _T_6707; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6718 = _T_4717 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6719 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_6721 = _T_6719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6723 = _T_6721 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6724 = _T_6718 | _T_6723; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6734 = _T_4593 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6737 = _T_6223 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6739 = _T_6737 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6740 = _T_6734 | _T_6739; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6750 = _T_4597 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6753 = _T_6239 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6755 = _T_6753 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6756 = _T_6750 | _T_6755; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6766 = _T_4601 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6769 = _T_6255 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6771 = _T_6769 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6772 = _T_6766 | _T_6771; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6782 = _T_4605 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6785 = _T_6271 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6787 = _T_6785 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6788 = _T_6782 | _T_6787; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6798 = _T_4609 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6801 = _T_6287 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6803 = _T_6801 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6804 = _T_6798 | _T_6803; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6814 = _T_4613 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6817 = _T_6303 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6819 = _T_6817 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6820 = _T_6814 | _T_6819; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6830 = _T_4617 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6833 = _T_6319 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6835 = _T_6833 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6836 = _T_6830 | _T_6835; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6846 = _T_4621 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6849 = _T_6335 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6851 = _T_6849 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6852 = _T_6846 | _T_6851; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6862 = _T_4625 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6865 = _T_6351 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6867 = _T_6865 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6868 = _T_6862 | _T_6867; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6878 = _T_4629 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6881 = _T_6367 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6883 = _T_6881 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6884 = _T_6878 | _T_6883; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6894 = _T_4633 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6897 = _T_6383 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6899 = _T_6897 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6900 = _T_6894 | _T_6899; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6910 = _T_4637 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6913 = _T_6399 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6915 = _T_6913 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6916 = _T_6910 | _T_6915; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6926 = _T_4641 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6929 = _T_6415 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6931 = _T_6929 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6932 = _T_6926 | _T_6931; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6942 = _T_4645 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6945 = _T_6431 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6947 = _T_6945 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6948 = _T_6942 | _T_6947; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6958 = _T_4649 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6961 = _T_6447 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6963 = _T_6961 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6964 = _T_6958 | _T_6963; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6974 = _T_4653 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6977 = _T_6463 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6979 = _T_6977 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6980 = _T_6974 | _T_6979; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_6990 = _T_4657 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_6993 = _T_6479 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_6995 = _T_6993 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_6996 = _T_6990 | _T_6995; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7006 = _T_4661 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7009 = _T_6495 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7011 = _T_7009 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7012 = _T_7006 | _T_7011; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7022 = _T_4665 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7025 = _T_6511 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7027 = _T_7025 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7028 = _T_7022 | _T_7027; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7038 = _T_4669 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7041 = _T_6527 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7043 = _T_7041 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7044 = _T_7038 | _T_7043; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7054 = _T_4673 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7057 = _T_6543 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7059 = _T_7057 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7060 = _T_7054 | _T_7059; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7070 = _T_4677 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7073 = _T_6559 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7075 = _T_7073 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7076 = _T_7070 | _T_7075; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7086 = _T_4681 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7089 = _T_6575 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7091 = _T_7089 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7092 = _T_7086 | _T_7091; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7102 = _T_4685 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7105 = _T_6591 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7107 = _T_7105 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7108 = _T_7102 | _T_7107; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7118 = _T_4689 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7121 = _T_6607 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7123 = _T_7121 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7124 = _T_7118 | _T_7123; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7134 = _T_4693 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7137 = _T_6623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7139 = _T_7137 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7140 = _T_7134 | _T_7139; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7150 = _T_4697 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7153 = _T_6639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7155 = _T_7153 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7156 = _T_7150 | _T_7155; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7166 = _T_4701 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7169 = _T_6655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7171 = _T_7169 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7172 = _T_7166 | _T_7171; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7182 = _T_4705 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7185 = _T_6671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7187 = _T_7185 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7188 = _T_7182 | _T_7187; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7198 = _T_4709 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7201 = _T_6687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7203 = _T_7201 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7204 = _T_7198 | _T_7203; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7214 = _T_4713 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7217 = _T_6703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7219 = _T_7217 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7220 = _T_7214 | _T_7219; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7230 = _T_4717 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7233 = _T_6719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7235 = _T_7233 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7236 = _T_7230 | _T_7235; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7246 = _T_4721 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire [6:0] _GEN_796 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7247 = _GEN_796 == 7'h40; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7249 = _T_7247 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7251 = _T_7249 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7252 = _T_7246 | _T_7251; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7262 = _T_4725 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7263 = _GEN_796 == 7'h41; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7265 = _T_7263 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7267 = _T_7265 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7268 = _T_7262 | _T_7267; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7278 = _T_4729 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7279 = _GEN_796 == 7'h42; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7281 = _T_7279 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7283 = _T_7281 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7284 = _T_7278 | _T_7283; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7294 = _T_4733 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7295 = _GEN_796 == 7'h43; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7297 = _T_7295 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7299 = _T_7297 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7300 = _T_7294 | _T_7299; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7310 = _T_4737 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7311 = _GEN_796 == 7'h44; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7313 = _T_7311 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7315 = _T_7313 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7316 = _T_7310 | _T_7315; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7326 = _T_4741 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7327 = _GEN_796 == 7'h45; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7329 = _T_7327 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7331 = _T_7329 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7332 = _T_7326 | _T_7331; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7342 = _T_4745 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7343 = _GEN_796 == 7'h46; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7345 = _T_7343 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7347 = _T_7345 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7348 = _T_7342 | _T_7347; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7358 = _T_4749 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7359 = _GEN_796 == 7'h47; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7361 = _T_7359 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7363 = _T_7361 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7364 = _T_7358 | _T_7363; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7374 = _T_4753 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7375 = _GEN_796 == 7'h48; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7377 = _T_7375 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7379 = _T_7377 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7380 = _T_7374 | _T_7379; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7390 = _T_4757 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7391 = _GEN_796 == 7'h49; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7393 = _T_7391 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7395 = _T_7393 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7396 = _T_7390 | _T_7395; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7406 = _T_4761 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7407 = _GEN_796 == 7'h4a; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7409 = _T_7407 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7411 = _T_7409 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7412 = _T_7406 | _T_7411; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7422 = _T_4765 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7423 = _GEN_796 == 7'h4b; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7425 = _T_7423 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7427 = _T_7425 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7428 = _T_7422 | _T_7427; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7438 = _T_4769 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7439 = _GEN_796 == 7'h4c; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7441 = _T_7439 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7443 = _T_7441 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7444 = _T_7438 | _T_7443; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7454 = _T_4773 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7455 = _GEN_796 == 7'h4d; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7457 = _T_7455 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7459 = _T_7457 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7460 = _T_7454 | _T_7459; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7470 = _T_4777 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7471 = _GEN_796 == 7'h4e; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7473 = _T_7471 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7475 = _T_7473 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7476 = _T_7470 | _T_7475; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7486 = _T_4781 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7487 = _GEN_796 == 7'h4f; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7489 = _T_7487 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7491 = _T_7489 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7492 = _T_7486 | _T_7491; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7502 = _T_4785 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7503 = _GEN_796 == 7'h50; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7505 = _T_7503 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7507 = _T_7505 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7508 = _T_7502 | _T_7507; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7518 = _T_4789 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7519 = _GEN_796 == 7'h51; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7521 = _T_7519 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7523 = _T_7521 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7524 = _T_7518 | _T_7523; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7534 = _T_4793 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7535 = _GEN_796 == 7'h52; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7537 = _T_7535 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7539 = _T_7537 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7540 = _T_7534 | _T_7539; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7550 = _T_4797 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7551 = _GEN_796 == 7'h53; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7553 = _T_7551 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7555 = _T_7553 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7556 = _T_7550 | _T_7555; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7566 = _T_4801 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7567 = _GEN_796 == 7'h54; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7569 = _T_7567 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7571 = _T_7569 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7572 = _T_7566 | _T_7571; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7582 = _T_4805 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7583 = _GEN_796 == 7'h55; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7585 = _T_7583 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7587 = _T_7585 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7588 = _T_7582 | _T_7587; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7598 = _T_4809 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7599 = _GEN_796 == 7'h56; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7601 = _T_7599 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7603 = _T_7601 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7604 = _T_7598 | _T_7603; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7614 = _T_4813 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7615 = _GEN_796 == 7'h57; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7617 = _T_7615 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7619 = _T_7617 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7620 = _T_7614 | _T_7619; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7630 = _T_4817 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7631 = _GEN_796 == 7'h58; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7633 = _T_7631 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7635 = _T_7633 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7636 = _T_7630 | _T_7635; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7646 = _T_4821 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7647 = _GEN_796 == 7'h59; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7649 = _T_7647 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7651 = _T_7649 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7652 = _T_7646 | _T_7651; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7662 = _T_4825 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7663 = _GEN_796 == 7'h5a; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7665 = _T_7663 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7667 = _T_7665 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7668 = _T_7662 | _T_7667; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7678 = _T_4829 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7679 = _GEN_796 == 7'h5b; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7681 = _T_7679 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7683 = _T_7681 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7684 = _T_7678 | _T_7683; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7694 = _T_4833 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7695 = _GEN_796 == 7'h5c; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7697 = _T_7695 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7699 = _T_7697 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7700 = _T_7694 | _T_7699; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7710 = _T_4837 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7711 = _GEN_796 == 7'h5d; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7713 = _T_7711 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7715 = _T_7713 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7716 = _T_7710 | _T_7715; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7726 = _T_4841 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7727 = _GEN_796 == 7'h5e; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7729 = _T_7727 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7731 = _T_7729 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7732 = _T_7726 | _T_7731; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7742 = _T_4845 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7743 = _GEN_796 == 7'h5f; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_7745 = _T_7743 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7747 = _T_7745 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7748 = _T_7742 | _T_7747; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7758 = _T_4721 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7761 = _T_7247 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7763 = _T_7761 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7764 = _T_7758 | _T_7763; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7774 = _T_4725 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7777 = _T_7263 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7779 = _T_7777 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7780 = _T_7774 | _T_7779; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7790 = _T_4729 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7793 = _T_7279 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7795 = _T_7793 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7796 = _T_7790 | _T_7795; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7806 = _T_4733 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7809 = _T_7295 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7811 = _T_7809 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7812 = _T_7806 | _T_7811; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7822 = _T_4737 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7825 = _T_7311 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7827 = _T_7825 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7828 = _T_7822 | _T_7827; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7838 = _T_4741 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7841 = _T_7327 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7843 = _T_7841 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7844 = _T_7838 | _T_7843; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7854 = _T_4745 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7857 = _T_7343 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7859 = _T_7857 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7860 = _T_7854 | _T_7859; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7870 = _T_4749 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7873 = _T_7359 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7875 = _T_7873 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7876 = _T_7870 | _T_7875; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7886 = _T_4753 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7889 = _T_7375 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7891 = _T_7889 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7892 = _T_7886 | _T_7891; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7902 = _T_4757 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7905 = _T_7391 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7907 = _T_7905 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7908 = _T_7902 | _T_7907; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7918 = _T_4761 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7921 = _T_7407 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7923 = _T_7921 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7924 = _T_7918 | _T_7923; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7934 = _T_4765 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7937 = _T_7423 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7939 = _T_7937 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7940 = _T_7934 | _T_7939; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7950 = _T_4769 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7953 = _T_7439 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7955 = _T_7953 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7956 = _T_7950 | _T_7955; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7966 = _T_4773 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7969 = _T_7455 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7971 = _T_7969 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7972 = _T_7966 | _T_7971; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7982 = _T_4777 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_7985 = _T_7471 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_7987 = _T_7985 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_7988 = _T_7982 | _T_7987; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_7998 = _T_4781 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8001 = _T_7487 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8003 = _T_8001 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8004 = _T_7998 | _T_8003; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8014 = _T_4785 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8017 = _T_7503 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8019 = _T_8017 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8020 = _T_8014 | _T_8019; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8030 = _T_4789 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8033 = _T_7519 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8035 = _T_8033 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8036 = _T_8030 | _T_8035; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8046 = _T_4793 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8049 = _T_7535 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8051 = _T_8049 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8052 = _T_8046 | _T_8051; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8062 = _T_4797 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8065 = _T_7551 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8067 = _T_8065 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8068 = _T_8062 | _T_8067; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8078 = _T_4801 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8081 = _T_7567 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8083 = _T_8081 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8084 = _T_8078 | _T_8083; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8094 = _T_4805 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8097 = _T_7583 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8099 = _T_8097 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8100 = _T_8094 | _T_8099; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8110 = _T_4809 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8113 = _T_7599 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8115 = _T_8113 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8116 = _T_8110 | _T_8115; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8126 = _T_4813 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8129 = _T_7615 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8131 = _T_8129 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8132 = _T_8126 | _T_8131; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8142 = _T_4817 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8145 = _T_7631 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8147 = _T_8145 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8148 = _T_8142 | _T_8147; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8158 = _T_4821 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8161 = _T_7647 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8163 = _T_8161 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8164 = _T_8158 | _T_8163; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8174 = _T_4825 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8177 = _T_7663 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8179 = _T_8177 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8180 = _T_8174 | _T_8179; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8190 = _T_4829 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8193 = _T_7679 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8195 = _T_8193 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8196 = _T_8190 | _T_8195; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8206 = _T_4833 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8209 = _T_7695 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8211 = _T_8209 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8212 = _T_8206 | _T_8211; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8222 = _T_4837 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8225 = _T_7711 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8227 = _T_8225 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8228 = _T_8222 | _T_8227; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8238 = _T_4841 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8241 = _T_7727 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8243 = _T_8241 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8244 = _T_8238 | _T_8243; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8254 = _T_4845 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8257 = _T_7743 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8259 = _T_8257 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8260 = _T_8254 | _T_8259; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8270 = _T_4849 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8271 = _GEN_796 == 7'h60; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8273 = _T_8271 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8275 = _T_8273 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8276 = _T_8270 | _T_8275; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8286 = _T_4853 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8287 = _GEN_796 == 7'h61; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8289 = _T_8287 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8291 = _T_8289 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8292 = _T_8286 | _T_8291; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8302 = _T_4857 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8303 = _GEN_796 == 7'h62; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8305 = _T_8303 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8307 = _T_8305 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8308 = _T_8302 | _T_8307; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8318 = _T_4861 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8319 = _GEN_796 == 7'h63; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8321 = _T_8319 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8323 = _T_8321 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8324 = _T_8318 | _T_8323; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8334 = _T_4865 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8335 = _GEN_796 == 7'h64; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8337 = _T_8335 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8339 = _T_8337 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8340 = _T_8334 | _T_8339; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8350 = _T_4869 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8351 = _GEN_796 == 7'h65; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8353 = _T_8351 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8355 = _T_8353 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8356 = _T_8350 | _T_8355; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8366 = _T_4873 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8367 = _GEN_796 == 7'h66; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8369 = _T_8367 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8371 = _T_8369 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8372 = _T_8366 | _T_8371; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8382 = _T_4877 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8383 = _GEN_796 == 7'h67; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8385 = _T_8383 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8387 = _T_8385 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8388 = _T_8382 | _T_8387; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8398 = _T_4881 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8399 = _GEN_796 == 7'h68; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8401 = _T_8399 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8403 = _T_8401 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8404 = _T_8398 | _T_8403; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8414 = _T_4885 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8415 = _GEN_796 == 7'h69; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8417 = _T_8415 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8419 = _T_8417 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8420 = _T_8414 | _T_8419; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8430 = _T_4889 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8431 = _GEN_796 == 7'h6a; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8433 = _T_8431 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8435 = _T_8433 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8436 = _T_8430 | _T_8435; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8446 = _T_4893 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8447 = _GEN_796 == 7'h6b; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8449 = _T_8447 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8451 = _T_8449 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8452 = _T_8446 | _T_8451; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8462 = _T_4897 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8463 = _GEN_796 == 7'h6c; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8465 = _T_8463 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8467 = _T_8465 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8468 = _T_8462 | _T_8467; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8478 = _T_4901 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8479 = _GEN_796 == 7'h6d; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8481 = _T_8479 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8483 = _T_8481 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8484 = _T_8478 | _T_8483; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8494 = _T_4905 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8495 = _GEN_796 == 7'h6e; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8497 = _T_8495 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8499 = _T_8497 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8500 = _T_8494 | _T_8499; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8510 = _T_4909 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8511 = _GEN_796 == 7'h6f; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8513 = _T_8511 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8515 = _T_8513 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8516 = _T_8510 | _T_8515; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8526 = _T_4913 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8527 = _GEN_796 == 7'h70; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8529 = _T_8527 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8531 = _T_8529 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8532 = _T_8526 | _T_8531; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8542 = _T_4917 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8543 = _GEN_796 == 7'h71; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8545 = _T_8543 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8547 = _T_8545 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8548 = _T_8542 | _T_8547; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8558 = _T_4921 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8559 = _GEN_796 == 7'h72; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8561 = _T_8559 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8563 = _T_8561 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8564 = _T_8558 | _T_8563; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8574 = _T_4925 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8575 = _GEN_796 == 7'h73; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8577 = _T_8575 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8579 = _T_8577 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8580 = _T_8574 | _T_8579; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8590 = _T_4929 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8591 = _GEN_796 == 7'h74; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8593 = _T_8591 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8595 = _T_8593 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8596 = _T_8590 | _T_8595; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8606 = _T_4933 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8607 = _GEN_796 == 7'h75; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8609 = _T_8607 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8611 = _T_8609 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8612 = _T_8606 | _T_8611; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8622 = _T_4937 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8623 = _GEN_796 == 7'h76; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8625 = _T_8623 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8627 = _T_8625 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8628 = _T_8622 | _T_8627; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8638 = _T_4941 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8639 = _GEN_796 == 7'h77; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8641 = _T_8639 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8643 = _T_8641 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8644 = _T_8638 | _T_8643; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8654 = _T_4945 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8655 = _GEN_796 == 7'h78; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8657 = _T_8655 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8659 = _T_8657 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8660 = _T_8654 | _T_8659; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8670 = _T_4949 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8671 = _GEN_796 == 7'h79; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8673 = _T_8671 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8675 = _T_8673 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8676 = _T_8670 | _T_8675; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8686 = _T_4953 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8687 = _GEN_796 == 7'h7a; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8689 = _T_8687 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8691 = _T_8689 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8692 = _T_8686 | _T_8691; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8702 = _T_4957 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8703 = _GEN_796 == 7'h7b; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8705 = _T_8703 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8707 = _T_8705 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8708 = _T_8702 | _T_8707; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8718 = _T_4961 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8719 = _GEN_796 == 7'h7c; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8721 = _T_8719 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8723 = _T_8721 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8724 = _T_8718 | _T_8723; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8734 = _T_4965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8735 = _GEN_796 == 7'h7d; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8737 = _T_8735 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8739 = _T_8737 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8740 = _T_8734 | _T_8739; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8750 = _T_4969 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8751 = _GEN_796 == 7'h7e; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8753 = _T_8751 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8755 = _T_8753 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8756 = _T_8750 | _T_8755; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8766 = _T_4973 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8767 = _GEN_796 == 7'h7f; // @[el2_ifu_mem_ctl.scala 736:101]
  wire  _T_8769 = _T_8767 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8771 = _T_8769 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8772 = _T_8766 | _T_8771; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8782 = _T_4849 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8785 = _T_8271 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8787 = _T_8785 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8788 = _T_8782 | _T_8787; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8798 = _T_4853 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8801 = _T_8287 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8803 = _T_8801 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8804 = _T_8798 | _T_8803; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8814 = _T_4857 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8817 = _T_8303 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8819 = _T_8817 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8820 = _T_8814 | _T_8819; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8830 = _T_4861 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8833 = _T_8319 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8835 = _T_8833 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8836 = _T_8830 | _T_8835; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8846 = _T_4865 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8849 = _T_8335 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8851 = _T_8849 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8852 = _T_8846 | _T_8851; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8862 = _T_4869 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8865 = _T_8351 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8867 = _T_8865 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8868 = _T_8862 | _T_8867; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8878 = _T_4873 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8881 = _T_8367 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8883 = _T_8881 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8884 = _T_8878 | _T_8883; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8894 = _T_4877 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8897 = _T_8383 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8899 = _T_8897 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8900 = _T_8894 | _T_8899; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8910 = _T_4881 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8913 = _T_8399 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8915 = _T_8913 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8916 = _T_8910 | _T_8915; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8926 = _T_4885 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8929 = _T_8415 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8931 = _T_8929 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8932 = _T_8926 | _T_8931; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8942 = _T_4889 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8945 = _T_8431 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8947 = _T_8945 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8948 = _T_8942 | _T_8947; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8958 = _T_4893 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8961 = _T_8447 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8963 = _T_8961 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8964 = _T_8958 | _T_8963; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8974 = _T_4897 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8977 = _T_8463 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8979 = _T_8977 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8980 = _T_8974 | _T_8979; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_8990 = _T_4901 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_8993 = _T_8479 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_8995 = _T_8993 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_8996 = _T_8990 | _T_8995; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9006 = _T_4905 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9009 = _T_8495 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9011 = _T_9009 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9012 = _T_9006 | _T_9011; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9022 = _T_4909 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9025 = _T_8511 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9027 = _T_9025 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9028 = _T_9022 | _T_9027; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9038 = _T_4913 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9041 = _T_8527 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9043 = _T_9041 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9044 = _T_9038 | _T_9043; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9054 = _T_4917 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9057 = _T_8543 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9059 = _T_9057 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9060 = _T_9054 | _T_9059; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9070 = _T_4921 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9073 = _T_8559 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9075 = _T_9073 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9076 = _T_9070 | _T_9075; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9086 = _T_4925 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9089 = _T_8575 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9091 = _T_9089 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9092 = _T_9086 | _T_9091; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9102 = _T_4929 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9105 = _T_8591 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9107 = _T_9105 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9108 = _T_9102 | _T_9107; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9118 = _T_4933 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9121 = _T_8607 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9123 = _T_9121 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9124 = _T_9118 | _T_9123; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9134 = _T_4937 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9137 = _T_8623 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9139 = _T_9137 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9140 = _T_9134 | _T_9139; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9150 = _T_4941 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9153 = _T_8639 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9155 = _T_9153 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9156 = _T_9150 | _T_9155; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9166 = _T_4945 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9169 = _T_8655 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9171 = _T_9169 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9172 = _T_9166 | _T_9171; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9182 = _T_4949 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9185 = _T_8671 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9187 = _T_9185 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9188 = _T_9182 | _T_9187; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9198 = _T_4953 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9201 = _T_8687 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9203 = _T_9201 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9204 = _T_9198 | _T_9203; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9214 = _T_4957 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9217 = _T_8703 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9219 = _T_9217 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9220 = _T_9214 | _T_9219; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9230 = _T_4961 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9233 = _T_8719 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9235 = _T_9233 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9236 = _T_9230 | _T_9235; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9246 = _T_4965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9249 = _T_8735 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9251 = _T_9249 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9252 = _T_9246 | _T_9251; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9262 = _T_4969 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9265 = _T_8751 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9267 = _T_9265 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9268 = _T_9262 | _T_9267; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_9278 = _T_4973 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:58]
  wire  _T_9281 = _T_8767 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 736:123]
  wire  _T_9283 = _T_9281 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 736:144]
  wire  _T_9284 = _T_9278 | _T_9283; // @[el2_ifu_mem_ctl.scala 736:80]
  wire  _T_10085 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 790:63]
  wire  _T_10086 = _T_10085 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 790:85]
  wire [1:0] _T_10088 = _T_10086 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10095; // @[el2_ifu_mem_ctl.scala 795:58]
  reg  _T_10096; // @[el2_ifu_mem_ctl.scala 796:58]
  reg  _T_10097; // @[el2_ifu_mem_ctl.scala 797:59]
  wire  _T_10098 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 798:78]
  wire  _T_10099 = ifu_bus_arvalid_ff & _T_10098; // @[el2_ifu_mem_ctl.scala 798:76]
  wire  _T_10100 = _T_10099 & miss_pending; // @[el2_ifu_mem_ctl.scala 798:98]
  reg  _T_10101; // @[el2_ifu_mem_ctl.scala 798:56]
  reg  _T_10102; // @[el2_ifu_mem_ctl.scala 799:57]
  wire  _T_10105 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 804:71]
  wire  _T_10107 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 804:124]
  wire  _T_10109 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 805:50]
  wire  _T_10111 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 805:103]
  wire [3:0] _T_10114 = {_T_10105,_T_10107,_T_10109,_T_10111}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 807:53]
  reg  _T_10125; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 319:26]
  assign io_ifu_ic_mb_empty = _T_317 | _T_222; // @[el2_ifu_mem_ctl.scala 318:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 185:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3920; // @[el2_ifu_mem_ctl.scala 686:21]
  assign io_ifu_pmu_ic_miss = _T_10102; // @[el2_ifu_mem_ctl.scala 799:22]
  assign io_ifu_pmu_ic_hit = _T_10101; // @[el2_ifu_mem_ctl.scala 798:21]
  assign io_ifu_pmu_bus_error = _T_10097; // @[el2_ifu_mem_ctl.scala 797:24]
  assign io_ifu_pmu_bus_busy = _T_10096; // @[el2_ifu_mem_ctl.scala 796:23]
  assign io_ifu_pmu_bus_trxn = _T_10095; // @[el2_ifu_mem_ctl.scala 795:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 136:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 135:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 130:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 134:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 132:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 143:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 145:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 138:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 131:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 129:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 127:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 128:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 146:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 141:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 548:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2514; // @[el2_ifu_mem_ctl.scala 549:19]
  assign io_ifu_axi_araddr = _T_2516 & _T_2518; // @[el2_ifu_mem_ctl.scala 550:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 553:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 142:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 551:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 554:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 552:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 144:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 139:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 555:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 645:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 643:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 647:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 638:20]
  assign io_iccm_ready = _T_2617 & _T_2611; // @[el2_ifu_mem_ctl.scala 618:17]
  assign io_ic_rw_addr = _T_331 | _T_332; // @[el2_ifu_mem_ctl.scala 328:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 685:15]
  assign io_ic_rd_en = _T_3898 | _T_3903; // @[el2_ifu_mem_ctl.scala 676:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 335:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 335:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 336:23]
  assign io_ifu_ic_debug_rd_data = _T_1202; // @[el2_ifu_mem_ctl.scala 344:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 800:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 802:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 803:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 801:25]
  assign io_ic_debug_way = _T_10114[1:0]; // @[el2_ifu_mem_ctl.scala 804:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10088; // @[el2_ifu_mem_ctl.scala 790:19]
  assign io_iccm_rw_addr = _T_3052[14:0]; // @[el2_ifu_mem_ctl.scala 649:19]
  assign io_iccm_wren = _T_2621 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 620:16]
  assign io_iccm_rden = _T_2625 | _T_2626; // @[el2_ifu_mem_ctl.scala 621:16]
  assign io_iccm_wr_data = _T_3027 ? _T_3028 : _T_3035; // @[el2_ifu_mem_ctl.scala 626:19]
  assign io_iccm_wr_size = _T_2631 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 623:19]
  assign io_ic_hit_f = _T_254 | _T_255; // @[el2_ifu_mem_ctl.scala 280:15]
  assign io_ic_access_fault_f = _T_2401 & _T_308; // @[el2_ifu_mem_ctl.scala 375:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1266; // @[el2_ifu_mem_ctl.scala 376:29]
  assign io_iccm_rd_ecc_single_err = _T_3843 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 662:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 663:29]
  assign io_ic_error_start = _T_1190 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 338:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 184:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 183:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 380:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 372:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 369:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 370:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10125; // @[el2_ifu_mem_ctl.scala 811:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2406; // @[el2_ifu_mem_ctl.scala 468:27]
  assign io_iccm_correction_state = _T_2434 ? 1'h0 : _GEN_59; // @[el2_ifu_mem_ctl.scala 503:28 el2_ifu_mem_ctl.scala 516:32 el2_ifu_mem_ctl.scala 523:32 el2_ifu_mem_ctl.scala 530:32]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_3[30:0];
  _RAND_4 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  perr_state = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  err_stop_state = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reset_all_tags = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  imb_ff = _RAND_16[30:0];
  _RAND_17 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_5108 = _RAND_19[6:0];
  _RAND_20 = {1{`RANDOM}};
  _T_4464 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4460 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_4456 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_4452 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_4448 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_4444 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_4440 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_4436 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_4432 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_4428 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_4424 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_4420 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_4416 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_4412 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_4408 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_4404 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_4400 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_4396 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_4392 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_4388 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_4384 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_4380 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_4376 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_4372 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_4368 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_4364 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_4360 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_4356 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_4352 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_4348 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_4344 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_4340 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_4336 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_4332 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_4328 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_4324 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_4320 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_4316 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_4312 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_4308 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_4304 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_4300 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_4296 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_4292 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_4288 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_4284 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_4280 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_4276 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_4272 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_4268 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_4264 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_4260 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_4256 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_4252 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_4248 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_4244 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_4240 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_4236 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_4232 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_4228 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_4224 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_4220 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_4216 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_4212 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_4208 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_4204 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_4200 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_4196 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_4192 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_4188 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_4184 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_4180 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_4176 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_4172 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_4168 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_4164 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_4160 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_4156 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_4152 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_4148 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_4144 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_4140 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_4136 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_4132 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_4128 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_4124 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_4120 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_4116 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_4112 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_4108 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_4104 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_4100 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_4096 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_4092 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_4088 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_4084 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_4080 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_4076 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_4072 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_4068 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_4064 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_4060 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_4056 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_4052 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_4048 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_4044 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_4040 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_4036 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_4032 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_4028 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_4024 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_4020 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_4016 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_4012 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_4008 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_4004 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_4000 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3996 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3992 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3988 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3984 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3980 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3976 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3972 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3968 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3964 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3960 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3956 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_148[30:0];
  _RAND_149 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  reset_ic_ff = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  miss_addr = _RAND_155[25:0];
  _RAND_156 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_157[2:0];
  _RAND_158 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_158[0:0];
  _RAND_159 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_159[63:0];
  _RAND_160 = {2{`RANDOM}};
  _T_1286 = _RAND_160[63:0];
  _RAND_161 = {2{`RANDOM}};
  _T_1288 = _RAND_161[63:0];
  _RAND_162 = {2{`RANDOM}};
  _T_1290 = _RAND_162[63:0];
  _RAND_163 = {2{`RANDOM}};
  _T_1292 = _RAND_163[63:0];
  _RAND_164 = {2{`RANDOM}};
  _T_1294 = _RAND_164[63:0];
  _RAND_165 = {2{`RANDOM}};
  _T_1296 = _RAND_165[63:0];
  _RAND_166 = {2{`RANDOM}};
  _T_1298 = _RAND_166[63:0];
  _RAND_167 = {2{`RANDOM}};
  _T_1300 = _RAND_167[63:0];
  _RAND_168 = {2{`RANDOM}};
  _T_1302 = _RAND_168[63:0];
  _RAND_169 = {2{`RANDOM}};
  _T_1304 = _RAND_169[63:0];
  _RAND_170 = {2{`RANDOM}};
  _T_1306 = _RAND_170[63:0];
  _RAND_171 = {2{`RANDOM}};
  _T_1308 = _RAND_171[63:0];
  _RAND_172 = {2{`RANDOM}};
  _T_1310 = _RAND_172[63:0];
  _RAND_173 = {2{`RANDOM}};
  _T_1312 = _RAND_173[63:0];
  _RAND_174 = {2{`RANDOM}};
  _T_1314 = _RAND_174[63:0];
  _RAND_175 = {2{`RANDOM}};
  _T_1316 = _RAND_175[63:0];
  _RAND_176 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_176[0:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_179[0:0];
  _RAND_180 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_435[1:0];
  _RAND_436 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_436[0:0];
  _RAND_437 = {3{`RANDOM}};
  _T_1202 = _RAND_437[70:0];
  _RAND_438 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_438[5:0];
  _RAND_439 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_440[0:0];
  _RAND_441 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_441[2:0];
  _RAND_442 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_442[0:0];
  _RAND_443 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_444[0:0];
  _RAND_445 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_445[38:0];
  _RAND_446 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_446[1:0];
  _RAND_447 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_447[2:0];
  _RAND_448 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_448[2:0];
  _RAND_449 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_449[0:0];
  _RAND_450 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_450[63:0];
  _RAND_451 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_451[13:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_452[0:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_453[13:0];
  _RAND_454 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_454[6:0];
  _RAND_455 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_455[0:0];
  _RAND_456 = {1{`RANDOM}};
  way_status_new_ff = _RAND_456[2:0];
  _RAND_457 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_457[1:0];
  _RAND_458 = {1{`RANDOM}};
  ic_valid_ff = _RAND_458[0:0];
  _RAND_459 = {1{`RANDOM}};
  _T_10095 = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  _T_10096 = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  _T_10097 = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  _T_10101 = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_10102 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10125 = _RAND_464[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_25) begin
        if (_T_27) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_32) begin
        if (_T_37) begin
          miss_state <= 3'h0;
        end else if (_T_41) begin
          miss_state <= 3'h3;
        end else if (_T_48) begin
          miss_state <= 3'h1;
        end else if (_T_52) begin
          miss_state <= 3'h0;
        end else if (_T_63) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h0;
        end else if (_T_76) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_93) begin
        miss_state <= 3'h0;
      end else if (_T_97) begin
        if (_T_104) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_112) begin
        if (_T_117) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_123) begin
        if (_T_128) begin
          miss_state <= 3'h5;
        end else if (_T_134) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_142) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_33) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_33) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      _T_4464 <= 3'h0;
    end else if (_T_4463) begin
      _T_4464 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4460 <= 3'h0;
    end else if (_T_4459) begin
      _T_4460 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4456 <= 3'h0;
    end else if (_T_4455) begin
      _T_4456 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4452 <= 3'h0;
    end else if (_T_4451) begin
      _T_4452 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4448 <= 3'h0;
    end else if (_T_4447) begin
      _T_4448 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4444 <= 3'h0;
    end else if (_T_4443) begin
      _T_4444 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4440 <= 3'h0;
    end else if (_T_4439) begin
      _T_4440 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4436 <= 3'h0;
    end else if (_T_4435) begin
      _T_4436 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4432 <= 3'h0;
    end else if (_T_4431) begin
      _T_4432 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4428 <= 3'h0;
    end else if (_T_4427) begin
      _T_4428 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4424 <= 3'h0;
    end else if (_T_4423) begin
      _T_4424 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4420 <= 3'h0;
    end else if (_T_4419) begin
      _T_4420 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4416 <= 3'h0;
    end else if (_T_4415) begin
      _T_4416 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4412 <= 3'h0;
    end else if (_T_4411) begin
      _T_4412 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4408 <= 3'h0;
    end else if (_T_4407) begin
      _T_4408 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4404 <= 3'h0;
    end else if (_T_4403) begin
      _T_4404 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4400 <= 3'h0;
    end else if (_T_4399) begin
      _T_4400 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4396 <= 3'h0;
    end else if (_T_4395) begin
      _T_4396 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4392 <= 3'h0;
    end else if (_T_4391) begin
      _T_4392 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4388 <= 3'h0;
    end else if (_T_4387) begin
      _T_4388 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4384 <= 3'h0;
    end else if (_T_4383) begin
      _T_4384 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4380 <= 3'h0;
    end else if (_T_4379) begin
      _T_4380 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4376 <= 3'h0;
    end else if (_T_4375) begin
      _T_4376 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4372 <= 3'h0;
    end else if (_T_4371) begin
      _T_4372 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4368 <= 3'h0;
    end else if (_T_4367) begin
      _T_4368 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4364 <= 3'h0;
    end else if (_T_4363) begin
      _T_4364 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4360 <= 3'h0;
    end else if (_T_4359) begin
      _T_4360 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4356 <= 3'h0;
    end else if (_T_4355) begin
      _T_4356 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4352 <= 3'h0;
    end else if (_T_4351) begin
      _T_4352 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4348 <= 3'h0;
    end else if (_T_4347) begin
      _T_4348 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4344 <= 3'h0;
    end else if (_T_4343) begin
      _T_4344 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4340 <= 3'h0;
    end else if (_T_4339) begin
      _T_4340 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4336 <= 3'h0;
    end else if (_T_4335) begin
      _T_4336 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4332 <= 3'h0;
    end else if (_T_4331) begin
      _T_4332 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4328 <= 3'h0;
    end else if (_T_4327) begin
      _T_4328 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4324 <= 3'h0;
    end else if (_T_4323) begin
      _T_4324 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4320 <= 3'h0;
    end else if (_T_4319) begin
      _T_4320 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4316 <= 3'h0;
    end else if (_T_4315) begin
      _T_4316 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4312 <= 3'h0;
    end else if (_T_4311) begin
      _T_4312 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4308 <= 3'h0;
    end else if (_T_4307) begin
      _T_4308 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4304 <= 3'h0;
    end else if (_T_4303) begin
      _T_4304 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4300 <= 3'h0;
    end else if (_T_4299) begin
      _T_4300 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4296 <= 3'h0;
    end else if (_T_4295) begin
      _T_4296 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4292 <= 3'h0;
    end else if (_T_4291) begin
      _T_4292 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4288 <= 3'h0;
    end else if (_T_4287) begin
      _T_4288 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4284 <= 3'h0;
    end else if (_T_4283) begin
      _T_4284 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4280 <= 3'h0;
    end else if (_T_4279) begin
      _T_4280 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4276 <= 3'h0;
    end else if (_T_4275) begin
      _T_4276 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4272 <= 3'h0;
    end else if (_T_4271) begin
      _T_4272 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4268 <= 3'h0;
    end else if (_T_4267) begin
      _T_4268 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4264 <= 3'h0;
    end else if (_T_4263) begin
      _T_4264 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4260 <= 3'h0;
    end else if (_T_4259) begin
      _T_4260 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4256 <= 3'h0;
    end else if (_T_4255) begin
      _T_4256 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4252 <= 3'h0;
    end else if (_T_4251) begin
      _T_4252 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4248 <= 3'h0;
    end else if (_T_4247) begin
      _T_4248 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4244 <= 3'h0;
    end else if (_T_4243) begin
      _T_4244 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4240 <= 3'h0;
    end else if (_T_4239) begin
      _T_4240 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4236 <= 3'h0;
    end else if (_T_4235) begin
      _T_4236 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4232 <= 3'h0;
    end else if (_T_4231) begin
      _T_4232 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4228 <= 3'h0;
    end else if (_T_4227) begin
      _T_4228 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4224 <= 3'h0;
    end else if (_T_4223) begin
      _T_4224 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4220 <= 3'h0;
    end else if (_T_4219) begin
      _T_4220 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4216 <= 3'h0;
    end else if (_T_4215) begin
      _T_4216 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4212 <= 3'h0;
    end else if (_T_4211) begin
      _T_4212 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4208 <= 3'h0;
    end else if (_T_4207) begin
      _T_4208 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4204 <= 3'h0;
    end else if (_T_4203) begin
      _T_4204 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4200 <= 3'h0;
    end else if (_T_4199) begin
      _T_4200 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4196 <= 3'h0;
    end else if (_T_4195) begin
      _T_4196 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4192 <= 3'h0;
    end else if (_T_4191) begin
      _T_4192 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4188 <= 3'h0;
    end else if (_T_4187) begin
      _T_4188 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4184 <= 3'h0;
    end else if (_T_4183) begin
      _T_4184 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4180 <= 3'h0;
    end else if (_T_4179) begin
      _T_4180 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4176 <= 3'h0;
    end else if (_T_4175) begin
      _T_4176 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4172 <= 3'h0;
    end else if (_T_4171) begin
      _T_4172 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4168 <= 3'h0;
    end else if (_T_4167) begin
      _T_4168 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4164 <= 3'h0;
    end else if (_T_4163) begin
      _T_4164 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4160 <= 3'h0;
    end else if (_T_4159) begin
      _T_4160 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4156 <= 3'h0;
    end else if (_T_4155) begin
      _T_4156 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4152 <= 3'h0;
    end else if (_T_4151) begin
      _T_4152 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4148 <= 3'h0;
    end else if (_T_4147) begin
      _T_4148 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4144 <= 3'h0;
    end else if (_T_4143) begin
      _T_4144 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4140 <= 3'h0;
    end else if (_T_4139) begin
      _T_4140 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4136 <= 3'h0;
    end else if (_T_4135) begin
      _T_4136 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4132 <= 3'h0;
    end else if (_T_4131) begin
      _T_4132 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4128 <= 3'h0;
    end else if (_T_4127) begin
      _T_4128 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4124 <= 3'h0;
    end else if (_T_4123) begin
      _T_4124 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4120 <= 3'h0;
    end else if (_T_4119) begin
      _T_4120 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4116 <= 3'h0;
    end else if (_T_4115) begin
      _T_4116 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4112 <= 3'h0;
    end else if (_T_4111) begin
      _T_4112 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4108 <= 3'h0;
    end else if (_T_4107) begin
      _T_4108 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4104 <= 3'h0;
    end else if (_T_4103) begin
      _T_4104 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4100 <= 3'h0;
    end else if (_T_4099) begin
      _T_4100 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4096 <= 3'h0;
    end else if (_T_4095) begin
      _T_4096 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4092 <= 3'h0;
    end else if (_T_4091) begin
      _T_4092 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4088 <= 3'h0;
    end else if (_T_4087) begin
      _T_4088 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4084 <= 3'h0;
    end else if (_T_4083) begin
      _T_4084 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4080 <= 3'h0;
    end else if (_T_4079) begin
      _T_4080 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4076 <= 3'h0;
    end else if (_T_4075) begin
      _T_4076 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4072 <= 3'h0;
    end else if (_T_4071) begin
      _T_4072 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4068 <= 3'h0;
    end else if (_T_4067) begin
      _T_4068 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4064 <= 3'h0;
    end else if (_T_4063) begin
      _T_4064 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4060 <= 3'h0;
    end else if (_T_4059) begin
      _T_4060 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4056 <= 3'h0;
    end else if (_T_4055) begin
      _T_4056 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4052 <= 3'h0;
    end else if (_T_4051) begin
      _T_4052 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4048 <= 3'h0;
    end else if (_T_4047) begin
      _T_4048 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4044 <= 3'h0;
    end else if (_T_4043) begin
      _T_4044 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4040 <= 3'h0;
    end else if (_T_4039) begin
      _T_4040 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4036 <= 3'h0;
    end else if (_T_4035) begin
      _T_4036 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4032 <= 3'h0;
    end else if (_T_4031) begin
      _T_4032 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4028 <= 3'h0;
    end else if (_T_4027) begin
      _T_4028 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4024 <= 3'h0;
    end else if (_T_4023) begin
      _T_4024 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4020 <= 3'h0;
    end else if (_T_4019) begin
      _T_4020 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4016 <= 3'h0;
    end else if (_T_4015) begin
      _T_4016 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4012 <= 3'h0;
    end else if (_T_4011) begin
      _T_4012 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4008 <= 3'h0;
    end else if (_T_4007) begin
      _T_4008 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4004 <= 3'h0;
    end else if (_T_4003) begin
      _T_4004 <= way_status_new_ff;
    end
    if (reset) begin
      _T_4000 <= 3'h0;
    end else if (_T_3999) begin
      _T_4000 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3996 <= 3'h0;
    end else if (_T_3995) begin
      _T_3996 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3992 <= 3'h0;
    end else if (_T_3991) begin
      _T_3992 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3988 <= 3'h0;
    end else if (_T_3987) begin
      _T_3988 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3984 <= 3'h0;
    end else if (_T_3983) begin
      _T_3984 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3980 <= 3'h0;
    end else if (_T_3979) begin
      _T_3980 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3976 <= 3'h0;
    end else if (_T_3975) begin
      _T_3976 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3972 <= 3'h0;
    end else if (_T_3971) begin
      _T_3972 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3968 <= 3'h0;
    end else if (_T_3967) begin
      _T_3968 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3964 <= 3'h0;
    end else if (_T_3963) begin
      _T_3964 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3960 <= 3'h0;
    end else if (_T_3959) begin
      _T_3960 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3956 <= 3'h0;
    end else if (_T_3955) begin
      _T_3956 <= way_status_new_ff;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    reset_ic_ff <= _T_289 & _T_290;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_222) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2557) begin
      if (_T_222) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2553;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1286 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1286 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1288 <= 64'h0;
    end else if (write_fill_data_0) begin
      _T_1288 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1290 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1290 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1292 <= 64'h0;
    end else if (write_fill_data_1) begin
      _T_1292 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1294 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1294 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1296 <= 64'h0;
    end else if (write_fill_data_2) begin
      _T_1296 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1298 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1298 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1300 <= 64'h0;
    end else if (write_fill_data_3) begin
      _T_1300 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1302 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1302 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1304 <= 64'h0;
    end else if (write_fill_data_4) begin
      _T_1304 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1306 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1306 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1308 <= 64'h0;
    end else if (write_fill_data_5) begin
      _T_1308 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1310 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1310 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1312 <= 64'h0;
    end else if (write_fill_data_6) begin
      _T_1312 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1314 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1314 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      _T_1316 <= 64'h0;
    end else if (write_fill_data_7) begin
      _T_1316 <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5716) begin
      ic_tag_valid_out_1_0 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5732) begin
      ic_tag_valid_out_1_1 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_5748) begin
      ic_tag_valid_out_1_2 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_5764) begin
      ic_tag_valid_out_1_3 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_5780) begin
      ic_tag_valid_out_1_4 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5796) begin
      ic_tag_valid_out_1_5 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5812) begin
      ic_tag_valid_out_1_6 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5828) begin
      ic_tag_valid_out_1_7 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5844) begin
      ic_tag_valid_out_1_8 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5860) begin
      ic_tag_valid_out_1_9 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5876) begin
      ic_tag_valid_out_1_10 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5892) begin
      ic_tag_valid_out_1_11 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5908) begin
      ic_tag_valid_out_1_12 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5924) begin
      ic_tag_valid_out_1_13 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5940) begin
      ic_tag_valid_out_1_14 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5956) begin
      ic_tag_valid_out_1_15 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5972) begin
      ic_tag_valid_out_1_16 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5988) begin
      ic_tag_valid_out_1_17 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6004) begin
      ic_tag_valid_out_1_18 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6020) begin
      ic_tag_valid_out_1_19 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6036) begin
      ic_tag_valid_out_1_20 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6052) begin
      ic_tag_valid_out_1_21 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6068) begin
      ic_tag_valid_out_1_22 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6084) begin
      ic_tag_valid_out_1_23 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6100) begin
      ic_tag_valid_out_1_24 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6116) begin
      ic_tag_valid_out_1_25 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6132) begin
      ic_tag_valid_out_1_26 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6148) begin
      ic_tag_valid_out_1_27 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6164) begin
      ic_tag_valid_out_1_28 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6180) begin
      ic_tag_valid_out_1_29 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6196) begin
      ic_tag_valid_out_1_30 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6212) begin
      ic_tag_valid_out_1_31 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_6740) begin
      ic_tag_valid_out_1_32 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_6756) begin
      ic_tag_valid_out_1_33 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_6772) begin
      ic_tag_valid_out_1_34 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6788) begin
      ic_tag_valid_out_1_35 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6804) begin
      ic_tag_valid_out_1_36 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6820) begin
      ic_tag_valid_out_1_37 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6836) begin
      ic_tag_valid_out_1_38 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6852) begin
      ic_tag_valid_out_1_39 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6868) begin
      ic_tag_valid_out_1_40 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6884) begin
      ic_tag_valid_out_1_41 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6900) begin
      ic_tag_valid_out_1_42 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6916) begin
      ic_tag_valid_out_1_43 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6932) begin
      ic_tag_valid_out_1_44 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6948) begin
      ic_tag_valid_out_1_45 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6964) begin
      ic_tag_valid_out_1_46 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6980) begin
      ic_tag_valid_out_1_47 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6996) begin
      ic_tag_valid_out_1_48 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7012) begin
      ic_tag_valid_out_1_49 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7028) begin
      ic_tag_valid_out_1_50 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7044) begin
      ic_tag_valid_out_1_51 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7060) begin
      ic_tag_valid_out_1_52 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7076) begin
      ic_tag_valid_out_1_53 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7092) begin
      ic_tag_valid_out_1_54 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7108) begin
      ic_tag_valid_out_1_55 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7124) begin
      ic_tag_valid_out_1_56 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7140) begin
      ic_tag_valid_out_1_57 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7156) begin
      ic_tag_valid_out_1_58 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7172) begin
      ic_tag_valid_out_1_59 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7188) begin
      ic_tag_valid_out_1_60 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7204) begin
      ic_tag_valid_out_1_61 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7220) begin
      ic_tag_valid_out_1_62 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7236) begin
      ic_tag_valid_out_1_63 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_7764) begin
      ic_tag_valid_out_1_64 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_7780) begin
      ic_tag_valid_out_1_65 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7796) begin
      ic_tag_valid_out_1_66 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7812) begin
      ic_tag_valid_out_1_67 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7828) begin
      ic_tag_valid_out_1_68 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7844) begin
      ic_tag_valid_out_1_69 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7860) begin
      ic_tag_valid_out_1_70 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7876) begin
      ic_tag_valid_out_1_71 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7892) begin
      ic_tag_valid_out_1_72 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7908) begin
      ic_tag_valid_out_1_73 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7924) begin
      ic_tag_valid_out_1_74 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7940) begin
      ic_tag_valid_out_1_75 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7956) begin
      ic_tag_valid_out_1_76 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7972) begin
      ic_tag_valid_out_1_77 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7988) begin
      ic_tag_valid_out_1_78 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8004) begin
      ic_tag_valid_out_1_79 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8020) begin
      ic_tag_valid_out_1_80 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8036) begin
      ic_tag_valid_out_1_81 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8052) begin
      ic_tag_valid_out_1_82 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8068) begin
      ic_tag_valid_out_1_83 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8084) begin
      ic_tag_valid_out_1_84 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8100) begin
      ic_tag_valid_out_1_85 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8116) begin
      ic_tag_valid_out_1_86 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8132) begin
      ic_tag_valid_out_1_87 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8148) begin
      ic_tag_valid_out_1_88 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8164) begin
      ic_tag_valid_out_1_89 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8180) begin
      ic_tag_valid_out_1_90 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8196) begin
      ic_tag_valid_out_1_91 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8212) begin
      ic_tag_valid_out_1_92 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8228) begin
      ic_tag_valid_out_1_93 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8244) begin
      ic_tag_valid_out_1_94 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8260) begin
      ic_tag_valid_out_1_95 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8788) begin
      ic_tag_valid_out_1_96 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8804) begin
      ic_tag_valid_out_1_97 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8820) begin
      ic_tag_valid_out_1_98 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8836) begin
      ic_tag_valid_out_1_99 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8852) begin
      ic_tag_valid_out_1_100 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8868) begin
      ic_tag_valid_out_1_101 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8884) begin
      ic_tag_valid_out_1_102 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8900) begin
      ic_tag_valid_out_1_103 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8916) begin
      ic_tag_valid_out_1_104 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8932) begin
      ic_tag_valid_out_1_105 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8948) begin
      ic_tag_valid_out_1_106 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8964) begin
      ic_tag_valid_out_1_107 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8980) begin
      ic_tag_valid_out_1_108 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8996) begin
      ic_tag_valid_out_1_109 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9012) begin
      ic_tag_valid_out_1_110 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9028) begin
      ic_tag_valid_out_1_111 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9044) begin
      ic_tag_valid_out_1_112 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9060) begin
      ic_tag_valid_out_1_113 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9076) begin
      ic_tag_valid_out_1_114 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9092) begin
      ic_tag_valid_out_1_115 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9108) begin
      ic_tag_valid_out_1_116 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9124) begin
      ic_tag_valid_out_1_117 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9140) begin
      ic_tag_valid_out_1_118 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9156) begin
      ic_tag_valid_out_1_119 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9172) begin
      ic_tag_valid_out_1_120 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9188) begin
      ic_tag_valid_out_1_121 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9204) begin
      ic_tag_valid_out_1_122 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9220) begin
      ic_tag_valid_out_1_123 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9236) begin
      ic_tag_valid_out_1_124 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9252) begin
      ic_tag_valid_out_1_125 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9268) begin
      ic_tag_valid_out_1_126 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9284) begin
      ic_tag_valid_out_1_127 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5204) begin
      ic_tag_valid_out_0_0 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5220) begin
      ic_tag_valid_out_0_1 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5236) begin
      ic_tag_valid_out_0_2 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5252) begin
      ic_tag_valid_out_0_3 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5268) begin
      ic_tag_valid_out_0_4 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5284) begin
      ic_tag_valid_out_0_5 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5300) begin
      ic_tag_valid_out_0_6 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5316) begin
      ic_tag_valid_out_0_7 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5332) begin
      ic_tag_valid_out_0_8 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5348) begin
      ic_tag_valid_out_0_9 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5364) begin
      ic_tag_valid_out_0_10 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5380) begin
      ic_tag_valid_out_0_11 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5396) begin
      ic_tag_valid_out_0_12 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5412) begin
      ic_tag_valid_out_0_13 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5428) begin
      ic_tag_valid_out_0_14 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5444) begin
      ic_tag_valid_out_0_15 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5460) begin
      ic_tag_valid_out_0_16 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5476) begin
      ic_tag_valid_out_0_17 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5492) begin
      ic_tag_valid_out_0_18 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5508) begin
      ic_tag_valid_out_0_19 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5524) begin
      ic_tag_valid_out_0_20 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5540) begin
      ic_tag_valid_out_0_21 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5556) begin
      ic_tag_valid_out_0_22 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5572) begin
      ic_tag_valid_out_0_23 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5588) begin
      ic_tag_valid_out_0_24 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5604) begin
      ic_tag_valid_out_0_25 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5620) begin
      ic_tag_valid_out_0_26 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5636) begin
      ic_tag_valid_out_0_27 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5652) begin
      ic_tag_valid_out_0_28 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5668) begin
      ic_tag_valid_out_0_29 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5684) begin
      ic_tag_valid_out_0_30 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5700) begin
      ic_tag_valid_out_0_31 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6228) begin
      ic_tag_valid_out_0_32 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6244) begin
      ic_tag_valid_out_0_33 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6260) begin
      ic_tag_valid_out_0_34 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6276) begin
      ic_tag_valid_out_0_35 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6292) begin
      ic_tag_valid_out_0_36 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6308) begin
      ic_tag_valid_out_0_37 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6324) begin
      ic_tag_valid_out_0_38 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6340) begin
      ic_tag_valid_out_0_39 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6356) begin
      ic_tag_valid_out_0_40 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6372) begin
      ic_tag_valid_out_0_41 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6388) begin
      ic_tag_valid_out_0_42 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6404) begin
      ic_tag_valid_out_0_43 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6420) begin
      ic_tag_valid_out_0_44 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6436) begin
      ic_tag_valid_out_0_45 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6452) begin
      ic_tag_valid_out_0_46 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6468) begin
      ic_tag_valid_out_0_47 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6484) begin
      ic_tag_valid_out_0_48 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6500) begin
      ic_tag_valid_out_0_49 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6516) begin
      ic_tag_valid_out_0_50 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6532) begin
      ic_tag_valid_out_0_51 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6548) begin
      ic_tag_valid_out_0_52 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6564) begin
      ic_tag_valid_out_0_53 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6580) begin
      ic_tag_valid_out_0_54 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6596) begin
      ic_tag_valid_out_0_55 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6612) begin
      ic_tag_valid_out_0_56 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6628) begin
      ic_tag_valid_out_0_57 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6644) begin
      ic_tag_valid_out_0_58 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6660) begin
      ic_tag_valid_out_0_59 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6676) begin
      ic_tag_valid_out_0_60 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_6692) begin
      ic_tag_valid_out_0_61 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_6708) begin
      ic_tag_valid_out_0_62 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_6724) begin
      ic_tag_valid_out_0_63 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7252) begin
      ic_tag_valid_out_0_64 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7268) begin
      ic_tag_valid_out_0_65 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7284) begin
      ic_tag_valid_out_0_66 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7300) begin
      ic_tag_valid_out_0_67 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7316) begin
      ic_tag_valid_out_0_68 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7332) begin
      ic_tag_valid_out_0_69 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7348) begin
      ic_tag_valid_out_0_70 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7364) begin
      ic_tag_valid_out_0_71 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7380) begin
      ic_tag_valid_out_0_72 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7396) begin
      ic_tag_valid_out_0_73 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7412) begin
      ic_tag_valid_out_0_74 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7428) begin
      ic_tag_valid_out_0_75 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7444) begin
      ic_tag_valid_out_0_76 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7460) begin
      ic_tag_valid_out_0_77 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7476) begin
      ic_tag_valid_out_0_78 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7492) begin
      ic_tag_valid_out_0_79 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7508) begin
      ic_tag_valid_out_0_80 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7524) begin
      ic_tag_valid_out_0_81 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7540) begin
      ic_tag_valid_out_0_82 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7556) begin
      ic_tag_valid_out_0_83 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7572) begin
      ic_tag_valid_out_0_84 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7588) begin
      ic_tag_valid_out_0_85 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7604) begin
      ic_tag_valid_out_0_86 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_7620) begin
      ic_tag_valid_out_0_87 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_7636) begin
      ic_tag_valid_out_0_88 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_7652) begin
      ic_tag_valid_out_0_89 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_7668) begin
      ic_tag_valid_out_0_90 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_7684) begin
      ic_tag_valid_out_0_91 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_7700) begin
      ic_tag_valid_out_0_92 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_7716) begin
      ic_tag_valid_out_0_93 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_7732) begin
      ic_tag_valid_out_0_94 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_7748) begin
      ic_tag_valid_out_0_95 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8276) begin
      ic_tag_valid_out_0_96 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8292) begin
      ic_tag_valid_out_0_97 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8308) begin
      ic_tag_valid_out_0_98 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8324) begin
      ic_tag_valid_out_0_99 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8340) begin
      ic_tag_valid_out_0_100 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8356) begin
      ic_tag_valid_out_0_101 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8372) begin
      ic_tag_valid_out_0_102 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8388) begin
      ic_tag_valid_out_0_103 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8404) begin
      ic_tag_valid_out_0_104 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8420) begin
      ic_tag_valid_out_0_105 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8436) begin
      ic_tag_valid_out_0_106 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8452) begin
      ic_tag_valid_out_0_107 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8468) begin
      ic_tag_valid_out_0_108 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8484) begin
      ic_tag_valid_out_0_109 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8500) begin
      ic_tag_valid_out_0_110 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8516) begin
      ic_tag_valid_out_0_111 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8532) begin
      ic_tag_valid_out_0_112 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8548) begin
      ic_tag_valid_out_0_113 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_8564) begin
      ic_tag_valid_out_0_114 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_8580) begin
      ic_tag_valid_out_0_115 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_8596) begin
      ic_tag_valid_out_0_116 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_8612) begin
      ic_tag_valid_out_0_117 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_8628) begin
      ic_tag_valid_out_0_118 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_8644) begin
      ic_tag_valid_out_0_119 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_8660) begin
      ic_tag_valid_out_0_120 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_8676) begin
      ic_tag_valid_out_0_121 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_8692) begin
      ic_tag_valid_out_0_122 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_8708) begin
      ic_tag_valid_out_0_123 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_8724) begin
      ic_tag_valid_out_0_124 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_8740) begin
      ic_tag_valid_out_0_125 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_8756) begin
      ic_tag_valid_out_0_126 <= _T_5195;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_8772) begin
      ic_tag_valid_out_0_127 <= _T_5195;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1202 <= 71'h0;
    end else if (ic_debug_ict_array_sel_ff) begin
      _T_1202 <= {{5'd0}, _T_1201};
    end else begin
      _T_1202 <= io_ic_debug_rd_data;
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2506) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2581) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2625;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2409) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2411) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2421) begin
        perr_state <= 3'h0;
      end else if (_T_2424) begin
        if (_T_2426) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2430) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2434) begin
        err_stop_state <= 2'h1;
      end else if (_T_2439) begin
        if (_T_2441) begin
          err_stop_state <= 2'h0;
        end else if (_T_2462) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2466) begin
        if (_T_2441) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2483) begin
        if (_T_2487) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1347;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_5108 <= 7'h0;
    end else if (_T_3929) begin
      _T_5108 <= io_ic_debug_addr[9:3];
    end else begin
      _T_5108 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1387;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3864;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_3039;
    end else begin
      iccm_dma_rdata <= _T_3040;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3860;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3929) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3932) begin
      way_status_new_ff <= _T_3936;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3932) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10125 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10125 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10095 <= 1'h0;
    end else begin
      _T_10095 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10096 <= 1'h0;
    end else begin
      _T_10096 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10097 <= 1'h0;
    end else begin
      _T_10097 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10101 <= 1'h0;
    end else begin
      _T_10101 <= _T_10100;
    end
    if (reset) begin
      _T_10102 <= 1'h0;
    end else begin
      _T_10102 <= bus_cmd_sent;
    end
  end
endmodule
