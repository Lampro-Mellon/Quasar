module rvecc_encode_64(
  input  [63:0] io_din,
  output [6:0]  io_ecc_out
);
  wire  w0_0 = io_din[0]; // @[el2_lib.scala 343:39]
  wire  w0_1 = io_din[1]; // @[el2_lib.scala 343:39]
  wire  w1_1 = io_din[2]; // @[el2_lib.scala 344:39]
  wire  w0_2 = io_din[3]; // @[el2_lib.scala 343:39]
  wire  w0_3 = io_din[4]; // @[el2_lib.scala 343:39]
  wire  w1_3 = io_din[5]; // @[el2_lib.scala 344:39]
  wire  w0_4 = io_din[6]; // @[el2_lib.scala 343:39]
  wire  w2_3 = io_din[7]; // @[el2_lib.scala 345:39]
  wire  w0_5 = io_din[8]; // @[el2_lib.scala 343:39]
  wire  w1_5 = io_din[9]; // @[el2_lib.scala 344:39]
  wire  w0_6 = io_din[10]; // @[el2_lib.scala 343:39]
  wire  w0_7 = io_din[11]; // @[el2_lib.scala 343:39]
  wire  w1_7 = io_din[12]; // @[el2_lib.scala 344:39]
  wire  w0_8 = io_din[13]; // @[el2_lib.scala 343:39]
  wire  w2_7 = io_din[14]; // @[el2_lib.scala 345:39]
  wire  w0_9 = io_din[15]; // @[el2_lib.scala 343:39]
  wire  w1_9 = io_din[16]; // @[el2_lib.scala 344:39]
  wire  w0_10 = io_din[17]; // @[el2_lib.scala 343:39]
  wire  w3_7 = io_din[18]; // @[el2_lib.scala 346:39]
  wire  w0_11 = io_din[19]; // @[el2_lib.scala 343:39]
  wire  w1_11 = io_din[20]; // @[el2_lib.scala 344:39]
  wire  w0_12 = io_din[21]; // @[el2_lib.scala 343:39]
  wire  w2_11 = io_din[22]; // @[el2_lib.scala 345:39]
  wire  w0_13 = io_din[23]; // @[el2_lib.scala 343:39]
  wire  w1_13 = io_din[24]; // @[el2_lib.scala 344:39]
  wire  w0_14 = io_din[25]; // @[el2_lib.scala 343:39]
  wire  w0_15 = io_din[26]; // @[el2_lib.scala 343:39]
  wire  w1_15 = io_din[27]; // @[el2_lib.scala 344:39]
  wire  w0_16 = io_din[28]; // @[el2_lib.scala 343:39]
  wire  w2_15 = io_din[29]; // @[el2_lib.scala 345:39]
  wire  w0_17 = io_din[30]; // @[el2_lib.scala 343:39]
  wire  w1_17 = io_din[31]; // @[el2_lib.scala 344:39]
  wire  w0_18 = io_din[32]; // @[el2_lib.scala 343:39]
  wire  w3_15 = io_din[33]; // @[el2_lib.scala 346:39]
  wire  w0_19 = io_din[34]; // @[el2_lib.scala 343:39]
  wire  w1_19 = io_din[35]; // @[el2_lib.scala 344:39]
  wire  w0_20 = io_din[36]; // @[el2_lib.scala 343:39]
  wire  w2_19 = io_din[37]; // @[el2_lib.scala 345:39]
  wire  w0_21 = io_din[38]; // @[el2_lib.scala 343:39]
  wire  w1_21 = io_din[39]; // @[el2_lib.scala 344:39]
  wire  w0_22 = io_din[40]; // @[el2_lib.scala 343:39]
  wire  w4_15 = io_din[41]; // @[el2_lib.scala 347:39]
  wire  w0_23 = io_din[42]; // @[el2_lib.scala 343:39]
  wire  w1_23 = io_din[43]; // @[el2_lib.scala 344:39]
  wire  w0_24 = io_din[44]; // @[el2_lib.scala 343:39]
  wire  w2_23 = io_din[45]; // @[el2_lib.scala 345:39]
  wire  w0_25 = io_din[46]; // @[el2_lib.scala 343:39]
  wire  w1_25 = io_din[47]; // @[el2_lib.scala 344:39]
  wire  w0_26 = io_din[48]; // @[el2_lib.scala 343:39]
  wire  w3_23 = io_din[49]; // @[el2_lib.scala 346:39]
  wire  w0_27 = io_din[50]; // @[el2_lib.scala 343:39]
  wire  w1_27 = io_din[51]; // @[el2_lib.scala 344:39]
  wire  w0_28 = io_din[52]; // @[el2_lib.scala 343:39]
  wire  w2_27 = io_din[53]; // @[el2_lib.scala 345:39]
  wire  w0_29 = io_din[54]; // @[el2_lib.scala 343:39]
  wire  w1_29 = io_din[55]; // @[el2_lib.scala 344:39]
  wire  w0_30 = io_din[56]; // @[el2_lib.scala 343:39]
  wire  w0_31 = io_din[57]; // @[el2_lib.scala 343:39]
  wire  w1_31 = io_din[58]; // @[el2_lib.scala 344:39]
  wire  w0_32 = io_din[59]; // @[el2_lib.scala 343:39]
  wire  w2_31 = io_din[60]; // @[el2_lib.scala 345:39]
  wire  w0_33 = io_din[61]; // @[el2_lib.scala 343:39]
  wire  w1_33 = io_din[62]; // @[el2_lib.scala 344:39]
  wire  w0_34 = io_din[63]; // @[el2_lib.scala 343:39]
  wire [6:0] _T_210 = {w0_34,w1_33,w0_33,w2_31,w0_32,w1_31,w0_31}; // @[el2_lib.scala 351:27]
  wire  _T_211 = ^_T_210; // @[el2_lib.scala 351:34]
  wire [6:0] _T_217 = {w0_18,w1_17,w0_17,w2_15,w0_16,w1_15,w0_15}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_224 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15}; // @[el2_lib.scala 351:44]
  wire [14:0] _T_225 = {w0_22,w1_21,w0_21,w2_19,w0_20,w1_19,w0_19,w3_15,_T_217}; // @[el2_lib.scala 351:44]
  wire [7:0] _T_232 = {w0_26,w1_25,w0_25,w2_23,w0_24,w1_23,w0_23,w4_15}; // @[el2_lib.scala 351:44]
  wire [30:0] _T_241 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_225}; // @[el2_lib.scala 351:44]
  wire  _T_242 = ^_T_241; // @[el2_lib.scala 351:51]
  wire [6:0] _T_248 = {w0_10,w1_9,w0_9,w2_7,w0_8,w1_7,w0_7}; // @[el2_lib.scala 351:61]
  wire [14:0] _T_256 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_248}; // @[el2_lib.scala 351:61]
  wire [30:0] _T_272 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_232,_T_256}; // @[el2_lib.scala 351:61]
  wire  _T_273 = ^_T_272; // @[el2_lib.scala 351:68]
  wire [6:0] _T_279 = {w0_6,w1_5,w0_5,w2_3,w0_4,w1_3,w0_3}; // @[el2_lib.scala 351:78]
  wire [14:0] _T_287 = {w0_14,w1_13,w0_13,w2_11,w0_12,w1_11,w0_11,w3_7,_T_279}; // @[el2_lib.scala 351:78]
  wire [30:0] _T_303 = {w0_30,w1_29,w0_29,w2_27,w0_28,w1_27,w0_27,w3_23,_T_224,_T_287}; // @[el2_lib.scala 351:78]
  wire  _T_304 = ^_T_303; // @[el2_lib.scala 351:85]
  wire [7:0] _T_311 = {w2_7,w0_6,w1_5,w0_5,w2_3,w0_2,w1_1,w0_1}; // @[el2_lib.scala 351:95]
  wire [16:0] _T_320 = {w0_17,w2_15,w0_14,w1_13,w0_13,w2_11,w0_10,w1_9,w0_9,_T_311}; // @[el2_lib.scala 351:95]
  wire [8:0] _T_328 = {w1_25,w0_25,w2_23,w0_22,w1_21,w0_21,w2_19,w0_18,w1_17}; // @[el2_lib.scala 351:95]
  wire [17:0] _T_337 = {w0_34,w1_33,w0_33,w2_31,w0_30,w1_29,w0_29,w2_27,w0_26,_T_328}; // @[el2_lib.scala 351:95]
  wire [34:0] _T_338 = {_T_337,_T_320}; // @[el2_lib.scala 351:95]
  wire  _T_339 = ^_T_338; // @[el2_lib.scala 351:102]
  wire [7:0] _T_346 = {w1_7,w0_6,w1_5,w0_4,w1_3,w0_2,w1_1,w0_0}; // @[el2_lib.scala 351:112]
  wire [16:0] _T_355 = {w0_16,w1_15,w0_14,w1_13,w0_12,w1_11,w0_10,w1_9,w0_8,_T_346}; // @[el2_lib.scala 351:112]
  wire [8:0] _T_363 = {w1_25,w0_24,w1_23,w0_22,w1_21,w0_20,w1_19,w0_18,w1_17}; // @[el2_lib.scala 351:112]
  wire [17:0] _T_372 = {w0_34,w1_33,w0_32,w1_31,w0_30,w1_29,w0_28,w1_27,w0_26,_T_363}; // @[el2_lib.scala 351:112]
  wire [34:0] _T_373 = {_T_372,_T_355}; // @[el2_lib.scala 351:112]
  wire  _T_374 = ^_T_373; // @[el2_lib.scala 351:119]
  wire [7:0] _T_381 = {w0_7,w0_6,w0_5,w0_4,w0_3,w0_2,w0_1,w0_0}; // @[el2_lib.scala 351:129]
  wire [16:0] _T_390 = {w0_16,w0_15,w0_14,w0_13,w0_12,w0_11,w0_10,w0_9,w0_8,_T_381}; // @[el2_lib.scala 351:129]
  wire [8:0] _T_398 = {w0_25,w0_24,w0_23,w0_22,w0_21,w0_20,w0_19,w0_18,w0_17}; // @[el2_lib.scala 351:129]
  wire [17:0] _T_407 = {w0_34,w0_33,w0_32,w0_31,w0_30,w0_29,w0_28,w0_27,w0_26,_T_398}; // @[el2_lib.scala 351:129]
  wire [34:0] _T_408 = {_T_407,_T_390}; // @[el2_lib.scala 351:129]
  wire  _T_409 = ^_T_408; // @[el2_lib.scala 351:136]
  wire [2:0] _T_411 = {_T_339,_T_374,_T_409}; // @[Cat.scala 29:58]
  wire [3:0] _T_414 = {_T_211,_T_242,_T_273,_T_304}; // @[Cat.scala 29:58]
  assign io_ecc_out = {_T_414,_T_411}; // @[el2_lib.scala 351:16]
endmodule
module el2_ifu_mem_ctl(
  input          clock,
  input          reset,
  input          io_free_clk,
  input          io_active_clk,
  input          io_exu_flush_final,
  input          io_dec_tlu_flush_lower_wb,
  input          io_dec_tlu_flush_err_wb,
  input          io_dec_tlu_i0_commit_cmt,
  input          io_dec_tlu_force_halt,
  input  [30:0]  io_ifc_fetch_addr_bf,
  input          io_ifc_fetch_uncacheable_bf,
  input          io_ifc_fetch_req_bf,
  input          io_ifc_fetch_req_bf_raw,
  input          io_ifc_iccm_access_bf,
  input          io_ifc_region_acc_fault_bf,
  input          io_ifc_dma_access_ok,
  input          io_dec_tlu_fence_i_wb,
  input          io_ifu_bp_hit_taken_f,
  input          io_ifu_bp_inst_mask_f,
  input          io_ifu_axi_arready,
  input          io_ifu_axi_rvalid,
  input  [2:0]   io_ifu_axi_rid,
  input  [63:0]  io_ifu_axi_rdata,
  input  [1:0]   io_ifu_axi_rresp,
  input          io_ifu_bus_clk_en,
  input          io_dma_iccm_req,
  input  [31:0]  io_dma_mem_addr,
  input  [2:0]   io_dma_mem_sz,
  input          io_dma_mem_write,
  input  [63:0]  io_dma_mem_wdata,
  input  [2:0]   io_dma_mem_tag,
  input  [63:0]  io_ic_rd_data,
  input  [70:0]  io_ic_debug_rd_data,
  input  [25:0]  io_ictag_debug_rd_data,
  input  [1:0]   io_ic_eccerr,
  input  [1:0]   io_ic_parerr,
  input  [1:0]   io_ic_rd_hit,
  input          io_ic_tag_perr,
  input  [63:0]  io_iccm_rd_data,
  input  [77:0]  io_iccm_rd_data_ecc,
  input  [1:0]   io_ifu_fetch_val,
  input  [70:0]  io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0]  io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input          io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input          io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output         io_ifu_miss_state_idle,
  output         io_ifu_ic_mb_empty,
  output         io_ic_dma_active,
  output         io_ic_write_stall,
  output         io_ifu_pmu_ic_miss,
  output         io_ifu_pmu_ic_hit,
  output         io_ifu_pmu_bus_error,
  output         io_ifu_pmu_bus_busy,
  output         io_ifu_pmu_bus_trxn,
  output         io_ifu_axi_awvalid,
  output [2:0]   io_ifu_axi_awid,
  output [31:0]  io_ifu_axi_awaddr,
  output [3:0]   io_ifu_axi_awregion,
  output [7:0]   io_ifu_axi_awlen,
  output [2:0]   io_ifu_axi_awsize,
  output [1:0]   io_ifu_axi_awburst,
  output         io_ifu_axi_awlock,
  output [3:0]   io_ifu_axi_awcache,
  output [2:0]   io_ifu_axi_awprot,
  output [3:0]   io_ifu_axi_awqos,
  output         io_ifu_axi_wvalid,
  output [63:0]  io_ifu_axi_wdata,
  output [7:0]   io_ifu_axi_wstrb,
  output         io_ifu_axi_wlast,
  output         io_ifu_axi_bready,
  output         io_ifu_axi_arvalid,
  output [2:0]   io_ifu_axi_arid,
  output [31:0]  io_ifu_axi_araddr,
  output [3:0]   io_ifu_axi_arregion,
  output [7:0]   io_ifu_axi_arlen,
  output [2:0]   io_ifu_axi_arsize,
  output [1:0]   io_ifu_axi_arburst,
  output         io_ifu_axi_arlock,
  output [3:0]   io_ifu_axi_arcache,
  output [2:0]   io_ifu_axi_arprot,
  output [3:0]   io_ifu_axi_arqos,
  output         io_ifu_axi_rready,
  output         io_iccm_dma_ecc_error,
  output         io_iccm_dma_rvalid,
  output [63:0]  io_iccm_dma_rdata,
  output [2:0]   io_iccm_dma_rtag,
  output         io_iccm_ready,
  output [30:0]  io_ic_rw_addr,
  output [1:0]   io_ic_wr_en,
  output         io_ic_rd_en,
  output [70:0]  io_ic_wr_data_0,
  output [70:0]  io_ic_wr_data_1,
  output [70:0]  io_ic_debug_wr_data,
  output [70:0]  io_ifu_ic_debug_rd_data,
  output [9:0]   io_ic_debug_addr,
  output         io_ic_debug_rd_en,
  output         io_ic_debug_wr_en,
  output         io_ic_debug_tag_array,
  output [1:0]   io_ic_debug_way,
  output [1:0]   io_ic_tag_valid,
  output [14:0]  io_iccm_rw_addr,
  output         io_iccm_wren,
  output         io_iccm_rden,
  output [77:0]  io_iccm_wr_data,
  output [2:0]   io_iccm_wr_size,
  output         io_ic_hit_f,
  output         io_ic_access_fault_f,
  output [1:0]   io_ic_access_fault_type_f,
  output         io_iccm_rd_ecc_single_err,
  output         io_iccm_rd_ecc_double_err,
  output         io_ic_error_start,
  output         io_ifu_async_error_start,
  output         io_iccm_dma_sb_error,
  output [1:0]   io_ic_fetch_val_f,
  output [31:0]  io_ic_data_f,
  output [63:0]  io_ic_premux_data,
  output         io_ic_sel_premux_data,
  input          io_dec_tlu_core_ecc_disable,
  output         io_ifu_ic_debug_rd_data_valid,
  output         io_iccm_buf_correct_ecc,
  output         io_iccm_correction_state,
  input          io_scan_mode,
  output [141:0] io_data,
  output [63:0]  io_ic_miss_buff_half,
  output [6:0]   io_ic_wr_ecc
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [63:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [95:0] _RAND_441;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [63:0] _RAND_449;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [63:0] _RAND_454;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] m1_io_din; // @[el2_ifu_mem_ctl.scala 346:18]
  wire [6:0] m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 346:18]
  wire [63:0] m2_io_din; // @[el2_ifu_mem_ctl.scala 347:18]
  wire [6:0] m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 347:18]
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 188:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 324:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 325:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 325:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 257:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 561:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 563:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 190:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 312:34]
  wire [4:0] _GEN_464 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 678:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_464 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 678:53]
  wire [1:0] _GEN_465 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 681:91]
  wire [1:0] _T_2278 = ic_fetch_val_shift_right[3:2] & _GEN_465; // @[el2_ifu_mem_ctl.scala 681:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 326:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 279:46]
  wire [1:0] _GEN_466 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 681:113]
  wire [1:0] _T_2279 = _T_2278 & _GEN_466; // @[el2_ifu_mem_ctl.scala 681:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 667:59]
  wire [1:0] _GEN_467 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 681:130]
  wire [1:0] _T_2280 = _T_2279 | _GEN_467; // @[el2_ifu_mem_ctl.scala 681:130]
  wire  _T_2281 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 681:154]
  wire [1:0] _GEN_468 = {{1'd0}, _T_2281}; // @[el2_ifu_mem_ctl.scala 681:152]
  wire [1:0] _T_2282 = _T_2280 & _GEN_468; // @[el2_ifu_mem_ctl.scala 681:152]
  wire [1:0] _T_2271 = ic_fetch_val_shift_right[1:0] & _GEN_465; // @[el2_ifu_mem_ctl.scala 681:91]
  wire [1:0] _T_2272 = _T_2271 & _GEN_466; // @[el2_ifu_mem_ctl.scala 681:113]
  wire [1:0] _T_2273 = _T_2272 | _GEN_467; // @[el2_ifu_mem_ctl.scala 681:130]
  wire [1:0] _T_2275 = _T_2273 & _GEN_468; // @[el2_ifu_mem_ctl.scala 681:152]
  wire [3:0] iccm_ecc_word_enable = {_T_2282,_T_2275}; // @[Cat.scala 29:58]
  wire  _T_2382 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 301:30]
  wire  _T_2383 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 301:44]
  wire  _T_2384 = _T_2382 ^ _T_2383; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2392 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 301:76]
  wire  _T_2393 = ^_T_2392; // @[el2_lib.scala 301:83]
  wire  _T_2394 = io_iccm_rd_data_ecc[37] ^ _T_2393; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2401 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2409 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2401}; // @[el2_lib.scala 301:103]
  wire  _T_2410 = ^_T_2409; // @[el2_lib.scala 301:110]
  wire  _T_2411 = io_iccm_rd_data_ecc[36] ^ _T_2410; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2418 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2426 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_2418}; // @[el2_lib.scala 301:130]
  wire  _T_2427 = ^_T_2426; // @[el2_lib.scala 301:137]
  wire  _T_2428 = io_iccm_rd_data_ecc[35] ^ _T_2427; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2437 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2446 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2437}; // @[el2_lib.scala 301:157]
  wire  _T_2447 = ^_T_2446; // @[el2_lib.scala 301:164]
  wire  _T_2448 = io_iccm_rd_data_ecc[34] ^ _T_2447; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2457 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2466 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_2457}; // @[el2_lib.scala 301:184]
  wire  _T_2467 = ^_T_2466; // @[el2_lib.scala 301:191]
  wire  _T_2468 = io_iccm_rd_data_ecc[33] ^ _T_2467; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2477 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2486 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_2477}; // @[el2_lib.scala 301:211]
  wire  _T_2487 = ^_T_2486; // @[el2_lib.scala 301:218]
  wire  _T_2488 = io_iccm_rd_data_ecc[32] ^ _T_2487; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2494 = {_T_2384,_T_2394,_T_2411,_T_2428,_T_2448,_T_2468,_T_2488}; // @[Cat.scala 29:58]
  wire  _T_2495 = _T_2494 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2496 = iccm_ecc_word_enable[0] & _T_2495; // @[el2_lib.scala 302:32]
  wire  _T_2498 = _T_2496 & _T_2494[6]; // @[el2_lib.scala 302:53]
  wire  _T_2767 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 301:30]
  wire  _T_2768 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 301:44]
  wire  _T_2769 = _T_2767 ^ _T_2768; // @[el2_lib.scala 301:35]
  wire [5:0] _T_2777 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 301:76]
  wire  _T_2778 = ^_T_2777; // @[el2_lib.scala 301:83]
  wire  _T_2779 = io_iccm_rd_data_ecc[76] ^ _T_2778; // @[el2_lib.scala 301:71]
  wire [6:0] _T_2786 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 301:103]
  wire [14:0] _T_2794 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2786}; // @[el2_lib.scala 301:103]
  wire  _T_2795 = ^_T_2794; // @[el2_lib.scala 301:110]
  wire  _T_2796 = io_iccm_rd_data_ecc[75] ^ _T_2795; // @[el2_lib.scala 301:98]
  wire [6:0] _T_2803 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 301:130]
  wire [14:0] _T_2811 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_2803}; // @[el2_lib.scala 301:130]
  wire  _T_2812 = ^_T_2811; // @[el2_lib.scala 301:137]
  wire  _T_2813 = io_iccm_rd_data_ecc[74] ^ _T_2812; // @[el2_lib.scala 301:125]
  wire [8:0] _T_2822 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 301:157]
  wire [17:0] _T_2831 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2822}; // @[el2_lib.scala 301:157]
  wire  _T_2832 = ^_T_2831; // @[el2_lib.scala 301:164]
  wire  _T_2833 = io_iccm_rd_data_ecc[73] ^ _T_2832; // @[el2_lib.scala 301:152]
  wire [8:0] _T_2842 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:184]
  wire [17:0] _T_2851 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_2842}; // @[el2_lib.scala 301:184]
  wire  _T_2852 = ^_T_2851; // @[el2_lib.scala 301:191]
  wire  _T_2853 = io_iccm_rd_data_ecc[72] ^ _T_2852; // @[el2_lib.scala 301:179]
  wire [8:0] _T_2862 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 301:211]
  wire [17:0] _T_2871 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_2862}; // @[el2_lib.scala 301:211]
  wire  _T_2872 = ^_T_2871; // @[el2_lib.scala 301:218]
  wire  _T_2873 = io_iccm_rd_data_ecc[71] ^ _T_2872; // @[el2_lib.scala 301:206]
  wire [6:0] _T_2879 = {_T_2769,_T_2779,_T_2796,_T_2813,_T_2833,_T_2853,_T_2873}; // @[Cat.scala 29:58]
  wire  _T_2880 = _T_2879 != 7'h0; // @[el2_lib.scala 302:44]
  wire  _T_2881 = iccm_ecc_word_enable[1] & _T_2880; // @[el2_lib.scala 302:32]
  wire  _T_2883 = _T_2881 & _T_2879[6]; // @[el2_lib.scala 302:53]
  wire [1:0] iccm_single_ecc_error = {_T_2498,_T_2883}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 193:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 645:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 194:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 195:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 490:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 195:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 195:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 195:72]
  wire  _T_1647 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1652 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1672 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 540:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 404:42]
  wire  _T_1674 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 540:79]
  wire  _T_1675 = _T_1672 | _T_1674; // @[el2_ifu_mem_ctl.scala 540:56]
  wire  _T_1676 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 540:122]
  wire  _T_1677 = ~_T_1676; // @[el2_ifu_mem_ctl.scala 540:101]
  wire  _T_1678 = _T_1675 & _T_1677; // @[el2_ifu_mem_ctl.scala 540:99]
  wire  _T_1679 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_1693 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 547:45]
  wire  _T_1694 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 547:69]
  wire  _T_1695 = _T_1693 & _T_1694; // @[el2_ifu_mem_ctl.scala 547:67]
  wire  _T_1696 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_1679 ? _T_1695 : _T_1696; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_1652 ? _T_1678 : _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_1647 ? 1'h0 : _GEN_59; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 195:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 197:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 197:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 287:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 287:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 713:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 287:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 278:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 278:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 328:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 278:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 278:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 287:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 287:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 287:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 287:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 287:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 560:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 602:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 629:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 314:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 610:56]
  wire  _T_1798 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 627:69]
  wire  _T_1799 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 627:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_1798 : _T_1799; // @[el2_ifu_mem_ctl.scala 627:28]
  wire  _T_1745 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 606:68]
  wire  _T_1746 = ic_act_miss_f | _T_1745; // @[el2_ifu_mem_ctl.scala 606:48]
  wire  bus_reset_data_beat_cnt = _T_1746 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 606:91]
  wire  _T_1742 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 605:50]
  wire  _T_1743 = bus_ifu_wr_en_ff & _T_1742; // @[el2_ifu_mem_ctl.scala 605:48]
  wire  _T_1744 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 605:72]
  wire  bus_inc_data_beat_cnt = _T_1743 & _T_1744; // @[el2_ifu_mem_ctl.scala 605:70]
  wire [2:0] _T_1750 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 609:115]
  wire [2:0] _T_1752 = bus_inc_data_beat_cnt ? _T_1750 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_1747 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 607:32]
  wire  _T_1748 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 607:57]
  wire  bus_hold_data_beat_cnt = _T_1747 & _T_1748; // @[el2_ifu_mem_ctl.scala 607:55]
  wire [2:0] _T_1753 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_1752 | _T_1753; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 197:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 197:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 198:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 197:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 198:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 204:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 204:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 440:45]
  wire  _T_1277 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 461:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 417:60]
  wire  _T_1308 = _T_1277 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1281 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 461:127]
  wire  _T_1309 = _T_1281 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1316 = _T_1308 | _T_1309; // @[Mux.scala 27:72]
  wire  _T_1285 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 461:127]
  wire  _T_1310 = _T_1285 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1317 = _T_1316 | _T_1310; // @[Mux.scala 27:72]
  wire  _T_1289 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 461:127]
  wire  _T_1311 = _T_1289 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1318 = _T_1317 | _T_1311; // @[Mux.scala 27:72]
  wire  _T_1293 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 461:127]
  wire  _T_1312 = _T_1293 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1319 = _T_1318 | _T_1312; // @[Mux.scala 27:72]
  wire  _T_1297 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 461:127]
  wire  _T_1313 = _T_1297 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1320 = _T_1319 | _T_1313; // @[Mux.scala 27:72]
  wire  _T_1301 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 461:127]
  wire  _T_1314 = _T_1301 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1321 = _T_1320 | _T_1314; // @[Mux.scala 27:72]
  wire  _T_1305 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 461:127]
  wire  _T_1315 = _T_1305 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_1321 | _T_1315; // @[Mux.scala 27:72]
  wire  _T_1363 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 463:69]
  wire  _T_1364 = ic_miss_buff_data_valid_bypass_index & _T_1363; // @[el2_ifu_mem_ctl.scala 463:67]
  wire  _T_1366 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 463:91]
  wire  _T_1367 = _T_1364 & _T_1366; // @[el2_ifu_mem_ctl.scala 463:89]
  wire  _T_1372 = _T_1364 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 464:65]
  wire  _T_1373 = _T_1367 | _T_1372; // @[el2_ifu_mem_ctl.scala 463:112]
  wire  _T_1375 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 465:43]
  wire  _T_1378 = _T_1375 & _T_1366; // @[el2_ifu_mem_ctl.scala 465:65]
  wire  _T_1379 = _T_1373 | _T_1378; // @[el2_ifu_mem_ctl.scala 464:88]
  wire  _T_1383 = _T_1375 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 466:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 443:75]
  wire  _T_1323 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1347 = _T_1323 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1326 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1348 = _T_1326 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1355 = _T_1347 | _T_1348; // @[Mux.scala 27:72]
  wire  _T_1329 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1349 = _T_1329 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1356 = _T_1355 | _T_1349; // @[Mux.scala 27:72]
  wire  _T_1332 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1350 = _T_1332 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1357 = _T_1356 | _T_1350; // @[Mux.scala 27:72]
  wire  _T_1335 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1351 = _T_1335 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1358 = _T_1357 | _T_1351; // @[Mux.scala 27:72]
  wire  _T_1338 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1352 = _T_1338 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1359 = _T_1358 | _T_1352; // @[Mux.scala 27:72]
  wire  _T_1341 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1353 = _T_1341 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1360 = _T_1359 | _T_1353; // @[Mux.scala 27:72]
  wire  _T_1344 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 462:110]
  wire  _T_1354 = _T_1344 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_1360 | _T_1354; // @[Mux.scala 27:72]
  wire  _T_1384 = _T_1383 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 466:87]
  wire  _T_1385 = _T_1379 | _T_1384; // @[el2_ifu_mem_ctl.scala 465:88]
  wire  _T_1389 = ic_miss_buff_data_valid_bypass_index & _T_1305; // @[el2_ifu_mem_ctl.scala 467:43]
  wire  miss_buff_hit_unq_f = _T_1385 | _T_1389; // @[el2_ifu_mem_ctl.scala 466:131]
  wire  _T_1405 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 472:55]
  wire  _T_1406 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 472:87]
  wire  _T_1407 = _T_1405 | _T_1406; // @[el2_ifu_mem_ctl.scala 472:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_1407; // @[el2_ifu_mem_ctl.scala 472:41]
  wire  _T_1390 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 469:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 315:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[6]; // @[el2_ifu_mem_ctl.scala 460:51]
  wire  _T_1391 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 469:68]
  wire  _T_1392 = miss_buff_hit_unq_f & _T_1391; // @[el2_ifu_mem_ctl.scala 469:66]
  wire  stream_hit_f = _T_1390 & _T_1392; // @[el2_ifu_mem_ctl.scala 469:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 282:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 282:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 282:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 612:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 639:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 208:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 208:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 208:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 208:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 208:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 209:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 209:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 209:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 210:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 210:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 210:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 210:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 211:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 212:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 212:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 212:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 200:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 212:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 212:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 213:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 213:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 213:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 213:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 214:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 215:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 215:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 215:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 214:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 213:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 212:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 211:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 210:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 209:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 208:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_1402 = byp_fetch_index[4:1] == 4'h7; // @[el2_ifu_mem_ctl.scala 471:60]
  wire  _T_1403 = _T_1402 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 471:92]
  wire  stream_eol_f = _T_1403 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 471:110]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 223:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 223:87]
  wire  _T_113 = _T_111 & _T_1744; // @[el2_ifu_mem_ctl.scala 223:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 223:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 227:48]
  wire  _T_126 = _T_124 & _T_1744; // @[el2_ifu_mem_ctl.scala 227:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 227:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 288:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 288:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 288:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 288:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 288:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 289:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 288:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 289:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 342:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 289:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 289:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 289:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 231:50]
  wire  _T_137 = _T_135 & _T_1744; // @[el2_ifu_mem_ctl.scala 231:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 290:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 291:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 291:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 290:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 232:35]
  wire  _T_143 = _T_141 & _T_1744; // @[el2_ifu_mem_ctl.scala 232:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 232:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 231:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 237:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 236:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 236:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 241:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 241:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 198:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 198:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 198:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 198:91]
  wire  _T_30 = ic_act_miss_f & _T_1744; // @[el2_ifu_mem_ctl.scala 205:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 216:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 216:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 216:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 216:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 216:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 216:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 220:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 220:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 220:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 224:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 224:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 228:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 228:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 233:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 233:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 233:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 238:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 238:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 258:95]
  wire  _T_175 = _T_1405 & _T_174; // @[el2_ifu_mem_ctl.scala 258:93]
  wire  crit_wd_byp_ok_ff = _T_1406 | _T_175; // @[el2_ifu_mem_ctl.scala 258:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 259:36]
  wire  _T_180 = _T_1405 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 259:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 259:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 259:70]
  wire  _T_184 = _T_1405 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 260:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 260:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 259:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 260:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 261:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 261:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 260:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 263:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 263:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 271:35]
  reg [6:0] _T_4323; // @[el2_ifu_mem_ctl.scala 741:14]
  wire [5:0] ifu_ic_rw_int_addr_ff = _T_4323[5:0]; // @[el2_ifu_mem_ctl.scala 740:27]
  wire [6:0] _GEN_473 = {{1'd0}, ifu_ic_rw_int_addr_ff}; // @[el2_ifu_mem_ctl.scala 737:121]
  wire  _T_4188 = _GEN_473 == 7'h7f; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4190 = _T_4188 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3679; // @[Reg.scala 27:20]
  wire  way_status_out_127 = _T_3679[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_474 = {{5'd0}, way_status_out_127}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4191 = _T_4190 & _GEN_474; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4184 = _GEN_473 == 7'h7e; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4186 = _T_4184 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3675; // @[Reg.scala 27:20]
  wire  way_status_out_126 = _T_3675[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_476 = {{5'd0}, way_status_out_126}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4187 = _T_4186 & _GEN_476; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4180 = _GEN_473 == 7'h7d; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4182 = _T_4180 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3671; // @[Reg.scala 27:20]
  wire  way_status_out_125 = _T_3671[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_478 = {{5'd0}, way_status_out_125}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4183 = _T_4182 & _GEN_478; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4176 = _GEN_473 == 7'h7c; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4178 = _T_4176 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3667; // @[Reg.scala 27:20]
  wire  way_status_out_124 = _T_3667[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_480 = {{5'd0}, way_status_out_124}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4179 = _T_4178 & _GEN_480; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4172 = _GEN_473 == 7'h7b; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4174 = _T_4172 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3663; // @[Reg.scala 27:20]
  wire  way_status_out_123 = _T_3663[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_482 = {{5'd0}, way_status_out_123}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4175 = _T_4174 & _GEN_482; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4168 = _GEN_473 == 7'h7a; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4170 = _T_4168 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3659; // @[Reg.scala 27:20]
  wire  way_status_out_122 = _T_3659[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_484 = {{5'd0}, way_status_out_122}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4171 = _T_4170 & _GEN_484; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4164 = _GEN_473 == 7'h79; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4166 = _T_4164 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3655; // @[Reg.scala 27:20]
  wire  way_status_out_121 = _T_3655[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_486 = {{5'd0}, way_status_out_121}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4167 = _T_4166 & _GEN_486; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4160 = _GEN_473 == 7'h78; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4162 = _T_4160 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3651; // @[Reg.scala 27:20]
  wire  way_status_out_120 = _T_3651[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_488 = {{5'd0}, way_status_out_120}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4163 = _T_4162 & _GEN_488; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4156 = _GEN_473 == 7'h77; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4158 = _T_4156 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3647; // @[Reg.scala 27:20]
  wire  way_status_out_119 = _T_3647[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_490 = {{5'd0}, way_status_out_119}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4159 = _T_4158 & _GEN_490; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4152 = _GEN_473 == 7'h76; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4154 = _T_4152 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3643; // @[Reg.scala 27:20]
  wire  way_status_out_118 = _T_3643[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_492 = {{5'd0}, way_status_out_118}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4155 = _T_4154 & _GEN_492; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [59:0] _T_4200 = {_T_4191,_T_4187,_T_4183,_T_4179,_T_4175,_T_4171,_T_4167,_T_4163,_T_4159,_T_4155}; // @[Cat.scala 29:58]
  wire  _T_4148 = _GEN_473 == 7'h75; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4150 = _T_4148 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3639; // @[Reg.scala 27:20]
  wire  way_status_out_117 = _T_3639[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_494 = {{5'd0}, way_status_out_117}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4151 = _T_4150 & _GEN_494; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4144 = _GEN_473 == 7'h74; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4146 = _T_4144 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3635; // @[Reg.scala 27:20]
  wire  way_status_out_116 = _T_3635[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_496 = {{5'd0}, way_status_out_116}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4147 = _T_4146 & _GEN_496; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4140 = _GEN_473 == 7'h73; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4142 = _T_4140 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3631; // @[Reg.scala 27:20]
  wire  way_status_out_115 = _T_3631[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_498 = {{5'd0}, way_status_out_115}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4143 = _T_4142 & _GEN_498; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4136 = _GEN_473 == 7'h72; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4138 = _T_4136 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3627; // @[Reg.scala 27:20]
  wire  way_status_out_114 = _T_3627[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_500 = {{5'd0}, way_status_out_114}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4139 = _T_4138 & _GEN_500; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4132 = _GEN_473 == 7'h71; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4134 = _T_4132 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3623; // @[Reg.scala 27:20]
  wire  way_status_out_113 = _T_3623[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_502 = {{5'd0}, way_status_out_113}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4135 = _T_4134 & _GEN_502; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4128 = _GEN_473 == 7'h70; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4130 = _T_4128 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3619; // @[Reg.scala 27:20]
  wire  way_status_out_112 = _T_3619[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_504 = {{5'd0}, way_status_out_112}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4131 = _T_4130 & _GEN_504; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4124 = _GEN_473 == 7'h6f; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4126 = _T_4124 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3615; // @[Reg.scala 27:20]
  wire  way_status_out_111 = _T_3615[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_506 = {{5'd0}, way_status_out_111}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4127 = _T_4126 & _GEN_506; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4120 = _GEN_473 == 7'h6e; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4122 = _T_4120 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3611; // @[Reg.scala 27:20]
  wire  way_status_out_110 = _T_3611[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_508 = {{5'd0}, way_status_out_110}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4123 = _T_4122 & _GEN_508; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4116 = _GEN_473 == 7'h6d; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4118 = _T_4116 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3607; // @[Reg.scala 27:20]
  wire  way_status_out_109 = _T_3607[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_510 = {{5'd0}, way_status_out_109}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4119 = _T_4118 & _GEN_510; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [113:0] _T_4209 = {_T_4200,_T_4151,_T_4147,_T_4143,_T_4139,_T_4135,_T_4131,_T_4127,_T_4123,_T_4119}; // @[Cat.scala 29:58]
  wire  _T_4112 = _GEN_473 == 7'h6c; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4114 = _T_4112 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3603; // @[Reg.scala 27:20]
  wire  way_status_out_108 = _T_3603[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_512 = {{5'd0}, way_status_out_108}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4115 = _T_4114 & _GEN_512; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4108 = _GEN_473 == 7'h6b; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4110 = _T_4108 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3599; // @[Reg.scala 27:20]
  wire  way_status_out_107 = _T_3599[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_514 = {{5'd0}, way_status_out_107}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4111 = _T_4110 & _GEN_514; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4104 = _GEN_473 == 7'h6a; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4106 = _T_4104 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3595; // @[Reg.scala 27:20]
  wire  way_status_out_106 = _T_3595[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_516 = {{5'd0}, way_status_out_106}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4107 = _T_4106 & _GEN_516; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4100 = _GEN_473 == 7'h69; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4102 = _T_4100 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3591; // @[Reg.scala 27:20]
  wire  way_status_out_105 = _T_3591[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_518 = {{5'd0}, way_status_out_105}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4103 = _T_4102 & _GEN_518; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4096 = _GEN_473 == 7'h68; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4098 = _T_4096 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3587; // @[Reg.scala 27:20]
  wire  way_status_out_104 = _T_3587[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_520 = {{5'd0}, way_status_out_104}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4099 = _T_4098 & _GEN_520; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4092 = _GEN_473 == 7'h67; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4094 = _T_4092 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3583; // @[Reg.scala 27:20]
  wire  way_status_out_103 = _T_3583[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_522 = {{5'd0}, way_status_out_103}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4095 = _T_4094 & _GEN_522; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4088 = _GEN_473 == 7'h66; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4090 = _T_4088 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3579; // @[Reg.scala 27:20]
  wire  way_status_out_102 = _T_3579[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_524 = {{5'd0}, way_status_out_102}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4091 = _T_4090 & _GEN_524; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4084 = _GEN_473 == 7'h65; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4086 = _T_4084 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3575; // @[Reg.scala 27:20]
  wire  way_status_out_101 = _T_3575[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_526 = {{5'd0}, way_status_out_101}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4087 = _T_4086 & _GEN_526; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4080 = _GEN_473 == 7'h64; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4082 = _T_4080 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3571; // @[Reg.scala 27:20]
  wire  way_status_out_100 = _T_3571[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_528 = {{5'd0}, way_status_out_100}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4083 = _T_4082 & _GEN_528; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [167:0] _T_4218 = {_T_4209,_T_4115,_T_4111,_T_4107,_T_4103,_T_4099,_T_4095,_T_4091,_T_4087,_T_4083}; // @[Cat.scala 29:58]
  wire  _T_4076 = _GEN_473 == 7'h63; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4078 = _T_4076 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3567; // @[Reg.scala 27:20]
  wire  way_status_out_99 = _T_3567[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_530 = {{5'd0}, way_status_out_99}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4079 = _T_4078 & _GEN_530; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4072 = _GEN_473 == 7'h62; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4074 = _T_4072 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3563; // @[Reg.scala 27:20]
  wire  way_status_out_98 = _T_3563[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_532 = {{5'd0}, way_status_out_98}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4075 = _T_4074 & _GEN_532; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4068 = _GEN_473 == 7'h61; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4070 = _T_4068 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3559; // @[Reg.scala 27:20]
  wire  way_status_out_97 = _T_3559[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_534 = {{5'd0}, way_status_out_97}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4071 = _T_4070 & _GEN_534; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4064 = _GEN_473 == 7'h60; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4066 = _T_4064 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3555; // @[Reg.scala 27:20]
  wire  way_status_out_96 = _T_3555[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_536 = {{5'd0}, way_status_out_96}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4067 = _T_4066 & _GEN_536; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4060 = _GEN_473 == 7'h5f; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4062 = _T_4060 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3551; // @[Reg.scala 27:20]
  wire  way_status_out_95 = _T_3551[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_538 = {{5'd0}, way_status_out_95}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4063 = _T_4062 & _GEN_538; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4056 = _GEN_473 == 7'h5e; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4058 = _T_4056 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3547; // @[Reg.scala 27:20]
  wire  way_status_out_94 = _T_3547[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_540 = {{5'd0}, way_status_out_94}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4059 = _T_4058 & _GEN_540; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4052 = _GEN_473 == 7'h5d; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4054 = _T_4052 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3543; // @[Reg.scala 27:20]
  wire  way_status_out_93 = _T_3543[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_542 = {{5'd0}, way_status_out_93}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4055 = _T_4054 & _GEN_542; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4048 = _GEN_473 == 7'h5c; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4050 = _T_4048 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3539; // @[Reg.scala 27:20]
  wire  way_status_out_92 = _T_3539[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_544 = {{5'd0}, way_status_out_92}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4051 = _T_4050 & _GEN_544; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4044 = _GEN_473 == 7'h5b; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4046 = _T_4044 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3535; // @[Reg.scala 27:20]
  wire  way_status_out_91 = _T_3535[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_546 = {{5'd0}, way_status_out_91}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4047 = _T_4046 & _GEN_546; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [221:0] _T_4227 = {_T_4218,_T_4079,_T_4075,_T_4071,_T_4067,_T_4063,_T_4059,_T_4055,_T_4051,_T_4047}; // @[Cat.scala 29:58]
  wire  _T_4040 = _GEN_473 == 7'h5a; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4042 = _T_4040 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3531; // @[Reg.scala 27:20]
  wire  way_status_out_90 = _T_3531[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_548 = {{5'd0}, way_status_out_90}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4043 = _T_4042 & _GEN_548; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4036 = _GEN_473 == 7'h59; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4038 = _T_4036 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3527; // @[Reg.scala 27:20]
  wire  way_status_out_89 = _T_3527[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_550 = {{5'd0}, way_status_out_89}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4039 = _T_4038 & _GEN_550; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4032 = _GEN_473 == 7'h58; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4034 = _T_4032 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3523; // @[Reg.scala 27:20]
  wire  way_status_out_88 = _T_3523[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_552 = {{5'd0}, way_status_out_88}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4035 = _T_4034 & _GEN_552; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4028 = _GEN_473 == 7'h57; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4030 = _T_4028 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3519; // @[Reg.scala 27:20]
  wire  way_status_out_87 = _T_3519[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_554 = {{5'd0}, way_status_out_87}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4031 = _T_4030 & _GEN_554; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4024 = _GEN_473 == 7'h56; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4026 = _T_4024 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3515; // @[Reg.scala 27:20]
  wire  way_status_out_86 = _T_3515[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_556 = {{5'd0}, way_status_out_86}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4027 = _T_4026 & _GEN_556; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4020 = _GEN_473 == 7'h55; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4022 = _T_4020 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3511; // @[Reg.scala 27:20]
  wire  way_status_out_85 = _T_3511[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_558 = {{5'd0}, way_status_out_85}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4023 = _T_4022 & _GEN_558; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4016 = _GEN_473 == 7'h54; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4018 = _T_4016 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3507; // @[Reg.scala 27:20]
  wire  way_status_out_84 = _T_3507[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_560 = {{5'd0}, way_status_out_84}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4019 = _T_4018 & _GEN_560; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4012 = _GEN_473 == 7'h53; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4014 = _T_4012 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3503; // @[Reg.scala 27:20]
  wire  way_status_out_83 = _T_3503[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_562 = {{5'd0}, way_status_out_83}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4015 = _T_4014 & _GEN_562; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4008 = _GEN_473 == 7'h52; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4010 = _T_4008 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3499; // @[Reg.scala 27:20]
  wire  way_status_out_82 = _T_3499[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_564 = {{5'd0}, way_status_out_82}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4011 = _T_4010 & _GEN_564; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [275:0] _T_4236 = {_T_4227,_T_4043,_T_4039,_T_4035,_T_4031,_T_4027,_T_4023,_T_4019,_T_4015,_T_4011}; // @[Cat.scala 29:58]
  wire  _T_4004 = _GEN_473 == 7'h51; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4006 = _T_4004 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3495; // @[Reg.scala 27:20]
  wire  way_status_out_81 = _T_3495[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_566 = {{5'd0}, way_status_out_81}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4007 = _T_4006 & _GEN_566; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_4000 = _GEN_473 == 7'h50; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_4002 = _T_4000 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3491; // @[Reg.scala 27:20]
  wire  way_status_out_80 = _T_3491[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_568 = {{5'd0}, way_status_out_80}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_4003 = _T_4002 & _GEN_568; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3996 = _GEN_473 == 7'h4f; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3998 = _T_3996 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3487; // @[Reg.scala 27:20]
  wire  way_status_out_79 = _T_3487[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_570 = {{5'd0}, way_status_out_79}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3999 = _T_3998 & _GEN_570; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3992 = _GEN_473 == 7'h4e; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3994 = _T_3992 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3483; // @[Reg.scala 27:20]
  wire  way_status_out_78 = _T_3483[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_572 = {{5'd0}, way_status_out_78}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3995 = _T_3994 & _GEN_572; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3988 = _GEN_473 == 7'h4d; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3990 = _T_3988 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3479; // @[Reg.scala 27:20]
  wire  way_status_out_77 = _T_3479[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_574 = {{5'd0}, way_status_out_77}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3991 = _T_3990 & _GEN_574; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3984 = _GEN_473 == 7'h4c; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3986 = _T_3984 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3475; // @[Reg.scala 27:20]
  wire  way_status_out_76 = _T_3475[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_576 = {{5'd0}, way_status_out_76}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3987 = _T_3986 & _GEN_576; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3980 = _GEN_473 == 7'h4b; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3982 = _T_3980 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3471; // @[Reg.scala 27:20]
  wire  way_status_out_75 = _T_3471[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_578 = {{5'd0}, way_status_out_75}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3983 = _T_3982 & _GEN_578; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3976 = _GEN_473 == 7'h4a; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3978 = _T_3976 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3467; // @[Reg.scala 27:20]
  wire  way_status_out_74 = _T_3467[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_580 = {{5'd0}, way_status_out_74}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3979 = _T_3978 & _GEN_580; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3972 = _GEN_473 == 7'h49; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3974 = _T_3972 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3463; // @[Reg.scala 27:20]
  wire  way_status_out_73 = _T_3463[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_582 = {{5'd0}, way_status_out_73}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3975 = _T_3974 & _GEN_582; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [329:0] _T_4245 = {_T_4236,_T_4007,_T_4003,_T_3999,_T_3995,_T_3991,_T_3987,_T_3983,_T_3979,_T_3975}; // @[Cat.scala 29:58]
  wire  _T_3968 = _GEN_473 == 7'h48; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3970 = _T_3968 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3459; // @[Reg.scala 27:20]
  wire  way_status_out_72 = _T_3459[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_584 = {{5'd0}, way_status_out_72}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3971 = _T_3970 & _GEN_584; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3964 = _GEN_473 == 7'h47; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3966 = _T_3964 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3455; // @[Reg.scala 27:20]
  wire  way_status_out_71 = _T_3455[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_586 = {{5'd0}, way_status_out_71}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3967 = _T_3966 & _GEN_586; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3960 = _GEN_473 == 7'h46; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3962 = _T_3960 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3451; // @[Reg.scala 27:20]
  wire  way_status_out_70 = _T_3451[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_588 = {{5'd0}, way_status_out_70}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3963 = _T_3962 & _GEN_588; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3956 = _GEN_473 == 7'h45; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3958 = _T_3956 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3447; // @[Reg.scala 27:20]
  wire  way_status_out_69 = _T_3447[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_590 = {{5'd0}, way_status_out_69}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3959 = _T_3958 & _GEN_590; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3952 = _GEN_473 == 7'h44; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3954 = _T_3952 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3443; // @[Reg.scala 27:20]
  wire  way_status_out_68 = _T_3443[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_592 = {{5'd0}, way_status_out_68}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3955 = _T_3954 & _GEN_592; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3948 = _GEN_473 == 7'h43; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3950 = _T_3948 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3439; // @[Reg.scala 27:20]
  wire  way_status_out_67 = _T_3439[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_594 = {{5'd0}, way_status_out_67}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3951 = _T_3950 & _GEN_594; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3944 = _GEN_473 == 7'h42; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3946 = _T_3944 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3435; // @[Reg.scala 27:20]
  wire  way_status_out_66 = _T_3435[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_596 = {{5'd0}, way_status_out_66}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3947 = _T_3946 & _GEN_596; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3940 = _GEN_473 == 7'h41; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3942 = _T_3940 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3431; // @[Reg.scala 27:20]
  wire  way_status_out_65 = _T_3431[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_598 = {{5'd0}, way_status_out_65}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3943 = _T_3942 & _GEN_598; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3936 = _GEN_473 == 7'h40; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3938 = _T_3936 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3427; // @[Reg.scala 27:20]
  wire  way_status_out_64 = _T_3427[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_600 = {{5'd0}, way_status_out_64}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3939 = _T_3938 & _GEN_600; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [383:0] _T_4254 = {_T_4245,_T_3971,_T_3967,_T_3963,_T_3959,_T_3955,_T_3951,_T_3947,_T_3943,_T_3939}; // @[Cat.scala 29:58]
  wire  _T_3932 = ifu_ic_rw_int_addr_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3934 = _T_3932 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3423; // @[Reg.scala 27:20]
  wire  way_status_out_63 = _T_3423[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_601 = {{5'd0}, way_status_out_63}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3935 = _T_3934 & _GEN_601; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3928 = ifu_ic_rw_int_addr_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3930 = _T_3928 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3419; // @[Reg.scala 27:20]
  wire  way_status_out_62 = _T_3419[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_602 = {{5'd0}, way_status_out_62}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3931 = _T_3930 & _GEN_602; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3924 = ifu_ic_rw_int_addr_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3926 = _T_3924 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3415; // @[Reg.scala 27:20]
  wire  way_status_out_61 = _T_3415[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_603 = {{5'd0}, way_status_out_61}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3927 = _T_3926 & _GEN_603; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3920 = ifu_ic_rw_int_addr_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3922 = _T_3920 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3411; // @[Reg.scala 27:20]
  wire  way_status_out_60 = _T_3411[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_604 = {{5'd0}, way_status_out_60}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3923 = _T_3922 & _GEN_604; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3916 = ifu_ic_rw_int_addr_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3918 = _T_3916 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3407; // @[Reg.scala 27:20]
  wire  way_status_out_59 = _T_3407[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_605 = {{5'd0}, way_status_out_59}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3919 = _T_3918 & _GEN_605; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3912 = ifu_ic_rw_int_addr_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3914 = _T_3912 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3403; // @[Reg.scala 27:20]
  wire  way_status_out_58 = _T_3403[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_606 = {{5'd0}, way_status_out_58}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3915 = _T_3914 & _GEN_606; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3908 = ifu_ic_rw_int_addr_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3910 = _T_3908 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3399; // @[Reg.scala 27:20]
  wire  way_status_out_57 = _T_3399[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_607 = {{5'd0}, way_status_out_57}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3911 = _T_3910 & _GEN_607; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3904 = ifu_ic_rw_int_addr_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3906 = _T_3904 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3395; // @[Reg.scala 27:20]
  wire  way_status_out_56 = _T_3395[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_608 = {{5'd0}, way_status_out_56}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3907 = _T_3906 & _GEN_608; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3900 = ifu_ic_rw_int_addr_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3902 = _T_3900 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3391; // @[Reg.scala 27:20]
  wire  way_status_out_55 = _T_3391[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_609 = {{5'd0}, way_status_out_55}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3903 = _T_3902 & _GEN_609; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [437:0] _T_4263 = {_T_4254,_T_3935,_T_3931,_T_3927,_T_3923,_T_3919,_T_3915,_T_3911,_T_3907,_T_3903}; // @[Cat.scala 29:58]
  wire  _T_3896 = ifu_ic_rw_int_addr_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3898 = _T_3896 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3387; // @[Reg.scala 27:20]
  wire  way_status_out_54 = _T_3387[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_610 = {{5'd0}, way_status_out_54}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3899 = _T_3898 & _GEN_610; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3892 = ifu_ic_rw_int_addr_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3894 = _T_3892 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3383; // @[Reg.scala 27:20]
  wire  way_status_out_53 = _T_3383[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_611 = {{5'd0}, way_status_out_53}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3895 = _T_3894 & _GEN_611; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3888 = ifu_ic_rw_int_addr_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3890 = _T_3888 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3379; // @[Reg.scala 27:20]
  wire  way_status_out_52 = _T_3379[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_612 = {{5'd0}, way_status_out_52}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3891 = _T_3890 & _GEN_612; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3884 = ifu_ic_rw_int_addr_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3886 = _T_3884 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3375; // @[Reg.scala 27:20]
  wire  way_status_out_51 = _T_3375[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_613 = {{5'd0}, way_status_out_51}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3887 = _T_3886 & _GEN_613; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3880 = ifu_ic_rw_int_addr_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3882 = _T_3880 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3371; // @[Reg.scala 27:20]
  wire  way_status_out_50 = _T_3371[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_614 = {{5'd0}, way_status_out_50}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3883 = _T_3882 & _GEN_614; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3876 = ifu_ic_rw_int_addr_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3878 = _T_3876 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3367; // @[Reg.scala 27:20]
  wire  way_status_out_49 = _T_3367[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_615 = {{5'd0}, way_status_out_49}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3879 = _T_3878 & _GEN_615; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3872 = ifu_ic_rw_int_addr_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3874 = _T_3872 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3363; // @[Reg.scala 27:20]
  wire  way_status_out_48 = _T_3363[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_616 = {{5'd0}, way_status_out_48}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3875 = _T_3874 & _GEN_616; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3868 = ifu_ic_rw_int_addr_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3870 = _T_3868 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3359; // @[Reg.scala 27:20]
  wire  way_status_out_47 = _T_3359[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_617 = {{5'd0}, way_status_out_47}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3871 = _T_3870 & _GEN_617; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3864 = ifu_ic_rw_int_addr_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3866 = _T_3864 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3355; // @[Reg.scala 27:20]
  wire  way_status_out_46 = _T_3355[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_618 = {{5'd0}, way_status_out_46}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3867 = _T_3866 & _GEN_618; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [491:0] _T_4272 = {_T_4263,_T_3899,_T_3895,_T_3891,_T_3887,_T_3883,_T_3879,_T_3875,_T_3871,_T_3867}; // @[Cat.scala 29:58]
  wire  _T_3860 = ifu_ic_rw_int_addr_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3862 = _T_3860 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3351; // @[Reg.scala 27:20]
  wire  way_status_out_45 = _T_3351[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_619 = {{5'd0}, way_status_out_45}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3863 = _T_3862 & _GEN_619; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3856 = ifu_ic_rw_int_addr_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3858 = _T_3856 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3347; // @[Reg.scala 27:20]
  wire  way_status_out_44 = _T_3347[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_620 = {{5'd0}, way_status_out_44}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3859 = _T_3858 & _GEN_620; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3852 = ifu_ic_rw_int_addr_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3854 = _T_3852 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3343; // @[Reg.scala 27:20]
  wire  way_status_out_43 = _T_3343[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_621 = {{5'd0}, way_status_out_43}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3855 = _T_3854 & _GEN_621; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3848 = ifu_ic_rw_int_addr_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3850 = _T_3848 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3339; // @[Reg.scala 27:20]
  wire  way_status_out_42 = _T_3339[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_622 = {{5'd0}, way_status_out_42}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3851 = _T_3850 & _GEN_622; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3844 = ifu_ic_rw_int_addr_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3846 = _T_3844 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3335; // @[Reg.scala 27:20]
  wire  way_status_out_41 = _T_3335[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_623 = {{5'd0}, way_status_out_41}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3847 = _T_3846 & _GEN_623; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3840 = ifu_ic_rw_int_addr_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3842 = _T_3840 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3331; // @[Reg.scala 27:20]
  wire  way_status_out_40 = _T_3331[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_624 = {{5'd0}, way_status_out_40}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3843 = _T_3842 & _GEN_624; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3836 = ifu_ic_rw_int_addr_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3838 = _T_3836 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3327; // @[Reg.scala 27:20]
  wire  way_status_out_39 = _T_3327[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_625 = {{5'd0}, way_status_out_39}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3839 = _T_3838 & _GEN_625; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3832 = ifu_ic_rw_int_addr_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3834 = _T_3832 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3323; // @[Reg.scala 27:20]
  wire  way_status_out_38 = _T_3323[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_626 = {{5'd0}, way_status_out_38}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3835 = _T_3834 & _GEN_626; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3828 = ifu_ic_rw_int_addr_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3830 = _T_3828 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3319; // @[Reg.scala 27:20]
  wire  way_status_out_37 = _T_3319[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_627 = {{5'd0}, way_status_out_37}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3831 = _T_3830 & _GEN_627; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [545:0] _T_4281 = {_T_4272,_T_3863,_T_3859,_T_3855,_T_3851,_T_3847,_T_3843,_T_3839,_T_3835,_T_3831}; // @[Cat.scala 29:58]
  wire  _T_3824 = ifu_ic_rw_int_addr_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3826 = _T_3824 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3315; // @[Reg.scala 27:20]
  wire  way_status_out_36 = _T_3315[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_628 = {{5'd0}, way_status_out_36}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3827 = _T_3826 & _GEN_628; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3820 = ifu_ic_rw_int_addr_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3822 = _T_3820 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3311; // @[Reg.scala 27:20]
  wire  way_status_out_35 = _T_3311[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_629 = {{5'd0}, way_status_out_35}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3823 = _T_3822 & _GEN_629; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3816 = ifu_ic_rw_int_addr_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3818 = _T_3816 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3307; // @[Reg.scala 27:20]
  wire  way_status_out_34 = _T_3307[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_630 = {{5'd0}, way_status_out_34}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3819 = _T_3818 & _GEN_630; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3812 = ifu_ic_rw_int_addr_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3814 = _T_3812 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3303; // @[Reg.scala 27:20]
  wire  way_status_out_33 = _T_3303[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_631 = {{5'd0}, way_status_out_33}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3815 = _T_3814 & _GEN_631; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3808 = ifu_ic_rw_int_addr_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3810 = _T_3808 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3299; // @[Reg.scala 27:20]
  wire  way_status_out_32 = _T_3299[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_632 = {{5'd0}, way_status_out_32}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3811 = _T_3810 & _GEN_632; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3804 = ifu_ic_rw_int_addr_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3806 = _T_3804 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3295; // @[Reg.scala 27:20]
  wire  way_status_out_31 = _T_3295[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_633 = {{5'd0}, way_status_out_31}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3807 = _T_3806 & _GEN_633; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3800 = ifu_ic_rw_int_addr_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3802 = _T_3800 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3291; // @[Reg.scala 27:20]
  wire  way_status_out_30 = _T_3291[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_634 = {{5'd0}, way_status_out_30}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3803 = _T_3802 & _GEN_634; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3796 = ifu_ic_rw_int_addr_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3798 = _T_3796 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3287; // @[Reg.scala 27:20]
  wire  way_status_out_29 = _T_3287[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_635 = {{5'd0}, way_status_out_29}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3799 = _T_3798 & _GEN_635; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3792 = ifu_ic_rw_int_addr_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3794 = _T_3792 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3283; // @[Reg.scala 27:20]
  wire  way_status_out_28 = _T_3283[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_636 = {{5'd0}, way_status_out_28}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3795 = _T_3794 & _GEN_636; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [599:0] _T_4290 = {_T_4281,_T_3827,_T_3823,_T_3819,_T_3815,_T_3811,_T_3807,_T_3803,_T_3799,_T_3795}; // @[Cat.scala 29:58]
  wire  _T_3788 = ifu_ic_rw_int_addr_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3790 = _T_3788 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3279; // @[Reg.scala 27:20]
  wire  way_status_out_27 = _T_3279[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_637 = {{5'd0}, way_status_out_27}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3791 = _T_3790 & _GEN_637; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3784 = ifu_ic_rw_int_addr_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3786 = _T_3784 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3275; // @[Reg.scala 27:20]
  wire  way_status_out_26 = _T_3275[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_638 = {{5'd0}, way_status_out_26}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3787 = _T_3786 & _GEN_638; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3780 = ifu_ic_rw_int_addr_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3782 = _T_3780 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3271; // @[Reg.scala 27:20]
  wire  way_status_out_25 = _T_3271[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_639 = {{5'd0}, way_status_out_25}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3783 = _T_3782 & _GEN_639; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3776 = ifu_ic_rw_int_addr_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3778 = _T_3776 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3267; // @[Reg.scala 27:20]
  wire  way_status_out_24 = _T_3267[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_640 = {{5'd0}, way_status_out_24}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3779 = _T_3778 & _GEN_640; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3772 = ifu_ic_rw_int_addr_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3774 = _T_3772 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3263; // @[Reg.scala 27:20]
  wire  way_status_out_23 = _T_3263[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_641 = {{5'd0}, way_status_out_23}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3775 = _T_3774 & _GEN_641; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3768 = ifu_ic_rw_int_addr_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3770 = _T_3768 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3259; // @[Reg.scala 27:20]
  wire  way_status_out_22 = _T_3259[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_642 = {{5'd0}, way_status_out_22}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3771 = _T_3770 & _GEN_642; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3764 = ifu_ic_rw_int_addr_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3766 = _T_3764 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3255; // @[Reg.scala 27:20]
  wire  way_status_out_21 = _T_3255[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_643 = {{5'd0}, way_status_out_21}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3767 = _T_3766 & _GEN_643; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3760 = ifu_ic_rw_int_addr_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3762 = _T_3760 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3251; // @[Reg.scala 27:20]
  wire  way_status_out_20 = _T_3251[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_644 = {{5'd0}, way_status_out_20}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3763 = _T_3762 & _GEN_644; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3756 = ifu_ic_rw_int_addr_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3758 = _T_3756 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3247; // @[Reg.scala 27:20]
  wire  way_status_out_19 = _T_3247[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_645 = {{5'd0}, way_status_out_19}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3759 = _T_3758 & _GEN_645; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [653:0] _T_4299 = {_T_4290,_T_3791,_T_3787,_T_3783,_T_3779,_T_3775,_T_3771,_T_3767,_T_3763,_T_3759}; // @[Cat.scala 29:58]
  wire  _T_3752 = ifu_ic_rw_int_addr_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3754 = _T_3752 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3243; // @[Reg.scala 27:20]
  wire  way_status_out_18 = _T_3243[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_646 = {{5'd0}, way_status_out_18}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3755 = _T_3754 & _GEN_646; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3748 = ifu_ic_rw_int_addr_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3750 = _T_3748 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3239; // @[Reg.scala 27:20]
  wire  way_status_out_17 = _T_3239[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_647 = {{5'd0}, way_status_out_17}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3751 = _T_3750 & _GEN_647; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3744 = ifu_ic_rw_int_addr_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3746 = _T_3744 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3235; // @[Reg.scala 27:20]
  wire  way_status_out_16 = _T_3235[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_648 = {{5'd0}, way_status_out_16}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3747 = _T_3746 & _GEN_648; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3740 = ifu_ic_rw_int_addr_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3742 = _T_3740 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3231; // @[Reg.scala 27:20]
  wire  way_status_out_15 = _T_3231[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_649 = {{5'd0}, way_status_out_15}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3743 = _T_3742 & _GEN_649; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3736 = ifu_ic_rw_int_addr_ff == 6'he; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3738 = _T_3736 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3227; // @[Reg.scala 27:20]
  wire  way_status_out_14 = _T_3227[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_650 = {{5'd0}, way_status_out_14}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3739 = _T_3738 & _GEN_650; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3732 = ifu_ic_rw_int_addr_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3734 = _T_3732 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3223; // @[Reg.scala 27:20]
  wire  way_status_out_13 = _T_3223[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_651 = {{5'd0}, way_status_out_13}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3735 = _T_3734 & _GEN_651; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3728 = ifu_ic_rw_int_addr_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3730 = _T_3728 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3219; // @[Reg.scala 27:20]
  wire  way_status_out_12 = _T_3219[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_652 = {{5'd0}, way_status_out_12}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3731 = _T_3730 & _GEN_652; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3724 = ifu_ic_rw_int_addr_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3726 = _T_3724 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3215; // @[Reg.scala 27:20]
  wire  way_status_out_11 = _T_3215[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_653 = {{5'd0}, way_status_out_11}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3727 = _T_3726 & _GEN_653; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3720 = ifu_ic_rw_int_addr_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3722 = _T_3720 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3211; // @[Reg.scala 27:20]
  wire  way_status_out_10 = _T_3211[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_654 = {{5'd0}, way_status_out_10}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3723 = _T_3722 & _GEN_654; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [707:0] _T_4308 = {_T_4299,_T_3755,_T_3751,_T_3747,_T_3743,_T_3739,_T_3735,_T_3731,_T_3727,_T_3723}; // @[Cat.scala 29:58]
  wire  _T_3716 = ifu_ic_rw_int_addr_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3718 = _T_3716 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3207; // @[Reg.scala 27:20]
  wire  way_status_out_9 = _T_3207[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_655 = {{5'd0}, way_status_out_9}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3719 = _T_3718 & _GEN_655; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3712 = ifu_ic_rw_int_addr_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3714 = _T_3712 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3203; // @[Reg.scala 27:20]
  wire  way_status_out_8 = _T_3203[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_656 = {{5'd0}, way_status_out_8}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3715 = _T_3714 & _GEN_656; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3708 = ifu_ic_rw_int_addr_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3710 = _T_3708 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3199; // @[Reg.scala 27:20]
  wire  way_status_out_7 = _T_3199[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_657 = {{5'd0}, way_status_out_7}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3711 = _T_3710 & _GEN_657; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3704 = ifu_ic_rw_int_addr_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3706 = _T_3704 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3195; // @[Reg.scala 27:20]
  wire  way_status_out_6 = _T_3195[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_658 = {{5'd0}, way_status_out_6}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3707 = _T_3706 & _GEN_658; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3700 = ifu_ic_rw_int_addr_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3702 = _T_3700 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3191; // @[Reg.scala 27:20]
  wire  way_status_out_5 = _T_3191[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_659 = {{5'd0}, way_status_out_5}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3703 = _T_3702 & _GEN_659; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3696 = ifu_ic_rw_int_addr_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3698 = _T_3696 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3187; // @[Reg.scala 27:20]
  wire  way_status_out_4 = _T_3187[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_660 = {{5'd0}, way_status_out_4}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3699 = _T_3698 & _GEN_660; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3692 = ifu_ic_rw_int_addr_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3694 = _T_3692 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3183; // @[Reg.scala 27:20]
  wire  way_status_out_3 = _T_3183[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_661 = {{5'd0}, way_status_out_3}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3695 = _T_3694 & _GEN_661; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3688 = ifu_ic_rw_int_addr_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3690 = _T_3688 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3179; // @[Reg.scala 27:20]
  wire  way_status_out_2 = _T_3179[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_662 = {{5'd0}, way_status_out_2}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3691 = _T_3690 & _GEN_662; // @[el2_ifu_mem_ctl.scala 737:130]
  wire  _T_3684 = ifu_ic_rw_int_addr_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3686 = _T_3684 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3175; // @[Reg.scala 27:20]
  wire  way_status_out_1 = _T_3175[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_663 = {{5'd0}, way_status_out_1}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3687 = _T_3686 & _GEN_663; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [761:0] _T_4317 = {_T_4308,_T_3719,_T_3715,_T_3711,_T_3707,_T_3703,_T_3699,_T_3695,_T_3691,_T_3687}; // @[Cat.scala 29:58]
  wire  _T_3680 = ifu_ic_rw_int_addr_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 737:121]
  wire [5:0] _T_3682 = _T_3680 ? 6'h3f : 6'h0; // @[Bitwise.scala 72:12]
  reg [2:0] _T_3171; // @[Reg.scala 27:20]
  wire  way_status_out_0 = _T_3171[0]; // @[el2_ifu_mem_ctl.scala 734:30 el2_ifu_mem_ctl.scala 736:33]
  wire [5:0] _GEN_664 = {{5'd0}, way_status_out_0}; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [5:0] _T_3683 = _T_3682 & _GEN_664; // @[el2_ifu_mem_ctl.scala 737:130]
  wire [767:0] _T_4318 = {_T_4317,_T_3683}; // @[Cat.scala 29:58]
  wire  way_status = _T_4318[0]; // @[el2_ifu_mem_ctl.scala 737:16]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 266:96]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 270:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 275:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 280:59]
  wire  _T_214 = _T_212 | _T_1390; // @[el2_ifu_mem_ctl.scala 280:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 280:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 286:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 286:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 286:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 286:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 293:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 293:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 293:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 294:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 294:32]
  wire  _T_274 = imb_ff[12:6] == imb_scnd_ff[12:6]; // @[el2_ifu_mem_ctl.scala 297:75]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 297:127]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_1819 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 635:48]
  wire  _T_1820 = _T_1819 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 635:52]
  wire  bus_ifu_wr_data_error_ff = _T_1820 & miss_pending; // @[el2_ifu_mem_ctl.scala 635:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 379:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 378:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 297:145]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 297:143]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 300:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 300:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 301:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 320:30]
  wire  _T_9268 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 790:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 321:24]
  wire  _T_9270 = _T_9268 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:51]
  wire  _T_9272 = _T_9270 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 790:67]
  wire  _T_9274 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 790:86]
  wire  replace_way_mb_any_0 = _T_9272 | _T_9274; // @[el2_ifu_mem_ctl.scala 790:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_9277 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 791:50]
  wire  _T_9279 = _T_9277 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 791:66]
  wire  _T_9281 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 791:85]
  wire  _T_9283 = _T_9281 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 791:100]
  wire  replace_way_mb_any_1 = _T_9279 | _T_9283; // @[el2_ifu_mem_ctl.scala 791:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 305:110]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 309:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 309:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 310:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 309:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 309:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 311:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 319:23]
  wire  _T_313 = _T_1405 & flush_final_f; // @[el2_ifu_mem_ctl.scala 323:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 323:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 323:53]
  wire  _T_1397 = ~_T_1392; // @[el2_ifu_mem_ctl.scala 470:46]
  wire  _T_1398 = _T_1390 & _T_1397; // @[el2_ifu_mem_ctl.scala 470:44]
  wire  stream_miss_f = _T_1398 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 470:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 323:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 323:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 329:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_1390; // @[el2_ifu_mem_ctl.scala 331:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 331:82]
  wire  _T_1411 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 475:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_1411}; // @[Cat.scala 29:58]
  wire  _T_1412 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1436 = _T_1412 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_1415 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1437 = _T_1415 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_1444 = _T_1436 | _T_1437; // @[Mux.scala 27:72]
  wire  _T_1418 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1438 = _T_1418 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1444 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1421 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1439 = _T_1421 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1424 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1440 = _T_1424 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1427 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1441 = _T_1427 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1430 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1442 = _T_1430 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1433 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 476:81]
  wire  _T_1443 = _T_1433 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 477:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 335:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 335:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 632:61]
  wire  _T_1813 = ic_act_miss_f_delayed & _T_1406; // @[el2_ifu_mem_ctl.scala 633:53]
  wire  reset_tag_valid_for_miss = _T_1813 & _T_17; // @[el2_ifu_mem_ctl.scala 633:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 335:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 337:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 339:84]
  wire  _T_1807 = ~_T_1819; // @[el2_ifu_mem_ctl.scala 630:84]
  wire  _T_1808 = _T_100 & _T_1807; // @[el2_ifu_mem_ctl.scala 630:82]
  wire  bus_ifu_wr_en_ff_q = _T_1808 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 630:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 339:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 340:31]
  wire [6:0] ic_wr_ecc = m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 349:13]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] ic_miss_buff_ecc = m2_io_ecc_out; // @[el2_ifu_mem_ctl.scala 353:20]
  wire [3:0] _T_1452 = {ifu_bus_rid_ff[2:1],_T_1411,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1453 = _T_1452 == 4'h0; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_1500 = _T_1453 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1456 = _T_1452 == 4'h1; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_1501 = _T_1456 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1516 = _T_1500 | _T_1501; // @[Mux.scala 27:72]
  wire  _T_1459 = _T_1452 == 4'h2; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_1502 = _T_1459 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1517 = _T_1516 | _T_1502; // @[Mux.scala 27:72]
  wire  _T_1462 = _T_1452 == 4'h3; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_1503 = _T_1462 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1518 = _T_1517 | _T_1503; // @[Mux.scala 27:72]
  wire  _T_1465 = _T_1452 == 4'h4; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_1504 = _T_1465 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1519 = _T_1518 | _T_1504; // @[Mux.scala 27:72]
  wire  _T_1468 = _T_1452 == 4'h5; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_1505 = _T_1468 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1520 = _T_1519 | _T_1505; // @[Mux.scala 27:72]
  wire  _T_1471 = _T_1452 == 4'h6; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_1506 = _T_1471 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1521 = _T_1520 | _T_1506; // @[Mux.scala 27:72]
  wire  _T_1474 = _T_1452 == 4'h7; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_1507 = _T_1474 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1522 = _T_1521 | _T_1507; // @[Mux.scala 27:72]
  wire  _T_1477 = _T_1452 == 4'h8; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_1508 = _T_1477 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1523 = _T_1522 | _T_1508; // @[Mux.scala 27:72]
  wire  _T_1480 = _T_1452 == 4'h9; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_1509 = _T_1480 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1524 = _T_1523 | _T_1509; // @[Mux.scala 27:72]
  wire  _T_1483 = _T_1452 == 4'ha; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_1510 = _T_1483 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1525 = _T_1524 | _T_1510; // @[Mux.scala 27:72]
  wire  _T_1486 = _T_1452 == 4'hb; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_1511 = _T_1486 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1526 = _T_1525 | _T_1511; // @[Mux.scala 27:72]
  wire  _T_1489 = _T_1452 == 4'hc; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_1512 = _T_1489 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1527 = _T_1526 | _T_1512; // @[Mux.scala 27:72]
  wire  _T_1492 = _T_1452 == 4'hd; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_1513 = _T_1492 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1528 = _T_1527 | _T_1513; // @[Mux.scala 27:72]
  wire  _T_1495 = _T_1452 == 4'he; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_1514 = _T_1495 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1529 = _T_1528 | _T_1514; // @[Mux.scala 27:72]
  wire  _T_1498 = _T_1452 == 4'hf; // @[el2_ifu_mem_ctl.scala 478:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_1515 = _T_1498 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1530 = _T_1529 | _T_1515; // @[Mux.scala 27:72]
  wire [3:0] _T_1532 = {ifu_bus_rid_ff[2:1],_T_1411,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1533 = _T_1532 == 4'h0; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1580 = _T_1533 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1536 = _T_1532 == 4'h1; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1581 = _T_1536 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1596 = _T_1580 | _T_1581; // @[Mux.scala 27:72]
  wire  _T_1539 = _T_1532 == 4'h2; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1582 = _T_1539 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1597 = _T_1596 | _T_1582; // @[Mux.scala 27:72]
  wire  _T_1542 = _T_1532 == 4'h3; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1583 = _T_1542 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1598 = _T_1597 | _T_1583; // @[Mux.scala 27:72]
  wire  _T_1545 = _T_1532 == 4'h4; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1584 = _T_1545 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1599 = _T_1598 | _T_1584; // @[Mux.scala 27:72]
  wire  _T_1548 = _T_1532 == 4'h5; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1585 = _T_1548 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1600 = _T_1599 | _T_1585; // @[Mux.scala 27:72]
  wire  _T_1551 = _T_1532 == 4'h6; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1586 = _T_1551 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1601 = _T_1600 | _T_1586; // @[Mux.scala 27:72]
  wire  _T_1554 = _T_1532 == 4'h7; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1587 = _T_1554 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1602 = _T_1601 | _T_1587; // @[Mux.scala 27:72]
  wire  _T_1557 = _T_1532 == 4'h8; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1588 = _T_1557 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1603 = _T_1602 | _T_1588; // @[Mux.scala 27:72]
  wire  _T_1560 = _T_1532 == 4'h9; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1589 = _T_1560 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1604 = _T_1603 | _T_1589; // @[Mux.scala 27:72]
  wire  _T_1563 = _T_1532 == 4'ha; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1590 = _T_1563 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1605 = _T_1604 | _T_1590; // @[Mux.scala 27:72]
  wire  _T_1566 = _T_1532 == 4'hb; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1591 = _T_1566 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1606 = _T_1605 | _T_1591; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1532 == 4'hc; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1592 = _T_1569 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1607 = _T_1606 | _T_1592; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1532 == 4'hd; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1593 = _T_1572 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1608 = _T_1607 | _T_1593; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1532 == 4'he; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1594 = _T_1575 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1609 = _T_1608 | _T_1594; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1532 == 4'hf; // @[el2_ifu_mem_ctl.scala 479:66]
  wire [31:0] _T_1595 = _T_1578 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1610 = _T_1609 | _T_1595; // @[Mux.scala 27:72]
  wire [141:0] _T_391 = {ic_wr_ecc,ifu_bus_rdata_ff,ic_miss_buff_ecc,_T_1530,_T_1610}; // @[Cat.scala 29:58]
  wire [141:0] _T_394 = {ic_miss_buff_ecc,_T_1530,_T_1610,ic_wr_ecc,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_391 : _T_394; // @[el2_ifu_mem_ctl.scala 369:28]
  wire  _T_353 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 359:56]
  wire  _T_354 = _T_353 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 359:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 425:28]
  wire  _T_570 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 628:35]
  wire  _T_439 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_439; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_496 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 416:118]
  wire  _T_497 = ic_miss_buff_data_valid[0] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_497; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_593 = _T_570 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_573 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  _T_440 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_440; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_500 = ic_miss_buff_data_valid[1] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_500; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_594 = _T_573 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_601 = _T_593 | _T_594; // @[Mux.scala 27:72]
  wire  _T_576 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  _T_441 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_441; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_503 = ic_miss_buff_data_valid[2] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_503; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_595 = _T_576 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_602 = _T_601 | _T_595; // @[Mux.scala 27:72]
  wire  _T_579 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  _T_442 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_442; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_506 = ic_miss_buff_data_valid[3] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_506; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_596 = _T_579 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_603 = _T_602 | _T_596; // @[Mux.scala 27:72]
  wire  _T_582 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  _T_443 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_443; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_509 = ic_miss_buff_data_valid[4] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_509; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_597 = _T_582 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_604 = _T_603 | _T_597; // @[Mux.scala 27:72]
  wire  _T_585 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  _T_444 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_444; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_512 = ic_miss_buff_data_valid[5] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_512; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_598 = _T_585 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_605 = _T_604 | _T_598; // @[Mux.scala 27:72]
  wire  _T_588 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  _T_445 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_445; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_515 = ic_miss_buff_data_valid[6] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_515; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_599 = _T_588 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_606 = _T_605 | _T_599; // @[Mux.scala 27:72]
  wire  _T_591 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 427:114]
  wire  _T_446 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 410:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_446; // @[el2_ifu_mem_ctl.scala 410:73]
  wire  _T_518 = ic_miss_buff_data_valid[7] & _T_496; // @[el2_ifu_mem_ctl.scala 416:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_518; // @[el2_ifu_mem_ctl.scala 416:88]
  wire  _T_600 = _T_591 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_606 | _T_600; // @[Mux.scala 27:72]
  wire  _T_609 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 428:58]
  wire  _T_610 = bypass_valid_value_check & _T_609; // @[el2_ifu_mem_ctl.scala 428:56]
  wire  _T_612 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 428:77]
  wire  _T_613 = _T_610 & _T_612; // @[el2_ifu_mem_ctl.scala 428:75]
  wire  _T_618 = _T_610 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 429:75]
  wire  _T_619 = _T_613 | _T_618; // @[el2_ifu_mem_ctl.scala 428:95]
  wire  _T_621 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 430:56]
  wire  _T_624 = _T_621 & _T_612; // @[el2_ifu_mem_ctl.scala 430:74]
  wire  _T_625 = _T_619 | _T_624; // @[el2_ifu_mem_ctl.scala 429:94]
  wire  _T_629 = _T_621 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 431:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 426:70]
  wire  _T_630 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_646 = _T_630 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_632 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_647 = _T_632 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_654 = _T_646 | _T_647; // @[Mux.scala 27:72]
  wire  _T_634 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_648 = _T_634 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_655 = _T_654 | _T_648; // @[Mux.scala 27:72]
  wire  _T_636 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_649 = _T_636 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_656 = _T_655 | _T_649; // @[Mux.scala 27:72]
  wire  _T_638 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_650 = _T_638 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_657 = _T_656 | _T_650; // @[Mux.scala 27:72]
  wire  _T_640 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_651 = _T_640 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_658 = _T_657 | _T_651; // @[Mux.scala 27:72]
  wire  _T_642 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_652 = _T_642 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_659 = _T_658 | _T_652; // @[Mux.scala 27:72]
  wire  _T_644 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 431:132]
  wire  _T_653 = _T_644 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_660 = _T_659 | _T_653; // @[Mux.scala 27:72]
  wire  _T_662 = _T_629 & _T_660; // @[el2_ifu_mem_ctl.scala 431:69]
  wire  _T_663 = _T_625 | _T_662; // @[el2_ifu_mem_ctl.scala 430:94]
  wire [4:0] _GEN_665 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 432:95]
  wire  _T_666 = _GEN_665 == 5'h1f; // @[el2_ifu_mem_ctl.scala 432:95]
  wire  _T_667 = bypass_valid_value_check & _T_666; // @[el2_ifu_mem_ctl.scala 432:56]
  wire  bypass_data_ready_in = _T_663 | _T_667; // @[el2_ifu_mem_ctl.scala 431:181]
  wire  _T_668 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 436:53]
  wire  _T_669 = _T_668 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 436:73]
  wire  _T_671 = _T_669 & _T_317; // @[el2_ifu_mem_ctl.scala 436:96]
  wire  _T_673 = _T_671 & _T_58; // @[el2_ifu_mem_ctl.scala 436:118]
  wire  _T_675 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 437:73]
  wire  _T_677 = _T_675 & _T_317; // @[el2_ifu_mem_ctl.scala 437:96]
  wire  _T_679 = _T_677 & _T_58; // @[el2_ifu_mem_ctl.scala 437:118]
  wire  _T_680 = _T_673 | _T_679; // @[el2_ifu_mem_ctl.scala 436:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 439:58]
  wire  _T_681 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 438:54]
  wire  _T_682 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 438:76]
  wire  _T_683 = _T_681 & _T_682; // @[el2_ifu_mem_ctl.scala 438:74]
  wire  _T_685 = _T_683 & _T_317; // @[el2_ifu_mem_ctl.scala 438:96]
  wire  ic_crit_wd_rdy_new_in = _T_680 | _T_685; // @[el2_ifu_mem_ctl.scala 437:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 638:43]
  wire  _T_406 = ic_crit_wd_rdy | _T_1390; // @[el2_ifu_mem_ctl.scala 383:38]
  wire  _T_408 = _T_406 | _T_1406; // @[el2_ifu_mem_ctl.scala 383:64]
  wire  _T_409 = ~_T_408; // @[el2_ifu_mem_ctl.scala 383:21]
  wire  _T_410 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 383:98]
  wire  sel_ic_data = _T_409 & _T_410; // @[el2_ifu_mem_ctl.scala 383:96]
  wire  _T_1613 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 483:44]
  wire  _T_779 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 450:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 422:60]
  wire  _T_723 = _T_570 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_724 = _T_573 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_731 = _T_723 | _T_724; // @[Mux.scala 27:72]
  wire  _T_725 = _T_576 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_732 = _T_731 | _T_725; // @[Mux.scala 27:72]
  wire  _T_726 = _T_579 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_733 = _T_732 | _T_726; // @[Mux.scala 27:72]
  wire  _T_727 = _T_582 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_734 = _T_733 | _T_727; // @[Mux.scala 27:72]
  wire  _T_728 = _T_585 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_735 = _T_734 | _T_728; // @[Mux.scala 27:72]
  wire  _T_729 = _T_588 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_736 = _T_735 | _T_729; // @[Mux.scala 27:72]
  wire  _T_730 = _T_591 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_736 | _T_730; // @[Mux.scala 27:72]
  wire  _T_762 = _T_1323 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_763 = _T_1326 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_770 = _T_762 | _T_763; // @[Mux.scala 27:72]
  wire  _T_764 = _T_1329 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_771 = _T_770 | _T_764; // @[Mux.scala 27:72]
  wire  _T_765 = _T_1332 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_772 = _T_771 | _T_765; // @[Mux.scala 27:72]
  wire  _T_766 = _T_1335 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_773 = _T_772 | _T_766; // @[Mux.scala 27:72]
  wire  _T_767 = _T_1338 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_774 = _T_773 | _T_767; // @[Mux.scala 27:72]
  wire  _T_768 = _T_1341 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_775 = _T_774 | _T_768; // @[Mux.scala 27:72]
  wire  _T_769 = _T_1344 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_775 | _T_769; // @[Mux.scala 27:72]
  wire  _T_780 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 452:70]
  wire  ifu_byp_data_err_new = _T_779 ? ic_miss_buff_data_error_bypass : _T_780; // @[el2_ifu_mem_ctl.scala 450:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 394:42]
  wire  _T_1614 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 483:91]
  wire  _T_1615 = ~_T_1614; // @[el2_ifu_mem_ctl.scala 483:60]
  wire  ic_rd_parity_final_err = _T_1613 & _T_1615; // @[el2_ifu_mem_ctl.scala 483:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_8886 = _T_3680 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 765:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_8888 = _T_3684 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9141 = _T_8886 | _T_8888; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_8890 = _T_3688 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9142 = _T_9141 | _T_8890; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_8892 = _T_3692 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9143 = _T_9142 | _T_8892; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_8894 = _T_3696 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9144 = _T_9143 | _T_8894; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_8896 = _T_3700 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9145 = _T_9144 | _T_8896; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_8898 = _T_3704 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9146 = _T_9145 | _T_8898; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_8900 = _T_3708 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9147 = _T_9146 | _T_8900; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_8902 = _T_3712 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9148 = _T_9147 | _T_8902; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_8904 = _T_3716 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9149 = _T_9148 | _T_8904; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_8906 = _T_3720 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9150 = _T_9149 | _T_8906; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_8908 = _T_3724 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9151 = _T_9150 | _T_8908; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_8910 = _T_3728 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9152 = _T_9151 | _T_8910; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_8912 = _T_3732 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9153 = _T_9152 | _T_8912; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_8914 = _T_3736 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9154 = _T_9153 | _T_8914; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_8916 = _T_3740 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9155 = _T_9154 | _T_8916; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_8918 = _T_3744 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9156 = _T_9155 | _T_8918; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_8920 = _T_3748 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9157 = _T_9156 | _T_8920; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_8922 = _T_3752 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9158 = _T_9157 | _T_8922; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_8924 = _T_3756 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9159 = _T_9158 | _T_8924; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_8926 = _T_3760 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9160 = _T_9159 | _T_8926; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_8928 = _T_3764 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9161 = _T_9160 | _T_8928; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_8930 = _T_3768 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9162 = _T_9161 | _T_8930; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_8932 = _T_3772 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9163 = _T_9162 | _T_8932; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_8934 = _T_3776 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9164 = _T_9163 | _T_8934; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_8936 = _T_3780 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9165 = _T_9164 | _T_8936; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_8938 = _T_3784 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9166 = _T_9165 | _T_8938; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_8940 = _T_3788 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9167 = _T_9166 | _T_8940; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_8942 = _T_3792 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9168 = _T_9167 | _T_8942; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_8944 = _T_3796 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9169 = _T_9168 | _T_8944; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_8946 = _T_3800 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9170 = _T_9169 | _T_8946; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_8948 = _T_3804 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9171 = _T_9170 | _T_8948; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_8950 = _T_3808 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9172 = _T_9171 | _T_8950; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_8952 = _T_3812 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9173 = _T_9172 | _T_8952; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_8954 = _T_3816 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9174 = _T_9173 | _T_8954; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_8956 = _T_3820 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9175 = _T_9174 | _T_8956; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_8958 = _T_3824 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9176 = _T_9175 | _T_8958; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_8960 = _T_3828 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9177 = _T_9176 | _T_8960; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_8962 = _T_3832 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9178 = _T_9177 | _T_8962; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_8964 = _T_3836 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9179 = _T_9178 | _T_8964; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_8966 = _T_3840 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9180 = _T_9179 | _T_8966; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_8968 = _T_3844 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9181 = _T_9180 | _T_8968; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_8970 = _T_3848 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9182 = _T_9181 | _T_8970; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_8972 = _T_3852 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9183 = _T_9182 | _T_8972; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_8974 = _T_3856 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9184 = _T_9183 | _T_8974; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_8976 = _T_3860 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9185 = _T_9184 | _T_8976; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_8978 = _T_3864 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9186 = _T_9185 | _T_8978; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_8980 = _T_3868 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9187 = _T_9186 | _T_8980; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_8982 = _T_3872 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9188 = _T_9187 | _T_8982; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_8984 = _T_3876 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9189 = _T_9188 | _T_8984; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_8986 = _T_3880 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9190 = _T_9189 | _T_8986; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_8988 = _T_3884 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9191 = _T_9190 | _T_8988; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_8990 = _T_3888 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9192 = _T_9191 | _T_8990; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_8992 = _T_3892 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9193 = _T_9192 | _T_8992; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_8994 = _T_3896 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9194 = _T_9193 | _T_8994; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_8996 = _T_3900 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9195 = _T_9194 | _T_8996; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_8998 = _T_3904 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9196 = _T_9195 | _T_8998; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_9000 = _T_3908 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9197 = _T_9196 | _T_9000; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_9002 = _T_3912 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9198 = _T_9197 | _T_9002; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_9004 = _T_3916 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9199 = _T_9198 | _T_9004; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_9006 = _T_3920 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9200 = _T_9199 | _T_9006; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_9008 = _T_3924 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9201 = _T_9200 | _T_9008; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_9010 = _T_3928 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9202 = _T_9201 | _T_9010; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_9012 = _T_3932 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9203 = _T_9202 | _T_9012; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_9014 = _T_3936 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9204 = _T_9203 | _T_9014; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_9016 = _T_3940 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9205 = _T_9204 | _T_9016; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_9018 = _T_3944 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9206 = _T_9205 | _T_9018; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_9020 = _T_3948 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9207 = _T_9206 | _T_9020; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_9022 = _T_3952 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9208 = _T_9207 | _T_9022; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_9024 = _T_3956 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9209 = _T_9208 | _T_9024; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_9026 = _T_3960 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9210 = _T_9209 | _T_9026; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_9028 = _T_3964 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9211 = _T_9210 | _T_9028; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_9030 = _T_3968 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9212 = _T_9211 | _T_9030; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_9032 = _T_3972 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9213 = _T_9212 | _T_9032; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_9034 = _T_3976 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9214 = _T_9213 | _T_9034; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_9036 = _T_3980 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9215 = _T_9214 | _T_9036; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_9038 = _T_3984 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9216 = _T_9215 | _T_9038; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_9040 = _T_3988 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9217 = _T_9216 | _T_9040; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_9042 = _T_3992 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9218 = _T_9217 | _T_9042; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_9044 = _T_3996 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9219 = _T_9218 | _T_9044; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_9046 = _T_4000 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9220 = _T_9219 | _T_9046; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_9048 = _T_4004 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9221 = _T_9220 | _T_9048; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_9050 = _T_4008 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9222 = _T_9221 | _T_9050; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_9052 = _T_4012 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9223 = _T_9222 | _T_9052; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_9054 = _T_4016 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9224 = _T_9223 | _T_9054; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_9056 = _T_4020 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9225 = _T_9224 | _T_9056; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_9058 = _T_4024 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9226 = _T_9225 | _T_9058; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_9060 = _T_4028 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9227 = _T_9226 | _T_9060; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_9062 = _T_4032 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9228 = _T_9227 | _T_9062; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_9064 = _T_4036 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9229 = _T_9228 | _T_9064; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_9066 = _T_4040 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9230 = _T_9229 | _T_9066; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_9068 = _T_4044 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9231 = _T_9230 | _T_9068; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_9070 = _T_4048 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9232 = _T_9231 | _T_9070; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_9072 = _T_4052 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9233 = _T_9232 | _T_9072; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_9074 = _T_4056 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9234 = _T_9233 | _T_9074; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_9076 = _T_4060 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9235 = _T_9234 | _T_9076; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_9078 = _T_4064 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9236 = _T_9235 | _T_9078; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_9080 = _T_4068 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9237 = _T_9236 | _T_9080; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_9082 = _T_4072 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9238 = _T_9237 | _T_9082; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_9084 = _T_4076 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9239 = _T_9238 | _T_9084; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_9086 = _T_4080 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9240 = _T_9239 | _T_9086; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_9088 = _T_4084 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9241 = _T_9240 | _T_9088; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_9090 = _T_4088 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9242 = _T_9241 | _T_9090; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_9092 = _T_4092 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9243 = _T_9242 | _T_9092; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_9094 = _T_4096 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9244 = _T_9243 | _T_9094; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_9096 = _T_4100 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9245 = _T_9244 | _T_9096; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_9098 = _T_4104 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9246 = _T_9245 | _T_9098; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_9100 = _T_4108 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9247 = _T_9246 | _T_9100; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_9102 = _T_4112 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9248 = _T_9247 | _T_9102; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_9104 = _T_4116 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9249 = _T_9248 | _T_9104; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_9106 = _T_4120 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9250 = _T_9249 | _T_9106; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_9108 = _T_4124 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9251 = _T_9250 | _T_9108; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_9110 = _T_4128 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9252 = _T_9251 | _T_9110; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_9112 = _T_4132 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9253 = _T_9252 | _T_9112; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_9114 = _T_4136 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9254 = _T_9253 | _T_9114; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_9116 = _T_4140 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9255 = _T_9254 | _T_9116; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_9118 = _T_4144 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9256 = _T_9255 | _T_9118; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_9120 = _T_4148 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9257 = _T_9256 | _T_9120; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_9122 = _T_4152 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9258 = _T_9257 | _T_9122; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_9124 = _T_4156 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9259 = _T_9258 | _T_9124; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_9126 = _T_4160 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9260 = _T_9259 | _T_9126; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_9128 = _T_4164 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9261 = _T_9260 | _T_9128; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_9130 = _T_4168 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9262 = _T_9261 | _T_9130; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_9132 = _T_4172 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9263 = _T_9262 | _T_9132; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_9134 = _T_4176 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9264 = _T_9263 | _T_9134; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_9136 = _T_4180 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9265 = _T_9264 | _T_9136; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_9138 = _T_4184 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9266 = _T_9265 | _T_9138; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_9140 = _T_4188 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_9267 = _T_9266 | _T_9140; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_8503 = _T_3680 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 765:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_8505 = _T_3684 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8758 = _T_8503 | _T_8505; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_8507 = _T_3688 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8759 = _T_8758 | _T_8507; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_8509 = _T_3692 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8760 = _T_8759 | _T_8509; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_8511 = _T_3696 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8761 = _T_8760 | _T_8511; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_8513 = _T_3700 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8762 = _T_8761 | _T_8513; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_8515 = _T_3704 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8763 = _T_8762 | _T_8515; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_8517 = _T_3708 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8764 = _T_8763 | _T_8517; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_8519 = _T_3712 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8765 = _T_8764 | _T_8519; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_8521 = _T_3716 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8766 = _T_8765 | _T_8521; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_8523 = _T_3720 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8767 = _T_8766 | _T_8523; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_8525 = _T_3724 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8768 = _T_8767 | _T_8525; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_8527 = _T_3728 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8769 = _T_8768 | _T_8527; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_8529 = _T_3732 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8770 = _T_8769 | _T_8529; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_8531 = _T_3736 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8771 = _T_8770 | _T_8531; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_8533 = _T_3740 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8772 = _T_8771 | _T_8533; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_8535 = _T_3744 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8773 = _T_8772 | _T_8535; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_8537 = _T_3748 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8774 = _T_8773 | _T_8537; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_8539 = _T_3752 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8775 = _T_8774 | _T_8539; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_8541 = _T_3756 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8776 = _T_8775 | _T_8541; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_8543 = _T_3760 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8777 = _T_8776 | _T_8543; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_8545 = _T_3764 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8778 = _T_8777 | _T_8545; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_8547 = _T_3768 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8779 = _T_8778 | _T_8547; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_8549 = _T_3772 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8780 = _T_8779 | _T_8549; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_8551 = _T_3776 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8781 = _T_8780 | _T_8551; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_8553 = _T_3780 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8782 = _T_8781 | _T_8553; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_8555 = _T_3784 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8783 = _T_8782 | _T_8555; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_8557 = _T_3788 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8784 = _T_8783 | _T_8557; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_8559 = _T_3792 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8785 = _T_8784 | _T_8559; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_8561 = _T_3796 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8786 = _T_8785 | _T_8561; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_8563 = _T_3800 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8787 = _T_8786 | _T_8563; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_8565 = _T_3804 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8788 = _T_8787 | _T_8565; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_8567 = _T_3808 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8789 = _T_8788 | _T_8567; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_8569 = _T_3812 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8790 = _T_8789 | _T_8569; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_8571 = _T_3816 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8791 = _T_8790 | _T_8571; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_8573 = _T_3820 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8792 = _T_8791 | _T_8573; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_8575 = _T_3824 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8793 = _T_8792 | _T_8575; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_8577 = _T_3828 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8794 = _T_8793 | _T_8577; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_8579 = _T_3832 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8795 = _T_8794 | _T_8579; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_8581 = _T_3836 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8796 = _T_8795 | _T_8581; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_8583 = _T_3840 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8797 = _T_8796 | _T_8583; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_8585 = _T_3844 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8798 = _T_8797 | _T_8585; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_8587 = _T_3848 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8799 = _T_8798 | _T_8587; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_8589 = _T_3852 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8800 = _T_8799 | _T_8589; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_8591 = _T_3856 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8801 = _T_8800 | _T_8591; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_8593 = _T_3860 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8802 = _T_8801 | _T_8593; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_8595 = _T_3864 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8803 = _T_8802 | _T_8595; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_8597 = _T_3868 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8804 = _T_8803 | _T_8597; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_8599 = _T_3872 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8805 = _T_8804 | _T_8599; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_8601 = _T_3876 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8806 = _T_8805 | _T_8601; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_8603 = _T_3880 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8807 = _T_8806 | _T_8603; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_8605 = _T_3884 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8808 = _T_8807 | _T_8605; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_8607 = _T_3888 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8809 = _T_8808 | _T_8607; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_8609 = _T_3892 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8810 = _T_8809 | _T_8609; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_8611 = _T_3896 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8811 = _T_8810 | _T_8611; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_8613 = _T_3900 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8812 = _T_8811 | _T_8613; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_8615 = _T_3904 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8813 = _T_8812 | _T_8615; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_8617 = _T_3908 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8814 = _T_8813 | _T_8617; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_8619 = _T_3912 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8815 = _T_8814 | _T_8619; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_8621 = _T_3916 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8816 = _T_8815 | _T_8621; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_8623 = _T_3920 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8817 = _T_8816 | _T_8623; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_8625 = _T_3924 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8818 = _T_8817 | _T_8625; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_8627 = _T_3928 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8819 = _T_8818 | _T_8627; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_8629 = _T_3932 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8820 = _T_8819 | _T_8629; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_8631 = _T_3936 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8821 = _T_8820 | _T_8631; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_8633 = _T_3940 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8822 = _T_8821 | _T_8633; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_8635 = _T_3944 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8823 = _T_8822 | _T_8635; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_8637 = _T_3948 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8824 = _T_8823 | _T_8637; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_8639 = _T_3952 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8825 = _T_8824 | _T_8639; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_8641 = _T_3956 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8826 = _T_8825 | _T_8641; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_8643 = _T_3960 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8827 = _T_8826 | _T_8643; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_8645 = _T_3964 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8828 = _T_8827 | _T_8645; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_8647 = _T_3968 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8829 = _T_8828 | _T_8647; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_8649 = _T_3972 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8830 = _T_8829 | _T_8649; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_8651 = _T_3976 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8831 = _T_8830 | _T_8651; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_8653 = _T_3980 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8832 = _T_8831 | _T_8653; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_8655 = _T_3984 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8833 = _T_8832 | _T_8655; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_8657 = _T_3988 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8834 = _T_8833 | _T_8657; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_8659 = _T_3992 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8835 = _T_8834 | _T_8659; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_8661 = _T_3996 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8836 = _T_8835 | _T_8661; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_8663 = _T_4000 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8837 = _T_8836 | _T_8663; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_8665 = _T_4004 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8838 = _T_8837 | _T_8665; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_8667 = _T_4008 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8839 = _T_8838 | _T_8667; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_8669 = _T_4012 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8840 = _T_8839 | _T_8669; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_8671 = _T_4016 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8841 = _T_8840 | _T_8671; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_8673 = _T_4020 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8842 = _T_8841 | _T_8673; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_8675 = _T_4024 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8843 = _T_8842 | _T_8675; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_8677 = _T_4028 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8844 = _T_8843 | _T_8677; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_8679 = _T_4032 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8845 = _T_8844 | _T_8679; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_8681 = _T_4036 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8846 = _T_8845 | _T_8681; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_8683 = _T_4040 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8847 = _T_8846 | _T_8683; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_8685 = _T_4044 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8848 = _T_8847 | _T_8685; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_8687 = _T_4048 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8849 = _T_8848 | _T_8687; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_8689 = _T_4052 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8850 = _T_8849 | _T_8689; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_8691 = _T_4056 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8851 = _T_8850 | _T_8691; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_8693 = _T_4060 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8852 = _T_8851 | _T_8693; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_8695 = _T_4064 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8853 = _T_8852 | _T_8695; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_8697 = _T_4068 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8854 = _T_8853 | _T_8697; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_8699 = _T_4072 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8855 = _T_8854 | _T_8699; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_8701 = _T_4076 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8856 = _T_8855 | _T_8701; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_8703 = _T_4080 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8857 = _T_8856 | _T_8703; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_8705 = _T_4084 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8858 = _T_8857 | _T_8705; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_8707 = _T_4088 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8859 = _T_8858 | _T_8707; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_8709 = _T_4092 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8860 = _T_8859 | _T_8709; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_8711 = _T_4096 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8861 = _T_8860 | _T_8711; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_8713 = _T_4100 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8862 = _T_8861 | _T_8713; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_8715 = _T_4104 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8863 = _T_8862 | _T_8715; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_8717 = _T_4108 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8864 = _T_8863 | _T_8717; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_8719 = _T_4112 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8865 = _T_8864 | _T_8719; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_8721 = _T_4116 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8866 = _T_8865 | _T_8721; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_8723 = _T_4120 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8867 = _T_8866 | _T_8723; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_8725 = _T_4124 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8868 = _T_8867 | _T_8725; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_8727 = _T_4128 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8869 = _T_8868 | _T_8727; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_8729 = _T_4132 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8870 = _T_8869 | _T_8729; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_8731 = _T_4136 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8871 = _T_8870 | _T_8731; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_8733 = _T_4140 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8872 = _T_8871 | _T_8733; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_8735 = _T_4144 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8873 = _T_8872 | _T_8735; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_8737 = _T_4148 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8874 = _T_8873 | _T_8737; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_8739 = _T_4152 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8875 = _T_8874 | _T_8739; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_8741 = _T_4156 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8876 = _T_8875 | _T_8741; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_8743 = _T_4160 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8877 = _T_8876 | _T_8743; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_8745 = _T_4164 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8878 = _T_8877 | _T_8745; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_8747 = _T_4168 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8879 = _T_8878 | _T_8747; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_8749 = _T_4172 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8880 = _T_8879 | _T_8749; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_8751 = _T_4176 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8881 = _T_8880 | _T_8751; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_8753 = _T_4180 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8882 = _T_8881 | _T_8753; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_8755 = _T_4184 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8883 = _T_8882 | _T_8755; // @[el2_ifu_mem_ctl.scala 765:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_8757 = _T_4188 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 765:10]
  wire  _T_8884 = _T_8883 | _T_8757; // @[el2_ifu_mem_ctl.scala 765:91]
  wire [1:0] ic_tag_valid_unq = {_T_9267,_T_8884}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 838:54]
  wire [1:0] _T_9306 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_9307 = ic_debug_way_ff & _T_9306; // @[el2_ifu_mem_ctl.scala 819:67]
  wire [1:0] _T_9308 = ic_tag_valid_unq & _T_9307; // @[el2_ifu_mem_ctl.scala 819:48]
  wire  ic_debug_tag_val_rd_out = |_T_9308; // @[el2_ifu_mem_ctl.scala 819:115]
  wire [65:0] _T_365 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_366; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_1748; // @[el2_ifu_mem_ctl.scala 377:80]
  wire  _T_404 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 382:98]
  wire  sel_byp_data = _T_408 & _T_404; // @[el2_ifu_mem_ctl.scala 382:96]
  wire [63:0] _T_415 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_416 = _T_415 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 389:64]
  wire [63:0] _T_418 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_1270 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 458:31]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_784 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_832 = _T_784 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_787 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_833 = _T_787 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_848 = _T_832 | _T_833; // @[Mux.scala 27:72]
  wire  _T_790 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_834 = _T_790 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_849 = _T_848 | _T_834; // @[Mux.scala 27:72]
  wire  _T_793 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_835 = _T_793 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_850 = _T_849 | _T_835; // @[Mux.scala 27:72]
  wire  _T_796 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_836 = _T_796 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_851 = _T_850 | _T_836; // @[Mux.scala 27:72]
  wire  _T_799 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_837 = _T_799 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_852 = _T_851 | _T_837; // @[Mux.scala 27:72]
  wire  _T_802 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_838 = _T_802 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_853 = _T_852 | _T_838; // @[Mux.scala 27:72]
  wire  _T_805 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_839 = _T_805 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_854 = _T_853 | _T_839; // @[Mux.scala 27:72]
  wire  _T_808 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_840 = _T_808 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_855 = _T_854 | _T_840; // @[Mux.scala 27:72]
  wire  _T_811 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_841 = _T_811 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_856 = _T_855 | _T_841; // @[Mux.scala 27:72]
  wire  _T_814 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_842 = _T_814 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_857 = _T_856 | _T_842; // @[Mux.scala 27:72]
  wire  _T_817 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_843 = _T_817 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_858 = _T_857 | _T_843; // @[Mux.scala 27:72]
  wire  _T_820 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_844 = _T_820 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_859 = _T_858 | _T_844; // @[Mux.scala 27:72]
  wire  _T_823 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_845 = _T_823 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_860 = _T_859 | _T_845; // @[Mux.scala 27:72]
  wire  _T_826 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_846 = _T_826 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_861 = _T_860 | _T_846; // @[Mux.scala 27:72]
  wire  _T_829 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 455:73]
  wire [15:0] _T_847 = _T_829 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_862 = _T_861 | _T_847; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_864 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_912 = _T_864 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_867 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_913 = _T_867 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_928 = _T_912 | _T_913; // @[Mux.scala 27:72]
  wire  _T_870 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_914 = _T_870 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_929 = _T_928 | _T_914; // @[Mux.scala 27:72]
  wire  _T_873 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_915 = _T_873 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_930 = _T_929 | _T_915; // @[Mux.scala 27:72]
  wire  _T_876 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_916 = _T_876 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_931 = _T_930 | _T_916; // @[Mux.scala 27:72]
  wire  _T_879 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_917 = _T_879 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_932 = _T_931 | _T_917; // @[Mux.scala 27:72]
  wire  _T_882 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_918 = _T_882 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_933 = _T_932 | _T_918; // @[Mux.scala 27:72]
  wire  _T_885 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_919 = _T_885 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_934 = _T_933 | _T_919; // @[Mux.scala 27:72]
  wire  _T_888 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_920 = _T_888 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_935 = _T_934 | _T_920; // @[Mux.scala 27:72]
  wire  _T_891 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_921 = _T_891 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_936 = _T_935 | _T_921; // @[Mux.scala 27:72]
  wire  _T_894 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_922 = _T_894 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_937 = _T_936 | _T_922; // @[Mux.scala 27:72]
  wire  _T_897 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_923 = _T_897 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_938 = _T_937 | _T_923; // @[Mux.scala 27:72]
  wire  _T_900 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_924 = _T_900 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_939 = _T_938 | _T_924; // @[Mux.scala 27:72]
  wire  _T_903 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_925 = _T_903 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_940 = _T_939 | _T_925; // @[Mux.scala 27:72]
  wire  _T_906 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_926 = _T_906 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_941 = _T_940 | _T_926; // @[Mux.scala 27:72]
  wire  _T_909 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 455:179]
  wire [31:0] _T_927 = _T_909 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_942 = _T_941 | _T_927; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_944 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_992 = _T_944 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_947 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_993 = _T_947 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1008 = _T_992 | _T_993; // @[Mux.scala 27:72]
  wire  _T_950 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_994 = _T_950 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1009 = _T_1008 | _T_994; // @[Mux.scala 27:72]
  wire  _T_953 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_995 = _T_953 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1010 = _T_1009 | _T_995; // @[Mux.scala 27:72]
  wire  _T_956 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_996 = _T_956 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1011 = _T_1010 | _T_996; // @[Mux.scala 27:72]
  wire  _T_959 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_997 = _T_959 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1012 = _T_1011 | _T_997; // @[Mux.scala 27:72]
  wire  _T_962 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_998 = _T_962 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1013 = _T_1012 | _T_998; // @[Mux.scala 27:72]
  wire  _T_965 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_999 = _T_965 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1014 = _T_1013 | _T_999; // @[Mux.scala 27:72]
  wire  _T_968 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1000 = _T_968 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1015 = _T_1014 | _T_1000; // @[Mux.scala 27:72]
  wire  _T_971 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1001 = _T_971 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1016 = _T_1015 | _T_1001; // @[Mux.scala 27:72]
  wire  _T_974 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1002 = _T_974 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1017 = _T_1016 | _T_1002; // @[Mux.scala 27:72]
  wire  _T_977 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1003 = _T_977 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1018 = _T_1017 | _T_1003; // @[Mux.scala 27:72]
  wire  _T_980 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1004 = _T_980 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1019 = _T_1018 | _T_1004; // @[Mux.scala 27:72]
  wire  _T_983 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1005 = _T_983 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1020 = _T_1019 | _T_1005; // @[Mux.scala 27:72]
  wire  _T_986 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1006 = _T_986 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1021 = _T_1020 | _T_1006; // @[Mux.scala 27:72]
  wire  _T_989 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 455:285]
  wire [31:0] _T_1007 = _T_989 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1022 = _T_1021 | _T_1007; // @[Mux.scala 27:72]
  wire [79:0] _T_1025 = {_T_862,_T_942,_T_1022}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1026 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1074 = _T_1026 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1029 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1075 = _T_1029 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1090 = _T_1074 | _T_1075; // @[Mux.scala 27:72]
  wire  _T_1032 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1076 = _T_1032 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1091 = _T_1090 | _T_1076; // @[Mux.scala 27:72]
  wire  _T_1035 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1077 = _T_1035 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1092 = _T_1091 | _T_1077; // @[Mux.scala 27:72]
  wire  _T_1038 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1078 = _T_1038 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1093 = _T_1092 | _T_1078; // @[Mux.scala 27:72]
  wire  _T_1041 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1079 = _T_1041 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1094 = _T_1093 | _T_1079; // @[Mux.scala 27:72]
  wire  _T_1044 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1080 = _T_1044 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1095 = _T_1094 | _T_1080; // @[Mux.scala 27:72]
  wire  _T_1047 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1081 = _T_1047 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1096 = _T_1095 | _T_1081; // @[Mux.scala 27:72]
  wire  _T_1050 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1082 = _T_1050 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1097 = _T_1096 | _T_1082; // @[Mux.scala 27:72]
  wire  _T_1053 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1083 = _T_1053 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1098 = _T_1097 | _T_1083; // @[Mux.scala 27:72]
  wire  _T_1056 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1084 = _T_1056 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1099 = _T_1098 | _T_1084; // @[Mux.scala 27:72]
  wire  _T_1059 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1085 = _T_1059 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1100 = _T_1099 | _T_1085; // @[Mux.scala 27:72]
  wire  _T_1062 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1086 = _T_1062 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1101 = _T_1100 | _T_1086; // @[Mux.scala 27:72]
  wire  _T_1065 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1087 = _T_1065 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1102 = _T_1101 | _T_1087; // @[Mux.scala 27:72]
  wire  _T_1068 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1088 = _T_1068 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1103 = _T_1102 | _T_1088; // @[Mux.scala 27:72]
  wire  _T_1071 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 456:73]
  wire [15:0] _T_1089 = _T_1071 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1104 = _T_1103 | _T_1089; // @[Mux.scala 27:72]
  wire [31:0] _T_1154 = _T_784 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1155 = _T_787 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1170 = _T_1154 | _T_1155; // @[Mux.scala 27:72]
  wire [31:0] _T_1156 = _T_790 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1171 = _T_1170 | _T_1156; // @[Mux.scala 27:72]
  wire [31:0] _T_1157 = _T_793 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1172 = _T_1171 | _T_1157; // @[Mux.scala 27:72]
  wire [31:0] _T_1158 = _T_796 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1173 = _T_1172 | _T_1158; // @[Mux.scala 27:72]
  wire [31:0] _T_1159 = _T_799 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1174 = _T_1173 | _T_1159; // @[Mux.scala 27:72]
  wire [31:0] _T_1160 = _T_802 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1175 = _T_1174 | _T_1160; // @[Mux.scala 27:72]
  wire [31:0] _T_1161 = _T_805 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1176 = _T_1175 | _T_1161; // @[Mux.scala 27:72]
  wire [31:0] _T_1162 = _T_808 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1177 = _T_1176 | _T_1162; // @[Mux.scala 27:72]
  wire [31:0] _T_1163 = _T_811 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1178 = _T_1177 | _T_1163; // @[Mux.scala 27:72]
  wire [31:0] _T_1164 = _T_814 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1179 = _T_1178 | _T_1164; // @[Mux.scala 27:72]
  wire [31:0] _T_1165 = _T_817 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1180 = _T_1179 | _T_1165; // @[Mux.scala 27:72]
  wire [31:0] _T_1166 = _T_820 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1181 = _T_1180 | _T_1166; // @[Mux.scala 27:72]
  wire [31:0] _T_1167 = _T_823 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1182 = _T_1181 | _T_1167; // @[Mux.scala 27:72]
  wire [31:0] _T_1168 = _T_826 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1183 = _T_1182 | _T_1168; // @[Mux.scala 27:72]
  wire [31:0] _T_1169 = _T_829 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1184 = _T_1183 | _T_1169; // @[Mux.scala 27:72]
  wire [79:0] _T_1267 = {_T_1104,_T_1184,_T_942}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1270 ? _T_1025 : _T_1267; // @[el2_ifu_mem_ctl.scala 454:37]
  wire [79:0] _T_1272 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_1270 ? ic_byp_data_only_pre_new : _T_1272; // @[el2_ifu_mem_ctl.scala 458:30]
  wire [79:0] _GEN_794 = {{16'd0}, _T_418}; // @[el2_ifu_mem_ctl.scala 389:109]
  wire [79:0] _T_419 = _GEN_794 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 389:109]
  wire [79:0] _GEN_795 = {{16'd0}, _T_416}; // @[el2_ifu_mem_ctl.scala 389:83]
  wire [79:0] ic_premux_data = _GEN_795 | _T_419; // @[el2_ifu_mem_ctl.scala 389:83]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 396:38]
  wire [1:0] _T_428 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 400:8]
  wire [7:0] _T_525 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_530 = ic_miss_buff_data_error[0] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  _T_1816 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 634:47]
  wire  _T_1817 = _T_1816 & _T_13; // @[el2_ifu_mem_ctl.scala 634:50]
  wire  bus_ifu_wr_data_error = _T_1817 & miss_pending; // @[el2_ifu_mem_ctl.scala 634:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_530; // @[el2_ifu_mem_ctl.scala 420:72]
  wire  _T_534 = ic_miss_buff_data_error[1] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_534; // @[el2_ifu_mem_ctl.scala 420:72]
  wire  _T_538 = ic_miss_buff_data_error[2] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_538; // @[el2_ifu_mem_ctl.scala 420:72]
  wire  _T_542 = ic_miss_buff_data_error[3] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_542; // @[el2_ifu_mem_ctl.scala 420:72]
  wire  _T_546 = ic_miss_buff_data_error[4] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_546; // @[el2_ifu_mem_ctl.scala 420:72]
  wire  _T_550 = ic_miss_buff_data_error[5] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_550; // @[el2_ifu_mem_ctl.scala 420:72]
  wire  _T_554 = ic_miss_buff_data_error[6] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_554; // @[el2_ifu_mem_ctl.scala 420:72]
  wire  _T_558 = ic_miss_buff_data_error[7] & _T_496; // @[el2_ifu_mem_ctl.scala 421:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_558; // @[el2_ifu_mem_ctl.scala 420:72]
  wire [7:0] _T_565 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [5:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_1622 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1630 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 503:65]
  wire  _T_1631 = _T_1630 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 503:88]
  wire  _T_1633 = _T_1631 & _T_1744; // @[el2_ifu_mem_ctl.scala 503:112]
  wire  _T_1634 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1635 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 508:50]
  wire  _T_1637 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1643 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_1645 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_1643 | _T_1645; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_1637 ? _T_1635 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_1634 ? _T_1635 : _GEN_41; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_1622 ? _T_1633 : _GEN_43; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_1622 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_1636 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 509:56]
  wire  _GEN_44 = _T_1634 & _T_1636; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_1622 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 494:58]
  wire  _T_1619 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 493:49]
  wire  _T_1624 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 502:87]
  wire  _T_1638 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 512:54]
  wire  _T_1639 = _T_1638 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 512:84]
  wire  _T_1648 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 533:66]
  wire  _T_1649 = io_dec_tlu_flush_err_wb & _T_1648; // @[el2_ifu_mem_ctl.scala 533:52]
  wire  _T_1651 = _T_1649 & _T_1744; // @[el2_ifu_mem_ctl.scala 533:81]
  wire  _T_1653 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 536:59]
  wire  _T_1654 = _T_1653 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 536:86]
  wire  _T_1668 = _T_1653 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 539:81]
  wire  _T_1669 = _T_1668 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 539:103]
  wire  _T_1670 = _T_1669 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 539:126]
  wire  _T_1690 = _T_1668 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 546:103]
  wire  _T_1697 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 551:62]
  wire  _T_1698 = io_dec_tlu_flush_lower_wb & _T_1697; // @[el2_ifu_mem_ctl.scala 551:60]
  wire  _T_1699 = _T_1698 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 551:88]
  wire  _T_1700 = _T_1699 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 551:115]
  wire  _GEN_51 = _T_1696 & _T_1654; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_1679 ? _T_1690 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_1679 | _T_1696; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_1652 ? _T_1670 : _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_1652 | _GEN_56; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_1647 ? _T_1651 : _GEN_58; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_1712 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 568:64]
  wire  _T_1714 = _T_1712 & _T_1744; // @[el2_ifu_mem_ctl.scala 568:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_1716 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 568:133]
  wire  _T_1717 = _T_1716 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 568:164]
  wire  _T_1718 = _T_1717 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 568:184]
  wire  _T_1719 = _T_1718 & miss_pending; // @[el2_ifu_mem_ctl.scala 568:204]
  wire  _T_1720 = ~_T_1719; // @[el2_ifu_mem_ctl.scala 568:112]
  wire  ifc_bus_ic_req_ff_in = _T_1714 & _T_1720; // @[el2_ifu_mem_ctl.scala 568:110]
  wire  _T_1721 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 569:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 600:45]
  wire  _T_1738 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 603:35]
  wire  _T_1739 = _T_1738 & miss_pending; // @[el2_ifu_mem_ctl.scala 603:53]
  wire  bus_cmd_sent = _T_1739 & _T_1744; // @[el2_ifu_mem_ctl.scala 603:68]
  wire [2:0] _T_1729 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_1731 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1733 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 601:51]
  wire  _T_1759 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 611:73]
  wire  _T_1760 = _T_1745 & _T_1759; // @[el2_ifu_mem_ctl.scala 611:71]
  wire  _T_1762 = last_data_recieved_ff & _T_496; // @[el2_ifu_mem_ctl.scala 611:114]
  wire  last_data_recieved_in = _T_1760 | _T_1762; // @[el2_ifu_mem_ctl.scala 611:89]
  wire [2:0] _T_1768 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 616:45]
  wire  _T_1771 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 617:81]
  wire  _T_1772 = _T_1771 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 617:97]
  wire  _T_1774 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 619:48]
  wire  _T_1775 = _T_1774 & miss_pending; // @[el2_ifu_mem_ctl.scala 619:68]
  wire  bus_inc_cmd_beat_cnt = _T_1775 & _T_1744; // @[el2_ifu_mem_ctl.scala 619:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 621:57]
  wire  _T_1779 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 622:31]
  wire  _T_1780 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 622:71]
  wire  _T_1781 = _T_1780 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 622:87]
  wire  _T_1782 = ~_T_1781; // @[el2_ifu_mem_ctl.scala 622:55]
  wire  bus_hold_cmd_beat_cnt = _T_1779 & _T_1782; // @[el2_ifu_mem_ctl.scala 622:53]
  wire  _T_1783 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 623:46]
  wire  bus_cmd_beat_en = _T_1783 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 623:62]
  wire [2:0] _T_1786 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 625:46]
  wire [2:0] _T_1788 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1789 = bus_inc_cmd_beat_cnt ? _T_1786 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1790 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_1792 = _T_1788 | _T_1789; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_1792 | _T_1790; // @[Mux.scala 27:72]
  wire  _T_1796 = _T_1772 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 626:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 637:62]
  wire  _T_1824 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 642:50]
  wire  _T_1825 = io_ifc_dma_access_ok & _T_1824; // @[el2_ifu_mem_ctl.scala 642:47]
  wire  _T_1826 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 642:70]
  wire  ifc_dma_access_ok_d = _T_1825 & _T_1826; // @[el2_ifu_mem_ctl.scala 642:68]
  wire  _T_1830 = _T_1825 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 643:72]
  wire  _T_1831 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 643:111]
  wire  _T_1832 = _T_1830 & _T_1831; // @[el2_ifu_mem_ctl.scala 643:97]
  wire  ifc_dma_access_q_ok = _T_1832 & _T_1826; // @[el2_ifu_mem_ctl.scala 643:127]
  wire  _T_1835 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 646:40]
  wire  _T_1836 = _T_1835 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 646:58]
  wire  _T_1839 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 647:60]
  wire  _T_1840 = _T_1835 & _T_1839; // @[el2_ifu_mem_ctl.scala 647:58]
  wire  _T_1841 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 647:104]
  wire [2:0] _T_1846 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [8:0] _T_1952 = {io_dma_mem_wdata[48],io_dma_mem_wdata[46],io_dma_mem_wdata[44],io_dma_mem_wdata[42],io_dma_mem_wdata[40],io_dma_mem_wdata[38],io_dma_mem_wdata[37],io_dma_mem_wdata[35],io_dma_mem_wdata[33]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_1961 = {io_dma_mem_wdata[63],io_dma_mem_wdata[62],io_dma_mem_wdata[60],io_dma_mem_wdata[59],io_dma_mem_wdata[57],io_dma_mem_wdata[55],io_dma_mem_wdata[53],io_dma_mem_wdata[52],io_dma_mem_wdata[50],_T_1952}; // @[el2_lib.scala 268:22]
  wire  _T_1962 = ^_T_1961; // @[el2_lib.scala 268:29]
  wire [8:0] _T_1970 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_1979 = {io_dma_mem_wdata[63],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[51],io_dma_mem_wdata[50],_T_1970}; // @[el2_lib.scala 268:39]
  wire  _T_1980 = ^_T_1979; // @[el2_lib.scala 268:46]
  wire [8:0] _T_1988 = {io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_1997 = {io_dma_mem_wdata[62],io_dma_mem_wdata[61],io_dma_mem_wdata[60],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[49],io_dma_mem_wdata[48],_T_1988}; // @[el2_lib.scala 268:56]
  wire  _T_1998 = ^_T_1997; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2004 = {io_dma_mem_wdata[44],io_dma_mem_wdata[43],io_dma_mem_wdata[42],io_dma_mem_wdata[41],io_dma_mem_wdata[40],io_dma_mem_wdata[39],io_dma_mem_wdata[38]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2012 = {io_dma_mem_wdata[59],io_dma_mem_wdata[58],io_dma_mem_wdata[57],io_dma_mem_wdata[56],io_dma_mem_wdata[55],io_dma_mem_wdata[54],io_dma_mem_wdata[53],io_dma_mem_wdata[45],_T_2004}; // @[el2_lib.scala 268:73]
  wire  _T_2013 = ^_T_2012; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2027 = {io_dma_mem_wdata[52],io_dma_mem_wdata[51],io_dma_mem_wdata[50],io_dma_mem_wdata[49],io_dma_mem_wdata[48],io_dma_mem_wdata[47],io_dma_mem_wdata[46],io_dma_mem_wdata[45],_T_2004}; // @[el2_lib.scala 268:90]
  wire  _T_2028 = ^_T_2027; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2033 = {io_dma_mem_wdata[37],io_dma_mem_wdata[36],io_dma_mem_wdata[35],io_dma_mem_wdata[34],io_dma_mem_wdata[33],io_dma_mem_wdata[32]}; // @[el2_lib.scala 268:107]
  wire  _T_2034 = ^_T_2033; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2039 = {_T_1962,_T_1980,_T_1998,_T_2013,_T_2028,_T_2034}; // @[Cat.scala 29:58]
  wire  _T_2040 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 269:13]
  wire  _T_2041 = ^_T_2039; // @[el2_lib.scala 269:23]
  wire  _T_2042 = _T_2040 ^ _T_2041; // @[el2_lib.scala 269:18]
  wire [8:0] _T_2148 = {io_dma_mem_wdata[16],io_dma_mem_wdata[14],io_dma_mem_wdata[12],io_dma_mem_wdata[10],io_dma_mem_wdata[8],io_dma_mem_wdata[6],io_dma_mem_wdata[5],io_dma_mem_wdata[3],io_dma_mem_wdata[1]}; // @[el2_lib.scala 268:22]
  wire [17:0] _T_2157 = {io_dma_mem_wdata[31],io_dma_mem_wdata[30],io_dma_mem_wdata[28],io_dma_mem_wdata[27],io_dma_mem_wdata[25],io_dma_mem_wdata[23],io_dma_mem_wdata[21],io_dma_mem_wdata[20],io_dma_mem_wdata[18],_T_2148}; // @[el2_lib.scala 268:22]
  wire  _T_2158 = ^_T_2157; // @[el2_lib.scala 268:29]
  wire [8:0] _T_2166 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:39]
  wire [17:0] _T_2175 = {io_dma_mem_wdata[31],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[19],io_dma_mem_wdata[18],_T_2166}; // @[el2_lib.scala 268:39]
  wire  _T_2176 = ^_T_2175; // @[el2_lib.scala 268:46]
  wire [8:0] _T_2184 = {io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:56]
  wire [17:0] _T_2193 = {io_dma_mem_wdata[30],io_dma_mem_wdata[29],io_dma_mem_wdata[28],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[17],io_dma_mem_wdata[16],_T_2184}; // @[el2_lib.scala 268:56]
  wire  _T_2194 = ^_T_2193; // @[el2_lib.scala 268:63]
  wire [6:0] _T_2200 = {io_dma_mem_wdata[12],io_dma_mem_wdata[11],io_dma_mem_wdata[10],io_dma_mem_wdata[9],io_dma_mem_wdata[8],io_dma_mem_wdata[7],io_dma_mem_wdata[6]}; // @[el2_lib.scala 268:73]
  wire [14:0] _T_2208 = {io_dma_mem_wdata[27],io_dma_mem_wdata[26],io_dma_mem_wdata[25],io_dma_mem_wdata[24],io_dma_mem_wdata[23],io_dma_mem_wdata[22],io_dma_mem_wdata[21],io_dma_mem_wdata[13],_T_2200}; // @[el2_lib.scala 268:73]
  wire  _T_2209 = ^_T_2208; // @[el2_lib.scala 268:80]
  wire [14:0] _T_2223 = {io_dma_mem_wdata[20],io_dma_mem_wdata[19],io_dma_mem_wdata[18],io_dma_mem_wdata[17],io_dma_mem_wdata[16],io_dma_mem_wdata[15],io_dma_mem_wdata[14],io_dma_mem_wdata[13],_T_2200}; // @[el2_lib.scala 268:90]
  wire  _T_2224 = ^_T_2223; // @[el2_lib.scala 268:97]
  wire [5:0] _T_2229 = {io_dma_mem_wdata[5],io_dma_mem_wdata[4],io_dma_mem_wdata[3],io_dma_mem_wdata[2],io_dma_mem_wdata[1],io_dma_mem_wdata[0]}; // @[el2_lib.scala 268:107]
  wire  _T_2230 = ^_T_2229; // @[el2_lib.scala 268:114]
  wire [5:0] _T_2235 = {_T_2158,_T_2176,_T_2194,_T_2209,_T_2224,_T_2230}; // @[Cat.scala 29:58]
  wire  _T_2236 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 269:13]
  wire  _T_2237 = ^_T_2235; // @[el2_lib.scala 269:23]
  wire  _T_2238 = _T_2236 ^ _T_2237; // @[el2_lib.scala 269:18]
  wire [6:0] _T_2239 = {_T_2238,_T_2158,_T_2176,_T_2194,_T_2209,_T_2224,_T_2230}; // @[Cat.scala 29:58]
  wire [13:0] dma_mem_ecc = {_T_2042,_T_1962,_T_1980,_T_1998,_T_2013,_T_2028,_T_2034,_T_2239}; // @[Cat.scala 29:58]
  wire  _T_2241 = ~_T_1835; // @[el2_ifu_mem_ctl.scala 652:45]
  wire  _T_2242 = iccm_correct_ecc & _T_2241; // @[el2_ifu_mem_ctl.scala 652:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_2243 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_2250 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 666:53]
  wire  _T_2582 = _T_2494[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2580 = _T_2494[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2578 = _T_2494[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2576 = _T_2494[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2574 = _T_2494[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2572 = _T_2494[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2570 = _T_2494[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2568 = _T_2494[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2566 = _T_2494[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2564 = _T_2494[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2640 = {_T_2582,_T_2580,_T_2578,_T_2576,_T_2574,_T_2572,_T_2570,_T_2568,_T_2566,_T_2564}; // @[el2_lib.scala 310:69]
  wire  _T_2562 = _T_2494[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2560 = _T_2494[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2558 = _T_2494[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2556 = _T_2494[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2554 = _T_2494[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2552 = _T_2494[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2550 = _T_2494[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2548 = _T_2494[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2546 = _T_2494[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2544 = _T_2494[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2631 = {_T_2562,_T_2560,_T_2558,_T_2556,_T_2554,_T_2552,_T_2550,_T_2548,_T_2546,_T_2544}; // @[el2_lib.scala 310:69]
  wire  _T_2542 = _T_2494[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2540 = _T_2494[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2538 = _T_2494[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2536 = _T_2494[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2534 = _T_2494[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2532 = _T_2494[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2530 = _T_2494[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2528 = _T_2494[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2526 = _T_2494[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2524 = _T_2494[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_2621 = {_T_2542,_T_2540,_T_2538,_T_2536,_T_2534,_T_2532,_T_2530,_T_2528,_T_2526,_T_2524}; // @[el2_lib.scala 310:69]
  wire  _T_2522 = _T_2494[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2520 = _T_2494[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2518 = _T_2494[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2516 = _T_2494[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2514 = _T_2494[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2512 = _T_2494[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2510 = _T_2494[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2508 = _T_2494[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2506 = _T_2494[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_2622 = {_T_2621,_T_2522,_T_2520,_T_2518,_T_2516,_T_2514,_T_2512,_T_2510,_T_2508,_T_2506}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_2642 = {_T_2640,_T_2631,_T_2622}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2597 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2603 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_2597}; // @[Cat.scala 29:58]
  wire [38:0] _T_2643 = _T_2642 ^ _T_2603; // @[el2_lib.scala 310:76]
  wire [38:0] _T_2644 = _T_2498 ? _T_2643 : _T_2603; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_0 = {_T_2644[37:32],_T_2644[30:16],_T_2644[14:8],_T_2644[6:4],_T_2644[2]}; // @[Cat.scala 29:58]
  wire  _T_2967 = _T_2879[5:0] == 6'h27; // @[el2_lib.scala 307:41]
  wire  _T_2965 = _T_2879[5:0] == 6'h26; // @[el2_lib.scala 307:41]
  wire  _T_2963 = _T_2879[5:0] == 6'h25; // @[el2_lib.scala 307:41]
  wire  _T_2961 = _T_2879[5:0] == 6'h24; // @[el2_lib.scala 307:41]
  wire  _T_2959 = _T_2879[5:0] == 6'h23; // @[el2_lib.scala 307:41]
  wire  _T_2957 = _T_2879[5:0] == 6'h22; // @[el2_lib.scala 307:41]
  wire  _T_2955 = _T_2879[5:0] == 6'h21; // @[el2_lib.scala 307:41]
  wire  _T_2953 = _T_2879[5:0] == 6'h20; // @[el2_lib.scala 307:41]
  wire  _T_2951 = _T_2879[5:0] == 6'h1f; // @[el2_lib.scala 307:41]
  wire  _T_2949 = _T_2879[5:0] == 6'h1e; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3025 = {_T_2967,_T_2965,_T_2963,_T_2961,_T_2959,_T_2957,_T_2955,_T_2953,_T_2951,_T_2949}; // @[el2_lib.scala 310:69]
  wire  _T_2947 = _T_2879[5:0] == 6'h1d; // @[el2_lib.scala 307:41]
  wire  _T_2945 = _T_2879[5:0] == 6'h1c; // @[el2_lib.scala 307:41]
  wire  _T_2943 = _T_2879[5:0] == 6'h1b; // @[el2_lib.scala 307:41]
  wire  _T_2941 = _T_2879[5:0] == 6'h1a; // @[el2_lib.scala 307:41]
  wire  _T_2939 = _T_2879[5:0] == 6'h19; // @[el2_lib.scala 307:41]
  wire  _T_2937 = _T_2879[5:0] == 6'h18; // @[el2_lib.scala 307:41]
  wire  _T_2935 = _T_2879[5:0] == 6'h17; // @[el2_lib.scala 307:41]
  wire  _T_2933 = _T_2879[5:0] == 6'h16; // @[el2_lib.scala 307:41]
  wire  _T_2931 = _T_2879[5:0] == 6'h15; // @[el2_lib.scala 307:41]
  wire  _T_2929 = _T_2879[5:0] == 6'h14; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3016 = {_T_2947,_T_2945,_T_2943,_T_2941,_T_2939,_T_2937,_T_2935,_T_2933,_T_2931,_T_2929}; // @[el2_lib.scala 310:69]
  wire  _T_2927 = _T_2879[5:0] == 6'h13; // @[el2_lib.scala 307:41]
  wire  _T_2925 = _T_2879[5:0] == 6'h12; // @[el2_lib.scala 307:41]
  wire  _T_2923 = _T_2879[5:0] == 6'h11; // @[el2_lib.scala 307:41]
  wire  _T_2921 = _T_2879[5:0] == 6'h10; // @[el2_lib.scala 307:41]
  wire  _T_2919 = _T_2879[5:0] == 6'hf; // @[el2_lib.scala 307:41]
  wire  _T_2917 = _T_2879[5:0] == 6'he; // @[el2_lib.scala 307:41]
  wire  _T_2915 = _T_2879[5:0] == 6'hd; // @[el2_lib.scala 307:41]
  wire  _T_2913 = _T_2879[5:0] == 6'hc; // @[el2_lib.scala 307:41]
  wire  _T_2911 = _T_2879[5:0] == 6'hb; // @[el2_lib.scala 307:41]
  wire  _T_2909 = _T_2879[5:0] == 6'ha; // @[el2_lib.scala 307:41]
  wire [9:0] _T_3006 = {_T_2927,_T_2925,_T_2923,_T_2921,_T_2919,_T_2917,_T_2915,_T_2913,_T_2911,_T_2909}; // @[el2_lib.scala 310:69]
  wire  _T_2907 = _T_2879[5:0] == 6'h9; // @[el2_lib.scala 307:41]
  wire  _T_2905 = _T_2879[5:0] == 6'h8; // @[el2_lib.scala 307:41]
  wire  _T_2903 = _T_2879[5:0] == 6'h7; // @[el2_lib.scala 307:41]
  wire  _T_2901 = _T_2879[5:0] == 6'h6; // @[el2_lib.scala 307:41]
  wire  _T_2899 = _T_2879[5:0] == 6'h5; // @[el2_lib.scala 307:41]
  wire  _T_2897 = _T_2879[5:0] == 6'h4; // @[el2_lib.scala 307:41]
  wire  _T_2895 = _T_2879[5:0] == 6'h3; // @[el2_lib.scala 307:41]
  wire  _T_2893 = _T_2879[5:0] == 6'h2; // @[el2_lib.scala 307:41]
  wire  _T_2891 = _T_2879[5:0] == 6'h1; // @[el2_lib.scala 307:41]
  wire [18:0] _T_3007 = {_T_3006,_T_2907,_T_2905,_T_2903,_T_2901,_T_2899,_T_2897,_T_2895,_T_2893,_T_2891}; // @[el2_lib.scala 310:69]
  wire [38:0] _T_3027 = {_T_3025,_T_3016,_T_3007}; // @[el2_lib.scala 310:69]
  wire [7:0] _T_2982 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_2988 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_2982}; // @[Cat.scala 29:58]
  wire [38:0] _T_3028 = _T_3027 ^ _T_2988; // @[el2_lib.scala 310:76]
  wire [38:0] _T_3029 = _T_2883 ? _T_3028 : _T_2988; // @[el2_lib.scala 310:31]
  wire [31:0] iccm_corrected_data_1 = {_T_3029[37:32],_T_3029[30:16],_T_3029[14:8],_T_3029[6:4],_T_3029[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 658:35]
  wire  _T_2502 = ~_T_2494[6]; // @[el2_lib.scala 303:55]
  wire  _T_2503 = _T_2496 & _T_2502; // @[el2_lib.scala 303:53]
  wire  _T_2887 = ~_T_2879[6]; // @[el2_lib.scala 303:55]
  wire  _T_2888 = _T_2881 & _T_2887; // @[el2_lib.scala 303:53]
  wire [1:0] iccm_double_ecc_error = {_T_2503,_T_2888}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 660:53]
  wire [63:0] _T_2254 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_2255 = {iccm_dma_rdata_1_muxed,_T_2644[37:32],_T_2644[30:16],_T_2644[14:8],_T_2644[6:4],_T_2644[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 662:54]
  reg [2:0] iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 663:69]
  reg  iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 668:71]
  reg [63:0] iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 672:70]
  wire  _T_2260 = _T_1835 & _T_1824; // @[el2_ifu_mem_ctl.scala 675:65]
  wire  _T_2263 = _T_2241 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 676:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_2264 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_2266 = _T_2263 ? {{1'd0}, _T_2264} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 676:8]
  wire [31:0] _T_2267 = _T_2260 ? io_dma_mem_addr : {{16'd0}, _T_2266}; // @[el2_ifu_mem_ctl.scala 675:25]
  wire  _T_2656 = _T_2494 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_2657 = _T_2644[38] ^ _T_2656; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_2657,_T_2644[31],_T_2644[15],_T_2644[7],_T_2644[3],_T_2644[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3041 = _T_2879 == 7'h40; // @[el2_lib.scala 313:62]
  wire  _T_3042 = _T_3029[38] ^ _T_3041; // @[el2_lib.scala 313:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_3042,_T_3029[31],_T_3029[15],_T_3029[7],_T_3029[3],_T_3029[1:0]}; // @[Cat.scala 29:58]
  wire  _T_3058 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 688:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 690:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 691:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 699:62]
  wire  _T_3066 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 693:76]
  wire  _T_3067 = io_iccm_rd_ecc_single_err & _T_3066; // @[el2_ifu_mem_ctl.scala 693:74]
  wire  _T_3069 = _T_3067 & _T_317; // @[el2_ifu_mem_ctl.scala 693:104]
  wire  iccm_ecc_write_status = _T_3069 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 693:127]
  wire  _T_3070 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 694:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_3070 & _T_317; // @[el2_ifu_mem_ctl.scala 694:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 698:51]
  wire [13:0] _T_3075 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 697:102]
  wire [38:0] _T_3079 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_3084 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 702:41]
  wire  _T_3085 = io_ifc_fetch_req_bf & _T_3084; // @[el2_ifu_mem_ctl.scala 702:39]
  wire  _T_3086 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 702:72]
  wire  _T_3087 = _T_3085 & _T_3086; // @[el2_ifu_mem_ctl.scala 702:70]
  wire  _T_3089 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 703:34]
  wire  _T_3090 = _T_1390 & _T_3089; // @[el2_ifu_mem_ctl.scala 703:32]
  wire  _T_3093 = _T_1406 & _T_3089; // @[el2_ifu_mem_ctl.scala 704:37]
  wire  _T_3094 = _T_3090 | _T_3093; // @[el2_ifu_mem_ctl.scala 703:88]
  wire  _T_3095 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 705:19]
  wire  _T_3097 = _T_3095 & _T_3089; // @[el2_ifu_mem_ctl.scala 705:41]
  wire  _T_3098 = _T_3094 | _T_3097; // @[el2_ifu_mem_ctl.scala 704:88]
  wire  _T_3099 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 706:19]
  wire  _T_3101 = _T_3099 & _T_3089; // @[el2_ifu_mem_ctl.scala 706:35]
  wire  _T_3102 = _T_3098 | _T_3101; // @[el2_ifu_mem_ctl.scala 705:88]
  wire  _T_3105 = _T_1405 & _T_3089; // @[el2_ifu_mem_ctl.scala 707:38]
  wire  _T_3106 = _T_3102 | _T_3105; // @[el2_ifu_mem_ctl.scala 706:88]
  wire  _T_3108 = _T_1406 & miss_state_en; // @[el2_ifu_mem_ctl.scala 708:37]
  wire  _T_3109 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 708:71]
  wire  _T_3110 = _T_3108 & _T_3109; // @[el2_ifu_mem_ctl.scala 708:54]
  wire  _T_3111 = _T_3106 | _T_3110; // @[el2_ifu_mem_ctl.scala 707:57]
  wire  _T_3112 = ~_T_3111; // @[el2_ifu_mem_ctl.scala 703:5]
  wire  _T_3113 = _T_3087 & _T_3112; // @[el2_ifu_mem_ctl.scala 702:96]
  wire  _T_3114 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 709:28]
  wire  _T_3116 = _T_3114 & _T_3084; // @[el2_ifu_mem_ctl.scala 709:50]
  wire  _T_3118 = _T_3116 & _T_3086; // @[el2_ifu_mem_ctl.scala 709:81]
  wire  _T_3127 = ~_T_108; // @[el2_ifu_mem_ctl.scala 712:106]
  wire  _T_3128 = _T_1390 & _T_3127; // @[el2_ifu_mem_ctl.scala 712:104]
  wire  _T_3129 = _T_1406 | _T_3128; // @[el2_ifu_mem_ctl.scala 712:77]
  wire  _T_3133 = ~_T_51; // @[el2_ifu_mem_ctl.scala 712:172]
  wire  _T_3134 = _T_3129 & _T_3133; // @[el2_ifu_mem_ctl.scala 712:170]
  wire  _T_3135 = ~_T_3134; // @[el2_ifu_mem_ctl.scala 712:44]
  wire  _T_3139 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 715:64]
  wire  _T_3140 = ~_T_3139; // @[el2_ifu_mem_ctl.scala 715:50]
  wire  _T_3141 = _T_276 & _T_3140; // @[el2_ifu_mem_ctl.scala 715:48]
  wire  _T_3142 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 715:81]
  wire  ic_valid = _T_3141 & _T_3142; // @[el2_ifu_mem_ctl.scala 715:79]
  wire  _T_3144 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 716:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 719:14]
  wire  _T_3147 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 722:74]
  wire  _T_9289 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 796:45]
  wire  way_status_wr_en = _T_9289 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 796:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_3147; // @[el2_ifu_mem_ctl.scala 722:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 724:14]
  wire [2:0] _T_3151 = {{2'd0}, io_ic_debug_wr_data[4]}; // @[el2_ifu_mem_ctl.scala 728:10]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 792:41]
  wire  way_status_new = _T_9289 ? replace_way_mb_any_0 : way_status_hit_new; // @[el2_ifu_mem_ctl.scala 795:26]
  reg [2:0] way_status_new_ff; // @[el2_ifu_mem_ctl.scala 730:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 732:132]
  wire  _T_3168 = ifu_status_wr_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3169 = _T_3168 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3170 = _T_3169 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3172 = ifu_status_wr_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3173 = _T_3172 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3174 = _T_3173 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3176 = ifu_status_wr_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3177 = _T_3176 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3178 = _T_3177 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3180 = ifu_status_wr_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3181 = _T_3180 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3182 = _T_3181 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3184 = ifu_status_wr_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3185 = _T_3184 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3186 = _T_3185 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3188 = ifu_status_wr_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3189 = _T_3188 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3190 = _T_3189 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3192 = ifu_status_wr_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3193 = _T_3192 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3194 = _T_3193 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3196 = ifu_status_wr_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 736:93]
  wire  _T_3197 = _T_3196 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 736:102]
  wire  _T_3198 = _T_3197 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3202 = _T_3169 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3206 = _T_3173 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3210 = _T_3177 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3214 = _T_3181 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3218 = _T_3185 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3222 = _T_3189 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3226 = _T_3193 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3230 = _T_3197 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3234 = _T_3169 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3238 = _T_3173 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3242 = _T_3177 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3246 = _T_3181 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3250 = _T_3185 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3254 = _T_3189 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3258 = _T_3193 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3262 = _T_3197 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3266 = _T_3169 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3270 = _T_3173 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3274 = _T_3177 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3278 = _T_3181 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3282 = _T_3185 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3286 = _T_3189 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3290 = _T_3193 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3294 = _T_3197 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3298 = _T_3169 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3302 = _T_3173 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3306 = _T_3177 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3310 = _T_3181 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3314 = _T_3185 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3318 = _T_3189 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3322 = _T_3193 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3326 = _T_3197 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3330 = _T_3169 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3334 = _T_3173 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3338 = _T_3177 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3342 = _T_3181 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3346 = _T_3185 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3350 = _T_3189 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3354 = _T_3193 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3358 = _T_3197 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3362 = _T_3169 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3366 = _T_3173 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3370 = _T_3177 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3374 = _T_3181 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3378 = _T_3185 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3382 = _T_3189 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3386 = _T_3193 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3390 = _T_3197 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3394 = _T_3169 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3398 = _T_3173 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3402 = _T_3177 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3406 = _T_3181 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3410 = _T_3185 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3414 = _T_3189 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3418 = _T_3193 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3422 = _T_3197 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3426 = _T_3169 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3430 = _T_3173 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3434 = _T_3177 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3438 = _T_3181 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3442 = _T_3185 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3446 = _T_3189 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3450 = _T_3193 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3454 = _T_3197 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3458 = _T_3169 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3462 = _T_3173 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3466 = _T_3177 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3470 = _T_3181 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3474 = _T_3185 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3478 = _T_3189 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3482 = _T_3193 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3486 = _T_3197 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3490 = _T_3169 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3494 = _T_3173 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3498 = _T_3177 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3502 = _T_3181 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3506 = _T_3185 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3510 = _T_3189 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3514 = _T_3193 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3518 = _T_3197 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3522 = _T_3169 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3526 = _T_3173 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3530 = _T_3177 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3534 = _T_3181 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3538 = _T_3185 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3542 = _T_3189 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3546 = _T_3193 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3550 = _T_3197 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3554 = _T_3169 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3558 = _T_3173 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3562 = _T_3177 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3566 = _T_3181 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3570 = _T_3185 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3574 = _T_3189 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3578 = _T_3193 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3582 = _T_3197 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3586 = _T_3169 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3590 = _T_3173 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3594 = _T_3177 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3598 = _T_3181 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3602 = _T_3185 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3606 = _T_3189 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3610 = _T_3193 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3614 = _T_3197 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3618 = _T_3169 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3622 = _T_3173 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3626 = _T_3177 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3630 = _T_3181 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3634 = _T_3185 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3638 = _T_3189 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3642 = _T_3193 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3646 = _T_3197 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3650 = _T_3169 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3654 = _T_3173 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3658 = _T_3177 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3662 = _T_3181 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3666 = _T_3185 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3670 = _T_3189 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3674 = _T_3193 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_3678 = _T_3197 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 736:124]
  wire  _T_9295 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 799:84]
  wire  _T_9296 = _T_9295 & miss_pending; // @[el2_ifu_mem_ctl.scala 799:108]
  wire  bus_wren_last_1 = _T_9296 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 799:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 800:84]
  wire  _T_9298 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 801:73]
  wire  _T_9293 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 799:84]
  wire  _T_9294 = _T_9293 & miss_pending; // @[el2_ifu_mem_ctl.scala 799:108]
  wire  bus_wren_last_0 = _T_9294 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 799:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 800:84]
  wire  _T_9297 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 801:73]
  wire [1:0] ifu_tag_wren = {_T_9298,_T_9297}; // @[Cat.scala 29:58]
  wire [1:0] _T_9332 = _T_3147 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_9332 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 834:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 745:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 747:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 751:14]
  wire  _T_4327 = ifu_ic_rw_int_addr_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 755:82]
  wire  _T_4329 = _T_4327 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4331 = perr_ic_index_ff[5:4] == 2'h0; // @[el2_ifu_mem_ctl.scala 756:74]
  wire  _T_4333 = _T_4331 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4334 = _T_4329 | _T_4333; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4335 = _T_4334 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire  _T_4339 = _T_4327 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4343 = _T_4331 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4344 = _T_4339 | _T_4343; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4345 = _T_4344 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire [1:0] tag_valid_clken_0 = {_T_4335,_T_4345}; // @[Cat.scala 29:58]
  wire  _T_4347 = ifu_ic_rw_int_addr_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 755:82]
  wire  _T_4349 = _T_4347 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4351 = perr_ic_index_ff[5:4] == 2'h1; // @[el2_ifu_mem_ctl.scala 756:74]
  wire  _T_4353 = _T_4351 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4354 = _T_4349 | _T_4353; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4355 = _T_4354 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire  _T_4359 = _T_4347 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4363 = _T_4351 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4364 = _T_4359 | _T_4363; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4365 = _T_4364 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire [1:0] tag_valid_clken_1 = {_T_4355,_T_4365}; // @[Cat.scala 29:58]
  wire  _T_4367 = ifu_ic_rw_int_addr_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 755:82]
  wire  _T_4369 = _T_4367 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4371 = perr_ic_index_ff[5:4] == 2'h2; // @[el2_ifu_mem_ctl.scala 756:74]
  wire  _T_4373 = _T_4371 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4374 = _T_4369 | _T_4373; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4375 = _T_4374 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire  _T_4379 = _T_4367 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4383 = _T_4371 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4384 = _T_4379 | _T_4383; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4385 = _T_4384 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire [1:0] tag_valid_clken_2 = {_T_4375,_T_4385}; // @[Cat.scala 29:58]
  wire  _T_4387 = ifu_ic_rw_int_addr_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 755:82]
  wire  _T_4389 = _T_4387 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4391 = perr_ic_index_ff[5:4] == 2'h3; // @[el2_ifu_mem_ctl.scala 756:74]
  wire  _T_4393 = _T_4391 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4394 = _T_4389 | _T_4393; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4395 = _T_4394 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire  _T_4399 = _T_4387 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 755:91]
  wire  _T_4403 = _T_4391 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 756:83]
  wire  _T_4404 = _T_4399 | _T_4403; // @[el2_ifu_mem_ctl.scala 755:113]
  wire  _T_4405 = _T_4404 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 756:106]
  wire [1:0] tag_valid_clken_3 = {_T_4395,_T_4405}; // @[Cat.scala 29:58]
  wire  _T_4408 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 761:64]
  wire  _T_4409 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 761:91]
  wire  _T_4410 = _T_4408 & _T_4409; // @[el2_ifu_mem_ctl.scala 761:89]
  wire  _T_4413 = _T_3680 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4414 = perr_ic_index_ff == 6'h0; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4416 = _T_4414 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4418 = _T_4416 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4419 = _T_4413 | _T_4418; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4429 = _T_3684 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4430 = perr_ic_index_ff == 6'h1; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4432 = _T_4430 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4434 = _T_4432 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4435 = _T_4429 | _T_4434; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4445 = _T_3688 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4446 = perr_ic_index_ff == 6'h2; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4448 = _T_4446 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4450 = _T_4448 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4451 = _T_4445 | _T_4450; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4461 = _T_3692 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4462 = perr_ic_index_ff == 6'h3; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4464 = _T_4462 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4466 = _T_4464 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4467 = _T_4461 | _T_4466; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4477 = _T_3696 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4478 = perr_ic_index_ff == 6'h4; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4480 = _T_4478 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4482 = _T_4480 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4483 = _T_4477 | _T_4482; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4493 = _T_3700 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4494 = perr_ic_index_ff == 6'h5; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4496 = _T_4494 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4498 = _T_4496 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4499 = _T_4493 | _T_4498; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4509 = _T_3704 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4510 = perr_ic_index_ff == 6'h6; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4512 = _T_4510 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4514 = _T_4512 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4515 = _T_4509 | _T_4514; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4525 = _T_3708 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4526 = perr_ic_index_ff == 6'h7; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4528 = _T_4526 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4530 = _T_4528 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4531 = _T_4525 | _T_4530; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4541 = _T_3712 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4542 = perr_ic_index_ff == 6'h8; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4544 = _T_4542 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4546 = _T_4544 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4547 = _T_4541 | _T_4546; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4557 = _T_3716 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4558 = perr_ic_index_ff == 6'h9; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4560 = _T_4558 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4562 = _T_4560 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4563 = _T_4557 | _T_4562; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4573 = _T_3720 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4574 = perr_ic_index_ff == 6'ha; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4576 = _T_4574 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4578 = _T_4576 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4579 = _T_4573 | _T_4578; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4589 = _T_3724 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4590 = perr_ic_index_ff == 6'hb; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4592 = _T_4590 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4594 = _T_4592 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4595 = _T_4589 | _T_4594; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4605 = _T_3728 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4606 = perr_ic_index_ff == 6'hc; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4608 = _T_4606 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4610 = _T_4608 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4611 = _T_4605 | _T_4610; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4621 = _T_3732 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4622 = perr_ic_index_ff == 6'hd; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4624 = _T_4622 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4626 = _T_4624 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4627 = _T_4621 | _T_4626; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4637 = _T_3736 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4638 = perr_ic_index_ff == 6'he; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4640 = _T_4638 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4642 = _T_4640 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4643 = _T_4637 | _T_4642; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4653 = _T_3740 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4654 = perr_ic_index_ff == 6'hf; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4656 = _T_4654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4658 = _T_4656 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4659 = _T_4653 | _T_4658; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4669 = _T_3744 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4670 = perr_ic_index_ff == 6'h10; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4672 = _T_4670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4674 = _T_4672 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4675 = _T_4669 | _T_4674; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4685 = _T_3748 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4686 = perr_ic_index_ff == 6'h11; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4688 = _T_4686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4690 = _T_4688 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4691 = _T_4685 | _T_4690; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4701 = _T_3752 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4702 = perr_ic_index_ff == 6'h12; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4704 = _T_4702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4706 = _T_4704 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4707 = _T_4701 | _T_4706; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4717 = _T_3756 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4718 = perr_ic_index_ff == 6'h13; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4720 = _T_4718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4722 = _T_4720 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4723 = _T_4717 | _T_4722; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4733 = _T_3760 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4734 = perr_ic_index_ff == 6'h14; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4736 = _T_4734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4738 = _T_4736 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4739 = _T_4733 | _T_4738; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4749 = _T_3764 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4750 = perr_ic_index_ff == 6'h15; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4752 = _T_4750 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4754 = _T_4752 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4755 = _T_4749 | _T_4754; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4765 = _T_3768 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4766 = perr_ic_index_ff == 6'h16; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4768 = _T_4766 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4770 = _T_4768 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4771 = _T_4765 | _T_4770; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4781 = _T_3772 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4782 = perr_ic_index_ff == 6'h17; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4784 = _T_4782 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4786 = _T_4784 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4787 = _T_4781 | _T_4786; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4797 = _T_3776 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4798 = perr_ic_index_ff == 6'h18; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4800 = _T_4798 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4802 = _T_4800 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4803 = _T_4797 | _T_4802; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4813 = _T_3780 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4814 = perr_ic_index_ff == 6'h19; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4816 = _T_4814 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4818 = _T_4816 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4819 = _T_4813 | _T_4818; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4829 = _T_3784 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4830 = perr_ic_index_ff == 6'h1a; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4832 = _T_4830 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4834 = _T_4832 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4835 = _T_4829 | _T_4834; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4845 = _T_3788 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4846 = perr_ic_index_ff == 6'h1b; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4848 = _T_4846 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4850 = _T_4848 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4851 = _T_4845 | _T_4850; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4861 = _T_3792 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4862 = perr_ic_index_ff == 6'h1c; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4864 = _T_4862 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4866 = _T_4864 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4867 = _T_4861 | _T_4866; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4877 = _T_3796 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4878 = perr_ic_index_ff == 6'h1d; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4880 = _T_4878 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4882 = _T_4880 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4883 = _T_4877 | _T_4882; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4893 = _T_3800 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4894 = perr_ic_index_ff == 6'h1e; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4896 = _T_4894 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4898 = _T_4896 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4899 = _T_4893 | _T_4898; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4909 = _T_3804 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4910 = perr_ic_index_ff == 6'h1f; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_4912 = _T_4910 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4914 = _T_4912 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4915 = _T_4909 | _T_4914; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4925 = _T_3680 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4928 = _T_4414 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4930 = _T_4928 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4931 = _T_4925 | _T_4930; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4941 = _T_3684 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4944 = _T_4430 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4946 = _T_4944 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4947 = _T_4941 | _T_4946; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4957 = _T_3688 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4960 = _T_4446 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4962 = _T_4960 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4963 = _T_4957 | _T_4962; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4973 = _T_3692 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4976 = _T_4462 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4978 = _T_4976 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4979 = _T_4973 | _T_4978; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_4989 = _T_3696 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_4992 = _T_4478 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_4994 = _T_4992 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_4995 = _T_4989 | _T_4994; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5005 = _T_3700 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5008 = _T_4494 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5010 = _T_5008 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5011 = _T_5005 | _T_5010; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5021 = _T_3704 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5024 = _T_4510 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5026 = _T_5024 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5027 = _T_5021 | _T_5026; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5037 = _T_3708 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5040 = _T_4526 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5042 = _T_5040 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5043 = _T_5037 | _T_5042; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5053 = _T_3712 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5056 = _T_4542 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5058 = _T_5056 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5059 = _T_5053 | _T_5058; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5069 = _T_3716 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5072 = _T_4558 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5074 = _T_5072 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5075 = _T_5069 | _T_5074; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5085 = _T_3720 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5088 = _T_4574 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5090 = _T_5088 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5091 = _T_5085 | _T_5090; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5101 = _T_3724 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5104 = _T_4590 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5106 = _T_5104 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5107 = _T_5101 | _T_5106; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5117 = _T_3728 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5120 = _T_4606 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5122 = _T_5120 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5123 = _T_5117 | _T_5122; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5133 = _T_3732 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5136 = _T_4622 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5138 = _T_5136 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5139 = _T_5133 | _T_5138; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5149 = _T_3736 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5152 = _T_4638 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5154 = _T_5152 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5155 = _T_5149 | _T_5154; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5165 = _T_3740 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5168 = _T_4654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5170 = _T_5168 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5171 = _T_5165 | _T_5170; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5181 = _T_3744 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5184 = _T_4670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5186 = _T_5184 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5187 = _T_5181 | _T_5186; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5197 = _T_3748 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5200 = _T_4686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5202 = _T_5200 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5203 = _T_5197 | _T_5202; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5213 = _T_3752 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5216 = _T_4702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5218 = _T_5216 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5219 = _T_5213 | _T_5218; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5229 = _T_3756 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5232 = _T_4718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5234 = _T_5232 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5235 = _T_5229 | _T_5234; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5245 = _T_3760 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5248 = _T_4734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5250 = _T_5248 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5251 = _T_5245 | _T_5250; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5261 = _T_3764 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5264 = _T_4750 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5266 = _T_5264 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5267 = _T_5261 | _T_5266; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5277 = _T_3768 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5280 = _T_4766 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5282 = _T_5280 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5283 = _T_5277 | _T_5282; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5293 = _T_3772 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5296 = _T_4782 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5298 = _T_5296 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5299 = _T_5293 | _T_5298; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5309 = _T_3776 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5312 = _T_4798 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5314 = _T_5312 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5315 = _T_5309 | _T_5314; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5325 = _T_3780 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5328 = _T_4814 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5330 = _T_5328 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5331 = _T_5325 | _T_5330; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5341 = _T_3784 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5344 = _T_4830 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5346 = _T_5344 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5347 = _T_5341 | _T_5346; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5357 = _T_3788 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5360 = _T_4846 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5362 = _T_5360 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5363 = _T_5357 | _T_5362; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5373 = _T_3792 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5376 = _T_4862 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5378 = _T_5376 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5379 = _T_5373 | _T_5378; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5389 = _T_3796 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5392 = _T_4878 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5394 = _T_5392 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5395 = _T_5389 | _T_5394; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5405 = _T_3800 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5408 = _T_4894 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5410 = _T_5408 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5411 = _T_5405 | _T_5410; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5421 = _T_3804 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5424 = _T_4910 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5426 = _T_5424 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5427 = _T_5421 | _T_5426; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5437 = _T_3808 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5438 = perr_ic_index_ff == 6'h20; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5440 = _T_5438 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5442 = _T_5440 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5443 = _T_5437 | _T_5442; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5453 = _T_3812 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5454 = perr_ic_index_ff == 6'h21; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5456 = _T_5454 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5458 = _T_5456 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5459 = _T_5453 | _T_5458; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5469 = _T_3816 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5470 = perr_ic_index_ff == 6'h22; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5472 = _T_5470 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5474 = _T_5472 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5475 = _T_5469 | _T_5474; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5485 = _T_3820 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5486 = perr_ic_index_ff == 6'h23; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5488 = _T_5486 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5490 = _T_5488 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5491 = _T_5485 | _T_5490; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5501 = _T_3824 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5502 = perr_ic_index_ff == 6'h24; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5504 = _T_5502 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5506 = _T_5504 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5507 = _T_5501 | _T_5506; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5517 = _T_3828 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5518 = perr_ic_index_ff == 6'h25; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5520 = _T_5518 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5522 = _T_5520 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5523 = _T_5517 | _T_5522; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5533 = _T_3832 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5534 = perr_ic_index_ff == 6'h26; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5536 = _T_5534 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5538 = _T_5536 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5539 = _T_5533 | _T_5538; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5549 = _T_3836 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5550 = perr_ic_index_ff == 6'h27; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5552 = _T_5550 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5554 = _T_5552 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5555 = _T_5549 | _T_5554; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5565 = _T_3840 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5566 = perr_ic_index_ff == 6'h28; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5568 = _T_5566 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5570 = _T_5568 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5571 = _T_5565 | _T_5570; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5581 = _T_3844 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5582 = perr_ic_index_ff == 6'h29; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5584 = _T_5582 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5586 = _T_5584 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5587 = _T_5581 | _T_5586; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5597 = _T_3848 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5598 = perr_ic_index_ff == 6'h2a; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5600 = _T_5598 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5602 = _T_5600 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5603 = _T_5597 | _T_5602; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5613 = _T_3852 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5614 = perr_ic_index_ff == 6'h2b; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5616 = _T_5614 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5618 = _T_5616 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5619 = _T_5613 | _T_5618; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5629 = _T_3856 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5630 = perr_ic_index_ff == 6'h2c; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5632 = _T_5630 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5634 = _T_5632 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5635 = _T_5629 | _T_5634; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5645 = _T_3860 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5646 = perr_ic_index_ff == 6'h2d; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5648 = _T_5646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5650 = _T_5648 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5651 = _T_5645 | _T_5650; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5661 = _T_3864 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5662 = perr_ic_index_ff == 6'h2e; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5664 = _T_5662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5666 = _T_5664 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5667 = _T_5661 | _T_5666; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5677 = _T_3868 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5678 = perr_ic_index_ff == 6'h2f; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5680 = _T_5678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5682 = _T_5680 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5683 = _T_5677 | _T_5682; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5693 = _T_3872 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5694 = perr_ic_index_ff == 6'h30; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5696 = _T_5694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5698 = _T_5696 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5699 = _T_5693 | _T_5698; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5709 = _T_3876 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5710 = perr_ic_index_ff == 6'h31; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5712 = _T_5710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5714 = _T_5712 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5715 = _T_5709 | _T_5714; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5725 = _T_3880 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5726 = perr_ic_index_ff == 6'h32; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5728 = _T_5726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5730 = _T_5728 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5731 = _T_5725 | _T_5730; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5741 = _T_3884 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5742 = perr_ic_index_ff == 6'h33; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5744 = _T_5742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5746 = _T_5744 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5747 = _T_5741 | _T_5746; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5757 = _T_3888 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5758 = perr_ic_index_ff == 6'h34; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5760 = _T_5758 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5762 = _T_5760 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5763 = _T_5757 | _T_5762; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5773 = _T_3892 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5774 = perr_ic_index_ff == 6'h35; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5776 = _T_5774 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5778 = _T_5776 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5779 = _T_5773 | _T_5778; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5789 = _T_3896 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5790 = perr_ic_index_ff == 6'h36; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5792 = _T_5790 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5794 = _T_5792 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5795 = _T_5789 | _T_5794; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5805 = _T_3900 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5806 = perr_ic_index_ff == 6'h37; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5808 = _T_5806 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5810 = _T_5808 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5811 = _T_5805 | _T_5810; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5821 = _T_3904 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5822 = perr_ic_index_ff == 6'h38; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5824 = _T_5822 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5826 = _T_5824 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5827 = _T_5821 | _T_5826; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5837 = _T_3908 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5838 = perr_ic_index_ff == 6'h39; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5840 = _T_5838 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5842 = _T_5840 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5843 = _T_5837 | _T_5842; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5853 = _T_3912 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5854 = perr_ic_index_ff == 6'h3a; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5856 = _T_5854 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5858 = _T_5856 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5859 = _T_5853 | _T_5858; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5869 = _T_3916 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5870 = perr_ic_index_ff == 6'h3b; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5872 = _T_5870 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5874 = _T_5872 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5875 = _T_5869 | _T_5874; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5885 = _T_3920 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5886 = perr_ic_index_ff == 6'h3c; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5888 = _T_5886 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5890 = _T_5888 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5891 = _T_5885 | _T_5890; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5901 = _T_3924 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5902 = perr_ic_index_ff == 6'h3d; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5904 = _T_5902 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5906 = _T_5904 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5907 = _T_5901 | _T_5906; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5917 = _T_3928 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5918 = perr_ic_index_ff == 6'h3e; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5920 = _T_5918 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5922 = _T_5920 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5923 = _T_5917 | _T_5922; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5933 = _T_3932 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5934 = perr_ic_index_ff == 6'h3f; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_5936 = _T_5934 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5938 = _T_5936 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5939 = _T_5933 | _T_5938; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5949 = _T_3808 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5952 = _T_5438 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5954 = _T_5952 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5955 = _T_5949 | _T_5954; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5965 = _T_3812 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5968 = _T_5454 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5970 = _T_5968 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5971 = _T_5965 | _T_5970; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5981 = _T_3816 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_5984 = _T_5470 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_5986 = _T_5984 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_5987 = _T_5981 | _T_5986; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_5997 = _T_3820 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6000 = _T_5486 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6002 = _T_6000 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6003 = _T_5997 | _T_6002; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6013 = _T_3824 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6016 = _T_5502 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6018 = _T_6016 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6019 = _T_6013 | _T_6018; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6029 = _T_3828 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6032 = _T_5518 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6034 = _T_6032 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6035 = _T_6029 | _T_6034; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6045 = _T_3832 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6048 = _T_5534 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6050 = _T_6048 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6051 = _T_6045 | _T_6050; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6061 = _T_3836 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6064 = _T_5550 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6066 = _T_6064 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6067 = _T_6061 | _T_6066; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6077 = _T_3840 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6080 = _T_5566 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6082 = _T_6080 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6083 = _T_6077 | _T_6082; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6093 = _T_3844 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6096 = _T_5582 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6098 = _T_6096 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6099 = _T_6093 | _T_6098; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6109 = _T_3848 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6112 = _T_5598 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6114 = _T_6112 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6115 = _T_6109 | _T_6114; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6125 = _T_3852 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6128 = _T_5614 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6130 = _T_6128 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6131 = _T_6125 | _T_6130; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6141 = _T_3856 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6144 = _T_5630 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6146 = _T_6144 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6147 = _T_6141 | _T_6146; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6157 = _T_3860 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6160 = _T_5646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6162 = _T_6160 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6163 = _T_6157 | _T_6162; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6173 = _T_3864 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6176 = _T_5662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6178 = _T_6176 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6179 = _T_6173 | _T_6178; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6189 = _T_3868 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6192 = _T_5678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6194 = _T_6192 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6195 = _T_6189 | _T_6194; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6205 = _T_3872 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6208 = _T_5694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6210 = _T_6208 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6211 = _T_6205 | _T_6210; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6221 = _T_3876 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6224 = _T_5710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6226 = _T_6224 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6227 = _T_6221 | _T_6226; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6237 = _T_3880 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6240 = _T_5726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6242 = _T_6240 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6243 = _T_6237 | _T_6242; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6253 = _T_3884 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6256 = _T_5742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6258 = _T_6256 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6259 = _T_6253 | _T_6258; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6269 = _T_3888 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6272 = _T_5758 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6274 = _T_6272 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6275 = _T_6269 | _T_6274; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6285 = _T_3892 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6288 = _T_5774 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6290 = _T_6288 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6291 = _T_6285 | _T_6290; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6301 = _T_3896 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6304 = _T_5790 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6306 = _T_6304 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6307 = _T_6301 | _T_6306; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6317 = _T_3900 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6320 = _T_5806 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6322 = _T_6320 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6323 = _T_6317 | _T_6322; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6333 = _T_3904 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6336 = _T_5822 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6338 = _T_6336 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6339 = _T_6333 | _T_6338; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6349 = _T_3908 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6352 = _T_5838 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6354 = _T_6352 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6355 = _T_6349 | _T_6354; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6365 = _T_3912 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6368 = _T_5854 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6370 = _T_6368 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6371 = _T_6365 | _T_6370; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6381 = _T_3916 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6384 = _T_5870 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6386 = _T_6384 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6387 = _T_6381 | _T_6386; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6397 = _T_3920 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6400 = _T_5886 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6402 = _T_6400 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6403 = _T_6397 | _T_6402; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6413 = _T_3924 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6416 = _T_5902 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6418 = _T_6416 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6419 = _T_6413 | _T_6418; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6429 = _T_3928 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6432 = _T_5918 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6434 = _T_6432 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6435 = _T_6429 | _T_6434; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6445 = _T_3932 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6448 = _T_5934 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6450 = _T_6448 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6451 = _T_6445 | _T_6450; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6461 = _T_3936 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire [6:0] _GEN_797 = {{1'd0}, perr_ic_index_ff}; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6462 = _GEN_797 == 7'h40; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6464 = _T_6462 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6466 = _T_6464 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6467 = _T_6461 | _T_6466; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6477 = _T_3940 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6478 = _GEN_797 == 7'h41; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6480 = _T_6478 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6482 = _T_6480 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6483 = _T_6477 | _T_6482; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6493 = _T_3944 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6494 = _GEN_797 == 7'h42; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6496 = _T_6494 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6498 = _T_6496 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6499 = _T_6493 | _T_6498; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6509 = _T_3948 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6510 = _GEN_797 == 7'h43; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6512 = _T_6510 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6514 = _T_6512 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6515 = _T_6509 | _T_6514; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6525 = _T_3952 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6526 = _GEN_797 == 7'h44; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6528 = _T_6526 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6530 = _T_6528 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6531 = _T_6525 | _T_6530; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6541 = _T_3956 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6542 = _GEN_797 == 7'h45; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6544 = _T_6542 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6546 = _T_6544 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6547 = _T_6541 | _T_6546; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6557 = _T_3960 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6558 = _GEN_797 == 7'h46; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6560 = _T_6558 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6562 = _T_6560 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6563 = _T_6557 | _T_6562; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6573 = _T_3964 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6574 = _GEN_797 == 7'h47; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6576 = _T_6574 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6578 = _T_6576 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6579 = _T_6573 | _T_6578; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6589 = _T_3968 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6590 = _GEN_797 == 7'h48; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6592 = _T_6590 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6594 = _T_6592 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6595 = _T_6589 | _T_6594; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6605 = _T_3972 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6606 = _GEN_797 == 7'h49; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6608 = _T_6606 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6610 = _T_6608 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6611 = _T_6605 | _T_6610; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6621 = _T_3976 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6622 = _GEN_797 == 7'h4a; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6624 = _T_6622 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6626 = _T_6624 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6627 = _T_6621 | _T_6626; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6637 = _T_3980 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6638 = _GEN_797 == 7'h4b; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6640 = _T_6638 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6642 = _T_6640 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6643 = _T_6637 | _T_6642; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6653 = _T_3984 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6654 = _GEN_797 == 7'h4c; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6656 = _T_6654 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6658 = _T_6656 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6659 = _T_6653 | _T_6658; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6669 = _T_3988 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6670 = _GEN_797 == 7'h4d; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6672 = _T_6670 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6674 = _T_6672 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6675 = _T_6669 | _T_6674; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6685 = _T_3992 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6686 = _GEN_797 == 7'h4e; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6688 = _T_6686 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6690 = _T_6688 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6691 = _T_6685 | _T_6690; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6701 = _T_3996 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6702 = _GEN_797 == 7'h4f; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6704 = _T_6702 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6706 = _T_6704 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6707 = _T_6701 | _T_6706; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6717 = _T_4000 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6718 = _GEN_797 == 7'h50; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6720 = _T_6718 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6722 = _T_6720 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6723 = _T_6717 | _T_6722; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6733 = _T_4004 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6734 = _GEN_797 == 7'h51; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6736 = _T_6734 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6738 = _T_6736 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6739 = _T_6733 | _T_6738; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6749 = _T_4008 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6750 = _GEN_797 == 7'h52; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6752 = _T_6750 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6754 = _T_6752 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6755 = _T_6749 | _T_6754; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6765 = _T_4012 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6766 = _GEN_797 == 7'h53; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6768 = _T_6766 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6770 = _T_6768 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6771 = _T_6765 | _T_6770; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6781 = _T_4016 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6782 = _GEN_797 == 7'h54; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6784 = _T_6782 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6786 = _T_6784 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6787 = _T_6781 | _T_6786; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6797 = _T_4020 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6798 = _GEN_797 == 7'h55; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6800 = _T_6798 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6802 = _T_6800 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6803 = _T_6797 | _T_6802; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6813 = _T_4024 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6814 = _GEN_797 == 7'h56; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6816 = _T_6814 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6818 = _T_6816 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6819 = _T_6813 | _T_6818; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6829 = _T_4028 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6830 = _GEN_797 == 7'h57; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6832 = _T_6830 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6834 = _T_6832 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6835 = _T_6829 | _T_6834; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6845 = _T_4032 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6846 = _GEN_797 == 7'h58; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6848 = _T_6846 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6850 = _T_6848 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6851 = _T_6845 | _T_6850; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6861 = _T_4036 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6862 = _GEN_797 == 7'h59; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6864 = _T_6862 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6866 = _T_6864 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6867 = _T_6861 | _T_6866; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6877 = _T_4040 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6878 = _GEN_797 == 7'h5a; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6880 = _T_6878 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6882 = _T_6880 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6883 = _T_6877 | _T_6882; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6893 = _T_4044 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6894 = _GEN_797 == 7'h5b; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6896 = _T_6894 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6898 = _T_6896 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6899 = _T_6893 | _T_6898; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6909 = _T_4048 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6910 = _GEN_797 == 7'h5c; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6912 = _T_6910 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6914 = _T_6912 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6915 = _T_6909 | _T_6914; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6925 = _T_4052 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6926 = _GEN_797 == 7'h5d; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6928 = _T_6926 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6930 = _T_6928 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6931 = _T_6925 | _T_6930; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6941 = _T_4056 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6942 = _GEN_797 == 7'h5e; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6944 = _T_6942 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6946 = _T_6944 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6947 = _T_6941 | _T_6946; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6957 = _T_4060 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6958 = _GEN_797 == 7'h5f; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_6960 = _T_6958 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6962 = _T_6960 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6963 = _T_6957 | _T_6962; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6973 = _T_3936 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6976 = _T_6462 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6978 = _T_6976 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6979 = _T_6973 | _T_6978; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_6989 = _T_3940 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_6992 = _T_6478 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_6994 = _T_6992 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_6995 = _T_6989 | _T_6994; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7005 = _T_3944 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7008 = _T_6494 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7010 = _T_7008 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7011 = _T_7005 | _T_7010; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7021 = _T_3948 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7024 = _T_6510 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7026 = _T_7024 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7027 = _T_7021 | _T_7026; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7037 = _T_3952 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7040 = _T_6526 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7042 = _T_7040 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7043 = _T_7037 | _T_7042; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7053 = _T_3956 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7056 = _T_6542 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7058 = _T_7056 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7059 = _T_7053 | _T_7058; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7069 = _T_3960 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7072 = _T_6558 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7074 = _T_7072 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7075 = _T_7069 | _T_7074; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7085 = _T_3964 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7088 = _T_6574 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7090 = _T_7088 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7091 = _T_7085 | _T_7090; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7101 = _T_3968 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7104 = _T_6590 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7106 = _T_7104 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7107 = _T_7101 | _T_7106; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7117 = _T_3972 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7120 = _T_6606 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7122 = _T_7120 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7123 = _T_7117 | _T_7122; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7133 = _T_3976 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7136 = _T_6622 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7138 = _T_7136 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7139 = _T_7133 | _T_7138; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7149 = _T_3980 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7152 = _T_6638 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7154 = _T_7152 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7155 = _T_7149 | _T_7154; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7165 = _T_3984 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7168 = _T_6654 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7170 = _T_7168 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7171 = _T_7165 | _T_7170; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7181 = _T_3988 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7184 = _T_6670 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7186 = _T_7184 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7187 = _T_7181 | _T_7186; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7197 = _T_3992 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7200 = _T_6686 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7202 = _T_7200 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7203 = _T_7197 | _T_7202; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7213 = _T_3996 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7216 = _T_6702 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7218 = _T_7216 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7219 = _T_7213 | _T_7218; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7229 = _T_4000 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7232 = _T_6718 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7234 = _T_7232 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7235 = _T_7229 | _T_7234; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7245 = _T_4004 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7248 = _T_6734 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7250 = _T_7248 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7251 = _T_7245 | _T_7250; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7261 = _T_4008 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7264 = _T_6750 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7266 = _T_7264 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7267 = _T_7261 | _T_7266; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7277 = _T_4012 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7280 = _T_6766 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7282 = _T_7280 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7283 = _T_7277 | _T_7282; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7293 = _T_4016 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7296 = _T_6782 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7298 = _T_7296 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7299 = _T_7293 | _T_7298; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7309 = _T_4020 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7312 = _T_6798 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7314 = _T_7312 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7315 = _T_7309 | _T_7314; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7325 = _T_4024 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7328 = _T_6814 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7330 = _T_7328 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7331 = _T_7325 | _T_7330; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7341 = _T_4028 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7344 = _T_6830 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7346 = _T_7344 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7347 = _T_7341 | _T_7346; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7357 = _T_4032 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7360 = _T_6846 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7362 = _T_7360 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7363 = _T_7357 | _T_7362; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7373 = _T_4036 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7376 = _T_6862 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7378 = _T_7376 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7379 = _T_7373 | _T_7378; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7389 = _T_4040 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7392 = _T_6878 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7394 = _T_7392 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7395 = _T_7389 | _T_7394; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7405 = _T_4044 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7408 = _T_6894 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7410 = _T_7408 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7411 = _T_7405 | _T_7410; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7421 = _T_4048 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7424 = _T_6910 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7426 = _T_7424 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7427 = _T_7421 | _T_7426; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7437 = _T_4052 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7440 = _T_6926 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7442 = _T_7440 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7443 = _T_7437 | _T_7442; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7453 = _T_4056 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7456 = _T_6942 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7458 = _T_7456 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7459 = _T_7453 | _T_7458; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7469 = _T_4060 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7472 = _T_6958 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7474 = _T_7472 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7475 = _T_7469 | _T_7474; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7485 = _T_4064 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7486 = _GEN_797 == 7'h60; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7488 = _T_7486 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7490 = _T_7488 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7491 = _T_7485 | _T_7490; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7501 = _T_4068 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7502 = _GEN_797 == 7'h61; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7504 = _T_7502 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7506 = _T_7504 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7507 = _T_7501 | _T_7506; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7517 = _T_4072 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7518 = _GEN_797 == 7'h62; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7520 = _T_7518 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7522 = _T_7520 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7523 = _T_7517 | _T_7522; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7533 = _T_4076 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7534 = _GEN_797 == 7'h63; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7536 = _T_7534 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7538 = _T_7536 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7539 = _T_7533 | _T_7538; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7549 = _T_4080 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7550 = _GEN_797 == 7'h64; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7552 = _T_7550 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7554 = _T_7552 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7555 = _T_7549 | _T_7554; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7565 = _T_4084 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7566 = _GEN_797 == 7'h65; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7568 = _T_7566 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7570 = _T_7568 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7571 = _T_7565 | _T_7570; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7581 = _T_4088 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7582 = _GEN_797 == 7'h66; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7584 = _T_7582 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7586 = _T_7584 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7587 = _T_7581 | _T_7586; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7597 = _T_4092 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7598 = _GEN_797 == 7'h67; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7600 = _T_7598 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7602 = _T_7600 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7603 = _T_7597 | _T_7602; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7613 = _T_4096 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7614 = _GEN_797 == 7'h68; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7616 = _T_7614 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7618 = _T_7616 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7619 = _T_7613 | _T_7618; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7629 = _T_4100 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7630 = _GEN_797 == 7'h69; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7632 = _T_7630 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7634 = _T_7632 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7635 = _T_7629 | _T_7634; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7645 = _T_4104 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7646 = _GEN_797 == 7'h6a; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7648 = _T_7646 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7650 = _T_7648 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7651 = _T_7645 | _T_7650; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7661 = _T_4108 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7662 = _GEN_797 == 7'h6b; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7664 = _T_7662 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7666 = _T_7664 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7667 = _T_7661 | _T_7666; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7677 = _T_4112 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7678 = _GEN_797 == 7'h6c; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7680 = _T_7678 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7682 = _T_7680 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7683 = _T_7677 | _T_7682; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7693 = _T_4116 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7694 = _GEN_797 == 7'h6d; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7696 = _T_7694 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7698 = _T_7696 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7699 = _T_7693 | _T_7698; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7709 = _T_4120 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7710 = _GEN_797 == 7'h6e; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7712 = _T_7710 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7714 = _T_7712 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7715 = _T_7709 | _T_7714; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7725 = _T_4124 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7726 = _GEN_797 == 7'h6f; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7728 = _T_7726 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7730 = _T_7728 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7731 = _T_7725 | _T_7730; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7741 = _T_4128 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7742 = _GEN_797 == 7'h70; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7744 = _T_7742 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7746 = _T_7744 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7747 = _T_7741 | _T_7746; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7757 = _T_4132 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7758 = _GEN_797 == 7'h71; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7760 = _T_7758 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7762 = _T_7760 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7763 = _T_7757 | _T_7762; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7773 = _T_4136 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7774 = _GEN_797 == 7'h72; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7776 = _T_7774 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7778 = _T_7776 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7779 = _T_7773 | _T_7778; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7789 = _T_4140 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7790 = _GEN_797 == 7'h73; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7792 = _T_7790 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7794 = _T_7792 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7795 = _T_7789 | _T_7794; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7805 = _T_4144 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7806 = _GEN_797 == 7'h74; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7808 = _T_7806 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7810 = _T_7808 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7811 = _T_7805 | _T_7810; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7821 = _T_4148 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7822 = _GEN_797 == 7'h75; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7824 = _T_7822 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7826 = _T_7824 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7827 = _T_7821 | _T_7826; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7837 = _T_4152 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7838 = _GEN_797 == 7'h76; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7840 = _T_7838 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7842 = _T_7840 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7843 = _T_7837 | _T_7842; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7853 = _T_4156 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7854 = _GEN_797 == 7'h77; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7856 = _T_7854 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7858 = _T_7856 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7859 = _T_7853 | _T_7858; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7869 = _T_4160 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7870 = _GEN_797 == 7'h78; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7872 = _T_7870 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7874 = _T_7872 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7875 = _T_7869 | _T_7874; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7885 = _T_4164 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7886 = _GEN_797 == 7'h79; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7888 = _T_7886 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7890 = _T_7888 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7891 = _T_7885 | _T_7890; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7901 = _T_4168 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7902 = _GEN_797 == 7'h7a; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7904 = _T_7902 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7906 = _T_7904 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7907 = _T_7901 | _T_7906; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7917 = _T_4172 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7918 = _GEN_797 == 7'h7b; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7920 = _T_7918 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7922 = _T_7920 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7923 = _T_7917 | _T_7922; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7933 = _T_4176 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7934 = _GEN_797 == 7'h7c; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7936 = _T_7934 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7938 = _T_7936 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7939 = _T_7933 | _T_7938; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7949 = _T_4180 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7950 = _GEN_797 == 7'h7d; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7952 = _T_7950 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7954 = _T_7952 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7955 = _T_7949 | _T_7954; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7965 = _T_4184 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7966 = _GEN_797 == 7'h7e; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7968 = _T_7966 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7970 = _T_7968 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7971 = _T_7965 | _T_7970; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7981 = _T_4188 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_7982 = _GEN_797 == 7'h7f; // @[el2_ifu_mem_ctl.scala 762:101]
  wire  _T_7984 = _T_7982 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_7986 = _T_7984 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_7987 = _T_7981 | _T_7986; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_7997 = _T_4064 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8000 = _T_7486 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8002 = _T_8000 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8003 = _T_7997 | _T_8002; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8013 = _T_4068 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8016 = _T_7502 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8018 = _T_8016 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8019 = _T_8013 | _T_8018; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8029 = _T_4072 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8032 = _T_7518 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8034 = _T_8032 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8035 = _T_8029 | _T_8034; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8045 = _T_4076 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8048 = _T_7534 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8050 = _T_8048 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8051 = _T_8045 | _T_8050; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8061 = _T_4080 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8064 = _T_7550 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8066 = _T_8064 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8067 = _T_8061 | _T_8066; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8077 = _T_4084 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8080 = _T_7566 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8082 = _T_8080 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8083 = _T_8077 | _T_8082; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8093 = _T_4088 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8096 = _T_7582 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8098 = _T_8096 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8099 = _T_8093 | _T_8098; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8109 = _T_4092 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8112 = _T_7598 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8114 = _T_8112 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8115 = _T_8109 | _T_8114; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8125 = _T_4096 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8128 = _T_7614 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8130 = _T_8128 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8131 = _T_8125 | _T_8130; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8141 = _T_4100 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8144 = _T_7630 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8146 = _T_8144 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8147 = _T_8141 | _T_8146; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8157 = _T_4104 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8160 = _T_7646 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8162 = _T_8160 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8163 = _T_8157 | _T_8162; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8173 = _T_4108 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8176 = _T_7662 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8178 = _T_8176 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8179 = _T_8173 | _T_8178; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8189 = _T_4112 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8192 = _T_7678 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8194 = _T_8192 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8195 = _T_8189 | _T_8194; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8205 = _T_4116 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8208 = _T_7694 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8210 = _T_8208 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8211 = _T_8205 | _T_8210; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8221 = _T_4120 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8224 = _T_7710 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8226 = _T_8224 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8227 = _T_8221 | _T_8226; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8237 = _T_4124 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8240 = _T_7726 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8242 = _T_8240 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8243 = _T_8237 | _T_8242; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8253 = _T_4128 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8256 = _T_7742 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8258 = _T_8256 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8259 = _T_8253 | _T_8258; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8269 = _T_4132 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8272 = _T_7758 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8274 = _T_8272 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8275 = _T_8269 | _T_8274; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8285 = _T_4136 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8288 = _T_7774 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8290 = _T_8288 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8291 = _T_8285 | _T_8290; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8301 = _T_4140 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8304 = _T_7790 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8306 = _T_8304 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8307 = _T_8301 | _T_8306; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8317 = _T_4144 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8320 = _T_7806 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8322 = _T_8320 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8323 = _T_8317 | _T_8322; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8333 = _T_4148 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8336 = _T_7822 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8338 = _T_8336 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8339 = _T_8333 | _T_8338; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8349 = _T_4152 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8352 = _T_7838 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8354 = _T_8352 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8355 = _T_8349 | _T_8354; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8365 = _T_4156 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8368 = _T_7854 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8370 = _T_8368 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8371 = _T_8365 | _T_8370; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8381 = _T_4160 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8384 = _T_7870 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8386 = _T_8384 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8387 = _T_8381 | _T_8386; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8397 = _T_4164 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8400 = _T_7886 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8402 = _T_8400 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8403 = _T_8397 | _T_8402; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8413 = _T_4168 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8416 = _T_7902 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8418 = _T_8416 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8419 = _T_8413 | _T_8418; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8429 = _T_4172 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8432 = _T_7918 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8434 = _T_8432 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8435 = _T_8429 | _T_8434; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8445 = _T_4176 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8448 = _T_7934 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8450 = _T_8448 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8451 = _T_8445 | _T_8450; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8461 = _T_4180 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8464 = _T_7950 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8466 = _T_8464 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8467 = _T_8461 | _T_8466; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8477 = _T_4184 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8480 = _T_7966 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8482 = _T_8480 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8483 = _T_8477 | _T_8482; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_8493 = _T_4188 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:58]
  wire  _T_8496 = _T_7982 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 762:123]
  wire  _T_8498 = _T_8496 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 762:144]
  wire  _T_8499 = _T_8493 | _T_8498; // @[el2_ifu_mem_ctl.scala 762:80]
  wire  _T_9300 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 816:63]
  wire  _T_9301 = _T_9300 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 816:85]
  wire [1:0] _T_9303 = _T_9301 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_9310; // @[el2_ifu_mem_ctl.scala 821:57]
  reg  _T_9311; // @[el2_ifu_mem_ctl.scala 822:56]
  reg  _T_9312; // @[el2_ifu_mem_ctl.scala 823:59]
  wire  _T_9313 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 824:80]
  wire  _T_9314 = ifu_bus_arvalid_ff & _T_9313; // @[el2_ifu_mem_ctl.scala 824:78]
  wire  _T_9315 = _T_9314 & miss_pending; // @[el2_ifu_mem_ctl.scala 824:100]
  reg  _T_9316; // @[el2_ifu_mem_ctl.scala 824:58]
  reg  _T_9317; // @[el2_ifu_mem_ctl.scala 825:58]
  wire  _T_9320 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 832:71]
  wire  _T_9322 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 832:124]
  wire  _T_9324 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 833:50]
  wire  _T_9326 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 833:103]
  wire [3:0] _T_9329 = {_T_9320,_T_9322,_T_9324,_T_9326}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 835:53]
  reg  _T_9340; // @[Reg.scala 27:20]
  rvecc_encode_64 m1 ( // @[el2_ifu_mem_ctl.scala 346:18]
    .io_din(m1_io_din),
    .io_ecc_out(m1_io_ecc_out)
  );
  rvecc_encode_64 m2 ( // @[el2_ifu_mem_ctl.scala 347:18]
    .io_din(m2_io_din),
    .io_ecc_out(m2_io_ecc_out)
  );
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 332:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 331:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 195:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_3135; // @[el2_ifu_mem_ctl.scala 712:21]
  assign io_ifu_pmu_ic_miss = _T_9310; // @[el2_ifu_mem_ctl.scala 821:22]
  assign io_ifu_pmu_ic_hit = _T_9311; // @[el2_ifu_mem_ctl.scala 822:21]
  assign io_ifu_pmu_bus_error = _T_9312; // @[el2_ifu_mem_ctl.scala 823:24]
  assign io_ifu_pmu_bus_busy = _T_9316; // @[el2_ifu_mem_ctl.scala 824:23]
  assign io_ifu_pmu_bus_trxn = _T_9317; // @[el2_ifu_mem_ctl.scala 825:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 145:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 144:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 143:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 141:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 152:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 154:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 147:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 140:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 138:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 136:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 137:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 146:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 155:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 574:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_1729; // @[el2_ifu_mem_ctl.scala 575:19]
  assign io_ifu_axi_araddr = _T_1731 & _T_1733; // @[el2_ifu_mem_ctl.scala 576:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 579:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 151:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 577:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 580:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 142:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 578:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 153:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 581:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 671:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid; // @[el2_ifu_mem_ctl.scala 669:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata; // @[el2_ifu_mem_ctl.scala 673:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag; // @[el2_ifu_mem_ctl.scala 664:20]
  assign io_iccm_ready = _T_1832 & _T_1826; // @[el2_ifu_mem_ctl.scala 644:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 341:17]
  assign io_ic_wr_en = 2'h0; // @[el2_ifu_mem_ctl.scala 711:15]
  assign io_ic_rd_en = _T_3113 | _T_3118; // @[el2_ifu_mem_ctl.scala 702:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 356:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 356:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 357:23]
  assign io_ifu_ic_debug_rd_data = _T_366; // @[el2_ifu_mem_ctl.scala 365:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 828:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 830:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 831:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 829:25]
  assign io_ic_debug_way = _T_9329[1:0]; // @[el2_ifu_mem_ctl.scala 832:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_9303; // @[el2_ifu_mem_ctl.scala 816:19]
  assign io_iccm_rw_addr = _T_2267[14:0]; // @[el2_ifu_mem_ctl.scala 675:19]
  assign io_iccm_wren = _T_1836 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 646:16]
  assign io_iccm_rden = _T_1840 | _T_1841; // @[el2_ifu_mem_ctl.scala 647:16]
  assign io_iccm_wr_data = _T_2242 ? _T_2243 : _T_2250; // @[el2_ifu_mem_ctl.scala 652:19]
  assign io_iccm_wr_size = _T_1846 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 649:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 293:15]
  assign io_ic_access_fault_f = _T_1614 & _T_317; // @[el2_ifu_mem_ctl.scala 398:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_428; // @[el2_ifu_mem_ctl.scala 399:29]
  assign io_iccm_rd_ecc_single_err = _T_3058 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 688:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 689:29]
  assign io_ic_error_start = _T_354 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 359:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 194:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 193:24]
  assign io_ic_fetch_val_f = {1'h0,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 403:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 395:16]
  assign io_ic_premux_data = ic_premux_data[63:0]; // @[el2_ifu_mem_ctl.scala 392:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 393:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_9340; // @[el2_ifu_mem_ctl.scala 839:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_1619; // @[el2_ifu_mem_ctl.scala 493:27]
  assign io_iccm_correction_state = _T_1647 ? 1'h0 : _GEN_60; // @[el2_ifu_mem_ctl.scala 528:28 el2_ifu_mem_ctl.scala 541:32 el2_ifu_mem_ctl.scala 548:32 el2_ifu_mem_ctl.scala 555:32]
  assign io_data = {io_ic_wr_data_1,io_ic_wr_data_0}; // @[el2_ifu_mem_ctl.scala 354:11]
  assign io_ic_miss_buff_half = {_T_1530,_T_1610}; // @[el2_ifu_mem_ctl.scala 372:24]
  assign io_ic_wr_ecc = m1_io_ecc_out; // @[el2_ifu_mem_ctl.scala 350:16]
  assign m1_io_din = ifu_bus_rdata_ff; // @[el2_ifu_mem_ctl.scala 348:13]
  assign m2_io_din = {_T_1530,_T_1610}; // @[el2_ifu_mem_ctl.scala 352:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_4323 = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  _T_3679 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_3675 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  _T_3671 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  _T_3667 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  _T_3663 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  _T_3659 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  _T_3655 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  _T_3651 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  _T_3647 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  _T_3643 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  _T_3639 = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_3635 = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  _T_3631 = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  _T_3627 = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  _T_3623 = _RAND_36[2:0];
  _RAND_37 = {1{`RANDOM}};
  _T_3619 = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  _T_3615 = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  _T_3611 = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  _T_3607 = _RAND_40[2:0];
  _RAND_41 = {1{`RANDOM}};
  _T_3603 = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  _T_3599 = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  _T_3595 = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  _T_3591 = _RAND_44[2:0];
  _RAND_45 = {1{`RANDOM}};
  _T_3587 = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  _T_3583 = _RAND_46[2:0];
  _RAND_47 = {1{`RANDOM}};
  _T_3579 = _RAND_47[2:0];
  _RAND_48 = {1{`RANDOM}};
  _T_3575 = _RAND_48[2:0];
  _RAND_49 = {1{`RANDOM}};
  _T_3571 = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  _T_3567 = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  _T_3563 = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_3559 = _RAND_52[2:0];
  _RAND_53 = {1{`RANDOM}};
  _T_3555 = _RAND_53[2:0];
  _RAND_54 = {1{`RANDOM}};
  _T_3551 = _RAND_54[2:0];
  _RAND_55 = {1{`RANDOM}};
  _T_3547 = _RAND_55[2:0];
  _RAND_56 = {1{`RANDOM}};
  _T_3543 = _RAND_56[2:0];
  _RAND_57 = {1{`RANDOM}};
  _T_3539 = _RAND_57[2:0];
  _RAND_58 = {1{`RANDOM}};
  _T_3535 = _RAND_58[2:0];
  _RAND_59 = {1{`RANDOM}};
  _T_3531 = _RAND_59[2:0];
  _RAND_60 = {1{`RANDOM}};
  _T_3527 = _RAND_60[2:0];
  _RAND_61 = {1{`RANDOM}};
  _T_3523 = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  _T_3519 = _RAND_62[2:0];
  _RAND_63 = {1{`RANDOM}};
  _T_3515 = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  _T_3511 = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  _T_3507 = _RAND_65[2:0];
  _RAND_66 = {1{`RANDOM}};
  _T_3503 = _RAND_66[2:0];
  _RAND_67 = {1{`RANDOM}};
  _T_3499 = _RAND_67[2:0];
  _RAND_68 = {1{`RANDOM}};
  _T_3495 = _RAND_68[2:0];
  _RAND_69 = {1{`RANDOM}};
  _T_3491 = _RAND_69[2:0];
  _RAND_70 = {1{`RANDOM}};
  _T_3487 = _RAND_70[2:0];
  _RAND_71 = {1{`RANDOM}};
  _T_3483 = _RAND_71[2:0];
  _RAND_72 = {1{`RANDOM}};
  _T_3479 = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  _T_3475 = _RAND_73[2:0];
  _RAND_74 = {1{`RANDOM}};
  _T_3471 = _RAND_74[2:0];
  _RAND_75 = {1{`RANDOM}};
  _T_3467 = _RAND_75[2:0];
  _RAND_76 = {1{`RANDOM}};
  _T_3463 = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  _T_3459 = _RAND_77[2:0];
  _RAND_78 = {1{`RANDOM}};
  _T_3455 = _RAND_78[2:0];
  _RAND_79 = {1{`RANDOM}};
  _T_3451 = _RAND_79[2:0];
  _RAND_80 = {1{`RANDOM}};
  _T_3447 = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_3443 = _RAND_81[2:0];
  _RAND_82 = {1{`RANDOM}};
  _T_3439 = _RAND_82[2:0];
  _RAND_83 = {1{`RANDOM}};
  _T_3435 = _RAND_83[2:0];
  _RAND_84 = {1{`RANDOM}};
  _T_3431 = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  _T_3427 = _RAND_85[2:0];
  _RAND_86 = {1{`RANDOM}};
  _T_3423 = _RAND_86[2:0];
  _RAND_87 = {1{`RANDOM}};
  _T_3419 = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  _T_3415 = _RAND_88[2:0];
  _RAND_89 = {1{`RANDOM}};
  _T_3411 = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  _T_3407 = _RAND_90[2:0];
  _RAND_91 = {1{`RANDOM}};
  _T_3403 = _RAND_91[2:0];
  _RAND_92 = {1{`RANDOM}};
  _T_3399 = _RAND_92[2:0];
  _RAND_93 = {1{`RANDOM}};
  _T_3395 = _RAND_93[2:0];
  _RAND_94 = {1{`RANDOM}};
  _T_3391 = _RAND_94[2:0];
  _RAND_95 = {1{`RANDOM}};
  _T_3387 = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  _T_3383 = _RAND_96[2:0];
  _RAND_97 = {1{`RANDOM}};
  _T_3379 = _RAND_97[2:0];
  _RAND_98 = {1{`RANDOM}};
  _T_3375 = _RAND_98[2:0];
  _RAND_99 = {1{`RANDOM}};
  _T_3371 = _RAND_99[2:0];
  _RAND_100 = {1{`RANDOM}};
  _T_3367 = _RAND_100[2:0];
  _RAND_101 = {1{`RANDOM}};
  _T_3363 = _RAND_101[2:0];
  _RAND_102 = {1{`RANDOM}};
  _T_3359 = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  _T_3355 = _RAND_103[2:0];
  _RAND_104 = {1{`RANDOM}};
  _T_3351 = _RAND_104[2:0];
  _RAND_105 = {1{`RANDOM}};
  _T_3347 = _RAND_105[2:0];
  _RAND_106 = {1{`RANDOM}};
  _T_3343 = _RAND_106[2:0];
  _RAND_107 = {1{`RANDOM}};
  _T_3339 = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  _T_3335 = _RAND_108[2:0];
  _RAND_109 = {1{`RANDOM}};
  _T_3331 = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_3327 = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  _T_3323 = _RAND_111[2:0];
  _RAND_112 = {1{`RANDOM}};
  _T_3319 = _RAND_112[2:0];
  _RAND_113 = {1{`RANDOM}};
  _T_3315 = _RAND_113[2:0];
  _RAND_114 = {1{`RANDOM}};
  _T_3311 = _RAND_114[2:0];
  _RAND_115 = {1{`RANDOM}};
  _T_3307 = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  _T_3303 = _RAND_116[2:0];
  _RAND_117 = {1{`RANDOM}};
  _T_3299 = _RAND_117[2:0];
  _RAND_118 = {1{`RANDOM}};
  _T_3295 = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  _T_3291 = _RAND_119[2:0];
  _RAND_120 = {1{`RANDOM}};
  _T_3287 = _RAND_120[2:0];
  _RAND_121 = {1{`RANDOM}};
  _T_3283 = _RAND_121[2:0];
  _RAND_122 = {1{`RANDOM}};
  _T_3279 = _RAND_122[2:0];
  _RAND_123 = {1{`RANDOM}};
  _T_3275 = _RAND_123[2:0];
  _RAND_124 = {1{`RANDOM}};
  _T_3271 = _RAND_124[2:0];
  _RAND_125 = {1{`RANDOM}};
  _T_3267 = _RAND_125[2:0];
  _RAND_126 = {1{`RANDOM}};
  _T_3263 = _RAND_126[2:0];
  _RAND_127 = {1{`RANDOM}};
  _T_3259 = _RAND_127[2:0];
  _RAND_128 = {1{`RANDOM}};
  _T_3255 = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  _T_3251 = _RAND_129[2:0];
  _RAND_130 = {1{`RANDOM}};
  _T_3247 = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  _T_3243 = _RAND_131[2:0];
  _RAND_132 = {1{`RANDOM}};
  _T_3239 = _RAND_132[2:0];
  _RAND_133 = {1{`RANDOM}};
  _T_3235 = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  _T_3231 = _RAND_134[2:0];
  _RAND_135 = {1{`RANDOM}};
  _T_3227 = _RAND_135[2:0];
  _RAND_136 = {1{`RANDOM}};
  _T_3223 = _RAND_136[2:0];
  _RAND_137 = {1{`RANDOM}};
  _T_3219 = _RAND_137[2:0];
  _RAND_138 = {1{`RANDOM}};
  _T_3215 = _RAND_138[2:0];
  _RAND_139 = {1{`RANDOM}};
  _T_3211 = _RAND_139[2:0];
  _RAND_140 = {1{`RANDOM}};
  _T_3207 = _RAND_140[2:0];
  _RAND_141 = {1{`RANDOM}};
  _T_3203 = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  _T_3199 = _RAND_142[2:0];
  _RAND_143 = {1{`RANDOM}};
  _T_3195 = _RAND_143[2:0];
  _RAND_144 = {1{`RANDOM}};
  _T_3191 = _RAND_144[2:0];
  _RAND_145 = {1{`RANDOM}};
  _T_3187 = _RAND_145[2:0];
  _RAND_146 = {1{`RANDOM}};
  _T_3183 = _RAND_146[2:0];
  _RAND_147 = {1{`RANDOM}};
  _T_3179 = _RAND_147[2:0];
  _RAND_148 = {1{`RANDOM}};
  _T_3175 = _RAND_148[2:0];
  _RAND_149 = {1{`RANDOM}};
  _T_3171 = _RAND_149[2:0];
  _RAND_150 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_151[30:0];
  _RAND_152 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_152[2:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_156[1:0];
  _RAND_157 = {1{`RANDOM}};
  reset_ic_ff = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  miss_addr = _RAND_159[25:0];
  _RAND_160 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_161[2:0];
  _RAND_162 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_162[0:0];
  _RAND_163 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_163[63:0];
  _RAND_164 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_164[31:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_180[0:0];
  _RAND_181 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_439[1:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_440[0:0];
  _RAND_441 = {3{`RANDOM}};
  _T_366 = _RAND_441[70:0];
  _RAND_442 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_442[5:0];
  _RAND_443 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_443[0:0];
  _RAND_444 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_445[2:0];
  _RAND_446 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_446[0:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_448[0:0];
  _RAND_449 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_449[38:0];
  _RAND_450 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_450[1:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_451[2:0];
  _RAND_452 = {1{`RANDOM}};
  iccm_dma_rtag = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rvalid = _RAND_453[0:0];
  _RAND_454 = {2{`RANDOM}};
  iccm_dma_rdata = _RAND_454[63:0];
  _RAND_455 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_455[13:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_456[0:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_457[13:0];
  _RAND_458 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_458[6:0];
  _RAND_459 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_459[0:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_new_ff = _RAND_460[2:0];
  _RAND_461 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_461[1:0];
  _RAND_462 = {1{`RANDOM}};
  ic_valid_ff = _RAND_462[0:0];
  _RAND_463 = {1{`RANDOM}};
  _T_9310 = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_9311 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_9312 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_9316 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_9317 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_9340 = _RAND_468[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      _T_3679 <= 3'h0;
    end else if (_T_3678) begin
      _T_3679 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3675 <= 3'h0;
    end else if (_T_3674) begin
      _T_3675 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3671 <= 3'h0;
    end else if (_T_3670) begin
      _T_3671 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3667 <= 3'h0;
    end else if (_T_3666) begin
      _T_3667 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3663 <= 3'h0;
    end else if (_T_3662) begin
      _T_3663 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3659 <= 3'h0;
    end else if (_T_3658) begin
      _T_3659 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3655 <= 3'h0;
    end else if (_T_3654) begin
      _T_3655 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3651 <= 3'h0;
    end else if (_T_3650) begin
      _T_3651 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3647 <= 3'h0;
    end else if (_T_3646) begin
      _T_3647 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3643 <= 3'h0;
    end else if (_T_3642) begin
      _T_3643 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3639 <= 3'h0;
    end else if (_T_3638) begin
      _T_3639 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3635 <= 3'h0;
    end else if (_T_3634) begin
      _T_3635 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3631 <= 3'h0;
    end else if (_T_3630) begin
      _T_3631 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3627 <= 3'h0;
    end else if (_T_3626) begin
      _T_3627 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3623 <= 3'h0;
    end else if (_T_3622) begin
      _T_3623 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3619 <= 3'h0;
    end else if (_T_3618) begin
      _T_3619 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3615 <= 3'h0;
    end else if (_T_3614) begin
      _T_3615 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3611 <= 3'h0;
    end else if (_T_3610) begin
      _T_3611 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3607 <= 3'h0;
    end else if (_T_3606) begin
      _T_3607 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3603 <= 3'h0;
    end else if (_T_3602) begin
      _T_3603 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3599 <= 3'h0;
    end else if (_T_3598) begin
      _T_3599 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3595 <= 3'h0;
    end else if (_T_3594) begin
      _T_3595 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3591 <= 3'h0;
    end else if (_T_3590) begin
      _T_3591 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3587 <= 3'h0;
    end else if (_T_3586) begin
      _T_3587 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3583 <= 3'h0;
    end else if (_T_3582) begin
      _T_3583 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3579 <= 3'h0;
    end else if (_T_3578) begin
      _T_3579 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3575 <= 3'h0;
    end else if (_T_3574) begin
      _T_3575 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3571 <= 3'h0;
    end else if (_T_3570) begin
      _T_3571 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3567 <= 3'h0;
    end else if (_T_3566) begin
      _T_3567 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3563 <= 3'h0;
    end else if (_T_3562) begin
      _T_3563 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3559 <= 3'h0;
    end else if (_T_3558) begin
      _T_3559 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3555 <= 3'h0;
    end else if (_T_3554) begin
      _T_3555 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3551 <= 3'h0;
    end else if (_T_3550) begin
      _T_3551 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3547 <= 3'h0;
    end else if (_T_3546) begin
      _T_3547 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3543 <= 3'h0;
    end else if (_T_3542) begin
      _T_3543 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3539 <= 3'h0;
    end else if (_T_3538) begin
      _T_3539 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3535 <= 3'h0;
    end else if (_T_3534) begin
      _T_3535 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3531 <= 3'h0;
    end else if (_T_3530) begin
      _T_3531 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3527 <= 3'h0;
    end else if (_T_3526) begin
      _T_3527 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3523 <= 3'h0;
    end else if (_T_3522) begin
      _T_3523 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3519 <= 3'h0;
    end else if (_T_3518) begin
      _T_3519 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3515 <= 3'h0;
    end else if (_T_3514) begin
      _T_3515 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3511 <= 3'h0;
    end else if (_T_3510) begin
      _T_3511 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3507 <= 3'h0;
    end else if (_T_3506) begin
      _T_3507 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3503 <= 3'h0;
    end else if (_T_3502) begin
      _T_3503 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3499 <= 3'h0;
    end else if (_T_3498) begin
      _T_3499 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3495 <= 3'h0;
    end else if (_T_3494) begin
      _T_3495 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3491 <= 3'h0;
    end else if (_T_3490) begin
      _T_3491 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3487 <= 3'h0;
    end else if (_T_3486) begin
      _T_3487 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3483 <= 3'h0;
    end else if (_T_3482) begin
      _T_3483 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3479 <= 3'h0;
    end else if (_T_3478) begin
      _T_3479 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3475 <= 3'h0;
    end else if (_T_3474) begin
      _T_3475 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3471 <= 3'h0;
    end else if (_T_3470) begin
      _T_3471 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3467 <= 3'h0;
    end else if (_T_3466) begin
      _T_3467 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3463 <= 3'h0;
    end else if (_T_3462) begin
      _T_3463 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3459 <= 3'h0;
    end else if (_T_3458) begin
      _T_3459 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3455 <= 3'h0;
    end else if (_T_3454) begin
      _T_3455 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3451 <= 3'h0;
    end else if (_T_3450) begin
      _T_3451 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3447 <= 3'h0;
    end else if (_T_3446) begin
      _T_3447 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3443 <= 3'h0;
    end else if (_T_3442) begin
      _T_3443 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3439 <= 3'h0;
    end else if (_T_3438) begin
      _T_3439 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3435 <= 3'h0;
    end else if (_T_3434) begin
      _T_3435 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3431 <= 3'h0;
    end else if (_T_3430) begin
      _T_3431 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3427 <= 3'h0;
    end else if (_T_3426) begin
      _T_3427 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3423 <= 3'h0;
    end else if (_T_3422) begin
      _T_3423 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3419 <= 3'h0;
    end else if (_T_3418) begin
      _T_3419 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3415 <= 3'h0;
    end else if (_T_3414) begin
      _T_3415 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3411 <= 3'h0;
    end else if (_T_3410) begin
      _T_3411 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3407 <= 3'h0;
    end else if (_T_3406) begin
      _T_3407 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3403 <= 3'h0;
    end else if (_T_3402) begin
      _T_3403 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3399 <= 3'h0;
    end else if (_T_3398) begin
      _T_3399 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3395 <= 3'h0;
    end else if (_T_3394) begin
      _T_3395 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3391 <= 3'h0;
    end else if (_T_3390) begin
      _T_3391 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3387 <= 3'h0;
    end else if (_T_3386) begin
      _T_3387 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3383 <= 3'h0;
    end else if (_T_3382) begin
      _T_3383 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3379 <= 3'h0;
    end else if (_T_3378) begin
      _T_3379 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3375 <= 3'h0;
    end else if (_T_3374) begin
      _T_3375 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3371 <= 3'h0;
    end else if (_T_3370) begin
      _T_3371 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3367 <= 3'h0;
    end else if (_T_3366) begin
      _T_3367 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3363 <= 3'h0;
    end else if (_T_3362) begin
      _T_3363 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3359 <= 3'h0;
    end else if (_T_3358) begin
      _T_3359 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3355 <= 3'h0;
    end else if (_T_3354) begin
      _T_3355 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3351 <= 3'h0;
    end else if (_T_3350) begin
      _T_3351 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3347 <= 3'h0;
    end else if (_T_3346) begin
      _T_3347 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3343 <= 3'h0;
    end else if (_T_3342) begin
      _T_3343 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3339 <= 3'h0;
    end else if (_T_3338) begin
      _T_3339 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3335 <= 3'h0;
    end else if (_T_3334) begin
      _T_3335 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3331 <= 3'h0;
    end else if (_T_3330) begin
      _T_3331 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3327 <= 3'h0;
    end else if (_T_3326) begin
      _T_3327 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3323 <= 3'h0;
    end else if (_T_3322) begin
      _T_3323 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3319 <= 3'h0;
    end else if (_T_3318) begin
      _T_3319 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3315 <= 3'h0;
    end else if (_T_3314) begin
      _T_3315 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3311 <= 3'h0;
    end else if (_T_3310) begin
      _T_3311 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3307 <= 3'h0;
    end else if (_T_3306) begin
      _T_3307 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3303 <= 3'h0;
    end else if (_T_3302) begin
      _T_3303 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3299 <= 3'h0;
    end else if (_T_3298) begin
      _T_3299 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3295 <= 3'h0;
    end else if (_T_3294) begin
      _T_3295 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3291 <= 3'h0;
    end else if (_T_3290) begin
      _T_3291 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3287 <= 3'h0;
    end else if (_T_3286) begin
      _T_3287 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3283 <= 3'h0;
    end else if (_T_3282) begin
      _T_3283 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3279 <= 3'h0;
    end else if (_T_3278) begin
      _T_3279 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3275 <= 3'h0;
    end else if (_T_3274) begin
      _T_3275 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3271 <= 3'h0;
    end else if (_T_3270) begin
      _T_3271 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3267 <= 3'h0;
    end else if (_T_3266) begin
      _T_3267 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3263 <= 3'h0;
    end else if (_T_3262) begin
      _T_3263 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3259 <= 3'h0;
    end else if (_T_3258) begin
      _T_3259 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3255 <= 3'h0;
    end else if (_T_3254) begin
      _T_3255 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3251 <= 3'h0;
    end else if (_T_3250) begin
      _T_3251 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3247 <= 3'h0;
    end else if (_T_3246) begin
      _T_3247 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3243 <= 3'h0;
    end else if (_T_3242) begin
      _T_3243 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3239 <= 3'h0;
    end else if (_T_3238) begin
      _T_3239 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3235 <= 3'h0;
    end else if (_T_3234) begin
      _T_3235 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3231 <= 3'h0;
    end else if (_T_3230) begin
      _T_3231 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3227 <= 3'h0;
    end else if (_T_3226) begin
      _T_3227 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3223 <= 3'h0;
    end else if (_T_3222) begin
      _T_3223 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3219 <= 3'h0;
    end else if (_T_3218) begin
      _T_3219 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3215 <= 3'h0;
    end else if (_T_3214) begin
      _T_3215 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3211 <= 3'h0;
    end else if (_T_3210) begin
      _T_3211 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3207 <= 3'h0;
    end else if (_T_3206) begin
      _T_3207 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3203 <= 3'h0;
    end else if (_T_3202) begin
      _T_3203 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3199 <= 3'h0;
    end else if (_T_3198) begin
      _T_3199 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3195 <= 3'h0;
    end else if (_T_3194) begin
      _T_3195 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3191 <= 3'h0;
    end else if (_T_3190) begin
      _T_3191 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3187 <= 3'h0;
    end else if (_T_3186) begin
      _T_3187 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3183 <= 3'h0;
    end else if (_T_3182) begin
      _T_3183 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3179 <= 3'h0;
    end else if (_T_3178) begin
      _T_3179 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3175 <= 3'h0;
    end else if (_T_3174) begin
      _T_3175 <= way_status_new_ff;
    end
    if (reset) begin
      _T_3171 <= 3'h0;
    end else if (_T_3170) begin
      _T_3171 <= way_status_new_ff;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_289;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= 2'h0;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_1772) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_1768;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_4931) begin
      ic_tag_valid_out_1_0 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_4947) begin
      ic_tag_valid_out_1_1 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_4963) begin
      ic_tag_valid_out_1_2 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_4979) begin
      ic_tag_valid_out_1_3 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_4995) begin
      ic_tag_valid_out_1_4 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_5011) begin
      ic_tag_valid_out_1_5 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_5027) begin
      ic_tag_valid_out_1_6 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_5043) begin
      ic_tag_valid_out_1_7 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_5059) begin
      ic_tag_valid_out_1_8 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_5075) begin
      ic_tag_valid_out_1_9 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_5091) begin
      ic_tag_valid_out_1_10 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_5107) begin
      ic_tag_valid_out_1_11 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_5123) begin
      ic_tag_valid_out_1_12 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_5139) begin
      ic_tag_valid_out_1_13 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_5155) begin
      ic_tag_valid_out_1_14 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_5171) begin
      ic_tag_valid_out_1_15 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_5187) begin
      ic_tag_valid_out_1_16 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_5203) begin
      ic_tag_valid_out_1_17 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_5219) begin
      ic_tag_valid_out_1_18 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_5235) begin
      ic_tag_valid_out_1_19 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_5251) begin
      ic_tag_valid_out_1_20 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_5267) begin
      ic_tag_valid_out_1_21 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_5283) begin
      ic_tag_valid_out_1_22 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_5299) begin
      ic_tag_valid_out_1_23 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_5315) begin
      ic_tag_valid_out_1_24 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_5331) begin
      ic_tag_valid_out_1_25 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_5347) begin
      ic_tag_valid_out_1_26 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_5363) begin
      ic_tag_valid_out_1_27 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_5379) begin
      ic_tag_valid_out_1_28 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_5395) begin
      ic_tag_valid_out_1_29 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_5411) begin
      ic_tag_valid_out_1_30 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_5427) begin
      ic_tag_valid_out_1_31 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_5955) begin
      ic_tag_valid_out_1_32 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_5971) begin
      ic_tag_valid_out_1_33 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_5987) begin
      ic_tag_valid_out_1_34 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_6003) begin
      ic_tag_valid_out_1_35 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_6019) begin
      ic_tag_valid_out_1_36 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_6035) begin
      ic_tag_valid_out_1_37 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_6051) begin
      ic_tag_valid_out_1_38 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_6067) begin
      ic_tag_valid_out_1_39 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_6083) begin
      ic_tag_valid_out_1_40 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_6099) begin
      ic_tag_valid_out_1_41 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_6115) begin
      ic_tag_valid_out_1_42 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_6131) begin
      ic_tag_valid_out_1_43 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_6147) begin
      ic_tag_valid_out_1_44 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_6163) begin
      ic_tag_valid_out_1_45 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_6179) begin
      ic_tag_valid_out_1_46 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_6195) begin
      ic_tag_valid_out_1_47 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_6211) begin
      ic_tag_valid_out_1_48 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_6227) begin
      ic_tag_valid_out_1_49 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_6243) begin
      ic_tag_valid_out_1_50 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_6259) begin
      ic_tag_valid_out_1_51 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_6275) begin
      ic_tag_valid_out_1_52 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_6291) begin
      ic_tag_valid_out_1_53 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_6307) begin
      ic_tag_valid_out_1_54 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_6323) begin
      ic_tag_valid_out_1_55 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_6339) begin
      ic_tag_valid_out_1_56 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_6355) begin
      ic_tag_valid_out_1_57 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_6371) begin
      ic_tag_valid_out_1_58 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_6387) begin
      ic_tag_valid_out_1_59 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_6403) begin
      ic_tag_valid_out_1_60 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_6419) begin
      ic_tag_valid_out_1_61 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_6435) begin
      ic_tag_valid_out_1_62 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_6451) begin
      ic_tag_valid_out_1_63 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_6979) begin
      ic_tag_valid_out_1_64 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_6995) begin
      ic_tag_valid_out_1_65 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_7011) begin
      ic_tag_valid_out_1_66 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_7027) begin
      ic_tag_valid_out_1_67 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_7043) begin
      ic_tag_valid_out_1_68 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_7059) begin
      ic_tag_valid_out_1_69 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_7075) begin
      ic_tag_valid_out_1_70 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_7091) begin
      ic_tag_valid_out_1_71 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_7107) begin
      ic_tag_valid_out_1_72 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_7123) begin
      ic_tag_valid_out_1_73 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_7139) begin
      ic_tag_valid_out_1_74 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_7155) begin
      ic_tag_valid_out_1_75 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_7171) begin
      ic_tag_valid_out_1_76 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_7187) begin
      ic_tag_valid_out_1_77 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_7203) begin
      ic_tag_valid_out_1_78 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_7219) begin
      ic_tag_valid_out_1_79 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_7235) begin
      ic_tag_valid_out_1_80 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_7251) begin
      ic_tag_valid_out_1_81 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_7267) begin
      ic_tag_valid_out_1_82 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_7283) begin
      ic_tag_valid_out_1_83 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_7299) begin
      ic_tag_valid_out_1_84 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_7315) begin
      ic_tag_valid_out_1_85 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_7331) begin
      ic_tag_valid_out_1_86 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_7347) begin
      ic_tag_valid_out_1_87 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_7363) begin
      ic_tag_valid_out_1_88 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_7379) begin
      ic_tag_valid_out_1_89 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_7395) begin
      ic_tag_valid_out_1_90 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_7411) begin
      ic_tag_valid_out_1_91 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_7427) begin
      ic_tag_valid_out_1_92 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_7443) begin
      ic_tag_valid_out_1_93 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_7459) begin
      ic_tag_valid_out_1_94 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_7475) begin
      ic_tag_valid_out_1_95 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_8003) begin
      ic_tag_valid_out_1_96 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_8019) begin
      ic_tag_valid_out_1_97 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_8035) begin
      ic_tag_valid_out_1_98 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_8051) begin
      ic_tag_valid_out_1_99 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_8067) begin
      ic_tag_valid_out_1_100 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_8083) begin
      ic_tag_valid_out_1_101 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_8099) begin
      ic_tag_valid_out_1_102 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_8115) begin
      ic_tag_valid_out_1_103 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_8131) begin
      ic_tag_valid_out_1_104 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_8147) begin
      ic_tag_valid_out_1_105 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_8163) begin
      ic_tag_valid_out_1_106 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_8179) begin
      ic_tag_valid_out_1_107 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_8195) begin
      ic_tag_valid_out_1_108 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_8211) begin
      ic_tag_valid_out_1_109 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_8227) begin
      ic_tag_valid_out_1_110 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_8243) begin
      ic_tag_valid_out_1_111 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_8259) begin
      ic_tag_valid_out_1_112 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_8275) begin
      ic_tag_valid_out_1_113 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_8291) begin
      ic_tag_valid_out_1_114 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_8307) begin
      ic_tag_valid_out_1_115 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_8323) begin
      ic_tag_valid_out_1_116 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_8339) begin
      ic_tag_valid_out_1_117 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_8355) begin
      ic_tag_valid_out_1_118 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_8371) begin
      ic_tag_valid_out_1_119 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_8387) begin
      ic_tag_valid_out_1_120 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_8403) begin
      ic_tag_valid_out_1_121 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_8419) begin
      ic_tag_valid_out_1_122 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_8435) begin
      ic_tag_valid_out_1_123 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_8451) begin
      ic_tag_valid_out_1_124 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_8467) begin
      ic_tag_valid_out_1_125 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_8483) begin
      ic_tag_valid_out_1_126 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_8499) begin
      ic_tag_valid_out_1_127 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_4419) begin
      ic_tag_valid_out_0_0 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_4435) begin
      ic_tag_valid_out_0_1 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_4451) begin
      ic_tag_valid_out_0_2 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_4467) begin
      ic_tag_valid_out_0_3 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_4483) begin
      ic_tag_valid_out_0_4 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_4499) begin
      ic_tag_valid_out_0_5 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_4515) begin
      ic_tag_valid_out_0_6 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_4531) begin
      ic_tag_valid_out_0_7 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_4547) begin
      ic_tag_valid_out_0_8 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_4563) begin
      ic_tag_valid_out_0_9 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_4579) begin
      ic_tag_valid_out_0_10 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_4595) begin
      ic_tag_valid_out_0_11 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_4611) begin
      ic_tag_valid_out_0_12 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_4627) begin
      ic_tag_valid_out_0_13 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_4643) begin
      ic_tag_valid_out_0_14 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_4659) begin
      ic_tag_valid_out_0_15 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_4675) begin
      ic_tag_valid_out_0_16 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_4691) begin
      ic_tag_valid_out_0_17 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_4707) begin
      ic_tag_valid_out_0_18 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_4723) begin
      ic_tag_valid_out_0_19 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_4739) begin
      ic_tag_valid_out_0_20 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_4755) begin
      ic_tag_valid_out_0_21 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_4771) begin
      ic_tag_valid_out_0_22 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_4787) begin
      ic_tag_valid_out_0_23 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_4803) begin
      ic_tag_valid_out_0_24 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_4819) begin
      ic_tag_valid_out_0_25 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_4835) begin
      ic_tag_valid_out_0_26 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_4851) begin
      ic_tag_valid_out_0_27 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_4867) begin
      ic_tag_valid_out_0_28 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_4883) begin
      ic_tag_valid_out_0_29 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_4899) begin
      ic_tag_valid_out_0_30 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_4915) begin
      ic_tag_valid_out_0_31 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_5443) begin
      ic_tag_valid_out_0_32 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_5459) begin
      ic_tag_valid_out_0_33 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_5475) begin
      ic_tag_valid_out_0_34 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_5491) begin
      ic_tag_valid_out_0_35 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_5507) begin
      ic_tag_valid_out_0_36 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_5523) begin
      ic_tag_valid_out_0_37 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_5539) begin
      ic_tag_valid_out_0_38 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_5555) begin
      ic_tag_valid_out_0_39 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_5571) begin
      ic_tag_valid_out_0_40 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_5587) begin
      ic_tag_valid_out_0_41 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_5603) begin
      ic_tag_valid_out_0_42 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_5619) begin
      ic_tag_valid_out_0_43 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_5635) begin
      ic_tag_valid_out_0_44 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_5651) begin
      ic_tag_valid_out_0_45 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_5667) begin
      ic_tag_valid_out_0_46 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_5683) begin
      ic_tag_valid_out_0_47 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_5699) begin
      ic_tag_valid_out_0_48 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_5715) begin
      ic_tag_valid_out_0_49 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_5731) begin
      ic_tag_valid_out_0_50 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_5747) begin
      ic_tag_valid_out_0_51 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_5763) begin
      ic_tag_valid_out_0_52 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_5779) begin
      ic_tag_valid_out_0_53 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_5795) begin
      ic_tag_valid_out_0_54 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_5811) begin
      ic_tag_valid_out_0_55 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_5827) begin
      ic_tag_valid_out_0_56 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_5843) begin
      ic_tag_valid_out_0_57 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_5859) begin
      ic_tag_valid_out_0_58 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_5875) begin
      ic_tag_valid_out_0_59 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_5891) begin
      ic_tag_valid_out_0_60 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_5907) begin
      ic_tag_valid_out_0_61 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_5923) begin
      ic_tag_valid_out_0_62 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_5939) begin
      ic_tag_valid_out_0_63 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_6467) begin
      ic_tag_valid_out_0_64 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_6483) begin
      ic_tag_valid_out_0_65 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_6499) begin
      ic_tag_valid_out_0_66 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_6515) begin
      ic_tag_valid_out_0_67 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_6531) begin
      ic_tag_valid_out_0_68 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_6547) begin
      ic_tag_valid_out_0_69 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_6563) begin
      ic_tag_valid_out_0_70 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_6579) begin
      ic_tag_valid_out_0_71 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_6595) begin
      ic_tag_valid_out_0_72 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_6611) begin
      ic_tag_valid_out_0_73 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_6627) begin
      ic_tag_valid_out_0_74 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_6643) begin
      ic_tag_valid_out_0_75 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_6659) begin
      ic_tag_valid_out_0_76 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_6675) begin
      ic_tag_valid_out_0_77 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_6691) begin
      ic_tag_valid_out_0_78 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_6707) begin
      ic_tag_valid_out_0_79 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_6723) begin
      ic_tag_valid_out_0_80 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_6739) begin
      ic_tag_valid_out_0_81 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_6755) begin
      ic_tag_valid_out_0_82 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_6771) begin
      ic_tag_valid_out_0_83 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_6787) begin
      ic_tag_valid_out_0_84 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_6803) begin
      ic_tag_valid_out_0_85 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_6819) begin
      ic_tag_valid_out_0_86 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_6835) begin
      ic_tag_valid_out_0_87 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_6851) begin
      ic_tag_valid_out_0_88 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_6867) begin
      ic_tag_valid_out_0_89 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_6883) begin
      ic_tag_valid_out_0_90 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_6899) begin
      ic_tag_valid_out_0_91 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_6915) begin
      ic_tag_valid_out_0_92 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_6931) begin
      ic_tag_valid_out_0_93 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_6947) begin
      ic_tag_valid_out_0_94 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_6963) begin
      ic_tag_valid_out_0_95 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_7491) begin
      ic_tag_valid_out_0_96 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_7507) begin
      ic_tag_valid_out_0_97 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_7523) begin
      ic_tag_valid_out_0_98 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_7539) begin
      ic_tag_valid_out_0_99 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_7555) begin
      ic_tag_valid_out_0_100 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_7571) begin
      ic_tag_valid_out_0_101 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_7587) begin
      ic_tag_valid_out_0_102 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_7603) begin
      ic_tag_valid_out_0_103 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_7619) begin
      ic_tag_valid_out_0_104 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_7635) begin
      ic_tag_valid_out_0_105 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_7651) begin
      ic_tag_valid_out_0_106 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_7667) begin
      ic_tag_valid_out_0_107 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_7683) begin
      ic_tag_valid_out_0_108 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_7699) begin
      ic_tag_valid_out_0_109 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_7715) begin
      ic_tag_valid_out_0_110 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_7731) begin
      ic_tag_valid_out_0_111 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_7747) begin
      ic_tag_valid_out_0_112 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_7763) begin
      ic_tag_valid_out_0_113 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_7779) begin
      ic_tag_valid_out_0_114 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_7795) begin
      ic_tag_valid_out_0_115 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_7811) begin
      ic_tag_valid_out_0_116 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_7827) begin
      ic_tag_valid_out_0_117 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_7843) begin
      ic_tag_valid_out_0_118 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_7859) begin
      ic_tag_valid_out_0_119 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_7875) begin
      ic_tag_valid_out_0_120 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_7891) begin
      ic_tag_valid_out_0_121 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_7907) begin
      ic_tag_valid_out_0_122 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_7923) begin
      ic_tag_valid_out_0_123 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_7939) begin
      ic_tag_valid_out_0_124 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_7955) begin
      ic_tag_valid_out_0_125 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_7971) begin
      ic_tag_valid_out_0_126 <= _T_4410;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_7987) begin
      ic_tag_valid_out_0_127 <= _T_4410;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_366 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_366 <= {{5'd0}, _T_365};
      end else begin
        _T_366 <= io_ic_debug_rd_data;
      end
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_1721) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_1796) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_1840;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_1622) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_1624) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_1634) begin
        perr_state <= 3'h0;
      end else if (_T_1637) begin
        if (_T_1639) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_1643) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_1647) begin
        err_stop_state <= 2'h1;
      end else if (_T_1652) begin
        if (_T_1654) begin
          err_stop_state <= 2'h0;
        end else if (_T_1675) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_1679) begin
        if (_T_1654) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_1696) begin
        if (_T_1700) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_525;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      _T_4323 <= 7'h0;
    end else if (_T_3144) begin
      _T_4323 <= io_ic_debug_addr[9:3];
    end else begin
      _T_4323 <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_565;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_3079;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag <= 3'h0;
    end else begin
      iccm_dma_rtag <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid <= 1'h0;
    end else begin
      iccm_dma_rvalid <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata <= _T_2254;
    end else begin
      iccm_dma_rdata <= _T_2255;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_3075;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_3144) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 3'h0;
    end else if (_T_3147) begin
      way_status_new_ff <= _T_3151;
    end else begin
      way_status_new_ff <= {{2'd0}, way_status_new};
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_3147) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_9340 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_9340 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 6'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_9310 <= 1'h0;
    end else begin
      _T_9310 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_9311 <= 1'h0;
    end else begin
      _T_9311 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_9312 <= 1'h0;
    end else begin
      _T_9312 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_9316 <= 1'h0;
    end else begin
      _T_9316 <= _T_9315;
    end
    if (reset) begin
      _T_9317 <= 1'h0;
    end else begin
      _T_9317 <= bus_cmd_sent;
    end
  end
endmodule
