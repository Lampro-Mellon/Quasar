module el2_ifu_mem_ctl(
  input         clock,
  input         reset,
  input         io_free_clk,
  input         io_active_clk,
  input         io_exu_flush_final,
  input         io_dec_tlu_flush_lower_wb,
  input         io_dec_tlu_flush_err_wb,
  input         io_dec_tlu_i0_commit_cmt,
  input         io_dec_tlu_force_halt,
  input  [30:0] io_ifc_fetch_addr_bf,
  input         io_ifc_fetch_uncacheable_bf,
  input         io_ifc_fetch_req_bf,
  input         io_ifc_fetch_req_bf_raw,
  input         io_ifc_iccm_access_bf,
  input         io_ifc_region_acc_fault_bf,
  input         io_ifc_dma_access_ok,
  input         io_dec_tlu_fence_i_wb,
  input         io_ifu_bp_hit_taken_f,
  input         io_ifu_bp_inst_mask_f,
  input         io_ifu_axi_arready,
  input         io_ifu_axi_rvalid,
  input  [2:0]  io_ifu_axi_rid,
  input  [63:0] io_ifu_axi_rdata,
  input  [1:0]  io_ifu_axi_rresp,
  input         io_ifu_bus_clk_en,
  input         io_dma_iccm_req,
  input  [31:0] io_dma_mem_addr,
  input  [2:0]  io_dma_mem_sz,
  input         io_dma_mem_write,
  input  [63:0] io_dma_mem_wdata,
  input  [2:0]  io_dma_mem_tag,
  input  [63:0] io_ic_rd_data,
  input  [70:0] io_ic_debug_rd_data,
  input  [25:0] io_ictag_debug_rd_data,
  input  [1:0]  io_ic_eccerr,
  input  [1:0]  io_ic_parerr,
  input  [1:0]  io_ic_rd_hit,
  input         io_ic_tag_perr,
  input  [63:0] io_iccm_rd_data,
  input  [77:0] io_iccm_rd_data_ecc,
  input  [1:0]  io_ifu_fetch_val,
  input  [70:0] io_dec_tlu_ic_diag_pkt_icache_wrdata,
  input  [16:0] io_dec_tlu_ic_diag_pkt_icache_dicawics,
  input         io_dec_tlu_ic_diag_pkt_icache_rd_valid,
  input         io_dec_tlu_ic_diag_pkt_icache_wr_valid,
  output        io_ifu_miss_state_idle,
  output        io_ifu_ic_mb_empty,
  output        io_ic_dma_active,
  output        io_ic_write_stall,
  output        io_ifu_pmu_ic_miss,
  output        io_ifu_pmu_ic_hit,
  output        io_ifu_pmu_bus_error,
  output        io_ifu_pmu_bus_busy,
  output        io_ifu_pmu_bus_trxn,
  output        io_ifu_axi_awvalid,
  output [2:0]  io_ifu_axi_awid,
  output [31:0] io_ifu_axi_awaddr,
  output [3:0]  io_ifu_axi_awregion,
  output [7:0]  io_ifu_axi_awlen,
  output [2:0]  io_ifu_axi_awsize,
  output [1:0]  io_ifu_axi_awburst,
  output        io_ifu_axi_awlock,
  output [3:0]  io_ifu_axi_awcache,
  output [2:0]  io_ifu_axi_awprot,
  output [3:0]  io_ifu_axi_awqos,
  output        io_ifu_axi_wvalid,
  output [63:0] io_ifu_axi_wdata,
  output [7:0]  io_ifu_axi_wstrb,
  output        io_ifu_axi_wlast,
  output        io_ifu_axi_bready,
  output        io_ifu_axi_arvalid,
  output [2:0]  io_ifu_axi_arid,
  output [31:0] io_ifu_axi_araddr,
  output [3:0]  io_ifu_axi_arregion,
  output [7:0]  io_ifu_axi_arlen,
  output [2:0]  io_ifu_axi_arsize,
  output [1:0]  io_ifu_axi_arburst,
  output        io_ifu_axi_arlock,
  output [3:0]  io_ifu_axi_arcache,
  output [2:0]  io_ifu_axi_arprot,
  output [3:0]  io_ifu_axi_arqos,
  output        io_ifu_axi_rready,
  output        io_iccm_dma_ecc_error,
  output        io_iccm_dma_rvalid,
  output [63:0] io_iccm_dma_rdata,
  output [2:0]  io_iccm_dma_rtag,
  output        io_iccm_ready,
  output [30:0] io_ic_rw_addr,
  output [1:0]  io_ic_wr_en,
  output        io_ic_rd_en,
  output [70:0] io_ic_wr_data_0,
  output [70:0] io_ic_wr_data_1,
  output [70:0] io_ic_debug_wr_data,
  output [70:0] io_ifu_ic_debug_rd_data,
  output [9:0]  io_ic_debug_addr,
  output        io_ic_debug_rd_en,
  output        io_ic_debug_wr_en,
  output        io_ic_debug_tag_array,
  output [1:0]  io_ic_debug_way,
  output [1:0]  io_ic_tag_valid,
  output [14:0] io_iccm_rw_addr,
  output        io_iccm_wren,
  output        io_iccm_rden,
  output [77:0] io_iccm_wr_data,
  output [2:0]  io_iccm_wr_size,
  output        io_ic_hit_f,
  output        io_ic_access_fault_f,
  output [1:0]  io_ic_access_fault_type_f,
  output        io_iccm_rd_ecc_single_err,
  output        io_iccm_rd_ecc_double_err,
  output        io_ic_error_start,
  output        io_ifu_async_error_start,
  output        io_iccm_dma_sb_error,
  output [1:0]  io_ic_fetch_val_f,
  output [31:0] io_ic_data_f,
  output [63:0] io_ic_premux_data,
  output        io_ic_sel_premux_data,
  input         io_dec_tlu_core_ecc_disable,
  output        io_ifu_ic_debug_rd_data_valid,
  output        io_iccm_buf_correct_ecc,
  output        io_iccm_correction_state,
  input         io_scan_mode,
  output [6:0]  io_test
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [63:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_441;
  reg [95:0] _RAND_442;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_449;
  reg [63:0] _RAND_450;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_454;
  reg [63:0] _RAND_455;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_469;
`endif // RANDOMIZE_REG_INIT
  reg  flush_final_f; // @[el2_ifu_mem_ctl.scala 185:30]
  reg  ifc_fetch_req_f_raw; // @[el2_ifu_mem_ctl.scala 320:36]
  wire  _T_317 = ~io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 321:44]
  wire  ifc_fetch_req_f = ifc_fetch_req_f_raw & _T_317; // @[el2_ifu_mem_ctl.scala 321:42]
  reg [2:0] miss_state; // @[Reg.scala 27:20]
  wire  miss_pending = miss_state != 3'h0; // @[el2_ifu_mem_ctl.scala 253:30]
  reg  scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 547:52]
  wire  scnd_miss_req = scnd_miss_req_q & _T_317; // @[el2_ifu_mem_ctl.scala 549:36]
  wire  debug_c1_clken = io_ic_debug_rd_en | io_ic_debug_wr_en; // @[el2_ifu_mem_ctl.scala 187:42]
  wire [3:0] ic_fetch_val_int_f = {2'h0,io_ic_fetch_val_f}; // @[Cat.scala 29:58]
  reg [30:0] ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 308:34]
  wire [4:0] _GEN_464 = {{1'd0}, ic_fetch_val_int_f}; // @[el2_ifu_mem_ctl.scala 665:53]
  wire [4:0] ic_fetch_val_shift_right = _GEN_464 << ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 665:53]
  wire [1:0] _GEN_465 = {{1'd0}, _T_317}; // @[el2_ifu_mem_ctl.scala 668:91]
  wire [1:0] _T_3281 = ic_fetch_val_shift_right[3:2] & _GEN_465; // @[el2_ifu_mem_ctl.scala 668:91]
  reg  ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 322:31]
  wire  fetch_req_iccm_f = ifc_fetch_req_f & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 275:46]
  wire [1:0] _GEN_466 = {{1'd0}, fetch_req_iccm_f}; // @[el2_ifu_mem_ctl.scala 668:113]
  wire [1:0] _T_3282 = _T_3281 & _GEN_466; // @[el2_ifu_mem_ctl.scala 668:113]
  reg  iccm_dma_rvalid_in; // @[el2_ifu_mem_ctl.scala 654:59]
  wire [1:0] _GEN_467 = {{1'd0}, iccm_dma_rvalid_in}; // @[el2_ifu_mem_ctl.scala 668:130]
  wire [1:0] _T_3283 = _T_3282 | _GEN_467; // @[el2_ifu_mem_ctl.scala 668:130]
  wire  _T_3284 = ~io_dec_tlu_core_ecc_disable; // @[el2_ifu_mem_ctl.scala 668:154]
  wire [1:0] _GEN_468 = {{1'd0}, _T_3284}; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [1:0] _T_3285 = _T_3283 & _GEN_468; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [1:0] _T_3274 = ic_fetch_val_shift_right[1:0] & _GEN_465; // @[el2_ifu_mem_ctl.scala 668:91]
  wire [1:0] _T_3275 = _T_3274 & _GEN_466; // @[el2_ifu_mem_ctl.scala 668:113]
  wire [1:0] _T_3276 = _T_3275 | _GEN_467; // @[el2_ifu_mem_ctl.scala 668:130]
  wire [1:0] _T_3278 = _T_3276 & _GEN_468; // @[el2_ifu_mem_ctl.scala 668:152]
  wire [3:0] iccm_ecc_word_enable = {_T_3285,_T_3278}; // @[Cat.scala 29:58]
  wire  _T_3385 = ^io_iccm_rd_data_ecc[31:0]; // @[el2_lib.scala 318:30]
  wire  _T_3386 = ^io_iccm_rd_data_ecc[38:32]; // @[el2_lib.scala 318:44]
  wire  _T_3387 = _T_3385 ^ _T_3386; // @[el2_lib.scala 318:35]
  wire [5:0] _T_3395 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[26]}; // @[el2_lib.scala 318:76]
  wire  _T_3396 = ^_T_3395; // @[el2_lib.scala 318:83]
  wire  _T_3397 = io_iccm_rd_data_ecc[37] ^ _T_3396; // @[el2_lib.scala 318:71]
  wire [6:0] _T_3404 = {io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[11]}; // @[el2_lib.scala 318:103]
  wire [14:0] _T_3412 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3404}; // @[el2_lib.scala 318:103]
  wire  _T_3413 = ^_T_3412; // @[el2_lib.scala 318:110]
  wire  _T_3414 = io_iccm_rd_data_ecc[36] ^ _T_3413; // @[el2_lib.scala 318:98]
  wire [6:0] _T_3421 = {io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[4]}; // @[el2_lib.scala 318:130]
  wire [14:0] _T_3429 = {io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[18],_T_3421}; // @[el2_lib.scala 318:130]
  wire  _T_3430 = ^_T_3429; // @[el2_lib.scala 318:137]
  wire  _T_3431 = io_iccm_rd_data_ecc[35] ^ _T_3430; // @[el2_lib.scala 318:125]
  wire [8:0] _T_3440 = {io_iccm_rd_data_ecc[15],io_iccm_rd_data_ecc[14],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[7],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[1]}; // @[el2_lib.scala 318:157]
  wire [17:0] _T_3449 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[29],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[22],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3440}; // @[el2_lib.scala 318:157]
  wire  _T_3450 = ^_T_3449; // @[el2_lib.scala 318:164]
  wire  _T_3451 = io_iccm_rd_data_ecc[34] ^ _T_3450; // @[el2_lib.scala 318:152]
  wire [8:0] _T_3460 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[12],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[9],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[5],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[2],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 318:184]
  wire [17:0] _T_3469 = {io_iccm_rd_data_ecc[31],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[27],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[24],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[20],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[16],_T_3460}; // @[el2_lib.scala 318:184]
  wire  _T_3470 = ^_T_3469; // @[el2_lib.scala 318:191]
  wire  _T_3471 = io_iccm_rd_data_ecc[33] ^ _T_3470; // @[el2_lib.scala 318:179]
  wire [8:0] _T_3480 = {io_iccm_rd_data_ecc[13],io_iccm_rd_data_ecc[11],io_iccm_rd_data_ecc[10],io_iccm_rd_data_ecc[8],io_iccm_rd_data_ecc[6],io_iccm_rd_data_ecc[4],io_iccm_rd_data_ecc[3],io_iccm_rd_data_ecc[1],io_iccm_rd_data_ecc[0]}; // @[el2_lib.scala 318:211]
  wire [17:0] _T_3489 = {io_iccm_rd_data_ecc[30],io_iccm_rd_data_ecc[28],io_iccm_rd_data_ecc[26],io_iccm_rd_data_ecc[25],io_iccm_rd_data_ecc[23],io_iccm_rd_data_ecc[21],io_iccm_rd_data_ecc[19],io_iccm_rd_data_ecc[17],io_iccm_rd_data_ecc[15],_T_3480}; // @[el2_lib.scala 318:211]
  wire  _T_3490 = ^_T_3489; // @[el2_lib.scala 318:218]
  wire  _T_3491 = io_iccm_rd_data_ecc[32] ^ _T_3490; // @[el2_lib.scala 318:206]
  wire [6:0] _T_3497 = {_T_3387,_T_3397,_T_3414,_T_3431,_T_3451,_T_3471,_T_3491}; // @[Cat.scala 29:58]
  wire  _T_3498 = _T_3497 != 7'h0; // @[el2_lib.scala 319:44]
  wire  _T_3499 = iccm_ecc_word_enable[0] & _T_3498; // @[el2_lib.scala 319:32]
  wire  _T_3501 = _T_3499 & _T_3497[6]; // @[el2_lib.scala 319:53]
  wire  _T_3770 = ^io_iccm_rd_data_ecc[70:39]; // @[el2_lib.scala 318:30]
  wire  _T_3771 = ^io_iccm_rd_data_ecc[77:71]; // @[el2_lib.scala 318:44]
  wire  _T_3772 = _T_3770 ^ _T_3771; // @[el2_lib.scala 318:35]
  wire [5:0] _T_3780 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[65]}; // @[el2_lib.scala 318:76]
  wire  _T_3781 = ^_T_3780; // @[el2_lib.scala 318:83]
  wire  _T_3782 = io_iccm_rd_data_ecc[76] ^ _T_3781; // @[el2_lib.scala 318:71]
  wire [6:0] _T_3789 = {io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[50]}; // @[el2_lib.scala 318:103]
  wire [14:0] _T_3797 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3789}; // @[el2_lib.scala 318:103]
  wire  _T_3798 = ^_T_3797; // @[el2_lib.scala 318:110]
  wire  _T_3799 = io_iccm_rd_data_ecc[75] ^ _T_3798; // @[el2_lib.scala 318:98]
  wire [6:0] _T_3806 = {io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[43]}; // @[el2_lib.scala 318:130]
  wire [14:0] _T_3814 = {io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[57],_T_3806}; // @[el2_lib.scala 318:130]
  wire  _T_3815 = ^_T_3814; // @[el2_lib.scala 318:137]
  wire  _T_3816 = io_iccm_rd_data_ecc[74] ^ _T_3815; // @[el2_lib.scala 318:125]
  wire [8:0] _T_3825 = {io_iccm_rd_data_ecc[54],io_iccm_rd_data_ecc[53],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[46],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[40]}; // @[el2_lib.scala 318:157]
  wire [17:0] _T_3834 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[68],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[61],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3825}; // @[el2_lib.scala 318:157]
  wire  _T_3835 = ^_T_3834; // @[el2_lib.scala 318:164]
  wire  _T_3836 = io_iccm_rd_data_ecc[73] ^ _T_3835; // @[el2_lib.scala 318:152]
  wire [8:0] _T_3845 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[51],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[48],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[44],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[41],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 318:184]
  wire [17:0] _T_3854 = {io_iccm_rd_data_ecc[70],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[66],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[63],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[59],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[55],_T_3845}; // @[el2_lib.scala 318:184]
  wire  _T_3855 = ^_T_3854; // @[el2_lib.scala 318:191]
  wire  _T_3856 = io_iccm_rd_data_ecc[72] ^ _T_3855; // @[el2_lib.scala 318:179]
  wire [8:0] _T_3865 = {io_iccm_rd_data_ecc[52],io_iccm_rd_data_ecc[50],io_iccm_rd_data_ecc[49],io_iccm_rd_data_ecc[47],io_iccm_rd_data_ecc[45],io_iccm_rd_data_ecc[43],io_iccm_rd_data_ecc[42],io_iccm_rd_data_ecc[40],io_iccm_rd_data_ecc[39]}; // @[el2_lib.scala 318:211]
  wire [17:0] _T_3874 = {io_iccm_rd_data_ecc[69],io_iccm_rd_data_ecc[67],io_iccm_rd_data_ecc[65],io_iccm_rd_data_ecc[64],io_iccm_rd_data_ecc[62],io_iccm_rd_data_ecc[60],io_iccm_rd_data_ecc[58],io_iccm_rd_data_ecc[56],io_iccm_rd_data_ecc[54],_T_3865}; // @[el2_lib.scala 318:211]
  wire  _T_3875 = ^_T_3874; // @[el2_lib.scala 318:218]
  wire  _T_3876 = io_iccm_rd_data_ecc[71] ^ _T_3875; // @[el2_lib.scala 318:206]
  wire [6:0] _T_3882 = {_T_3772,_T_3782,_T_3799,_T_3816,_T_3836,_T_3856,_T_3876}; // @[Cat.scala 29:58]
  wire  _T_3883 = _T_3882 != 7'h0; // @[el2_lib.scala 319:44]
  wire  _T_3884 = iccm_ecc_word_enable[1] & _T_3883; // @[el2_lib.scala 319:32]
  wire  _T_3886 = _T_3884 & _T_3882[6]; // @[el2_lib.scala 319:53]
  wire [1:0] iccm_single_ecc_error = {_T_3501,_T_3886}; // @[Cat.scala 29:58]
  wire  _T_3 = |iccm_single_ecc_error; // @[el2_ifu_mem_ctl.scala 190:52]
  reg  dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 631:51]
  wire  _T_6 = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:57]
  reg [2:0] perr_state; // @[Reg.scala 27:20]
  wire  _T_7 = perr_state == 3'h4; // @[el2_ifu_mem_ctl.scala 192:54]
  wire  iccm_correct_ecc = perr_state == 3'h3; // @[el2_ifu_mem_ctl.scala 476:34]
  wire  _T_8 = iccm_correct_ecc | _T_7; // @[el2_ifu_mem_ctl.scala 192:40]
  reg [1:0] err_stop_state; // @[Reg.scala 27:20]
  wire  _T_9 = err_stop_state == 2'h3; // @[el2_ifu_mem_ctl.scala 192:90]
  wire  _T_10 = _T_8 | _T_9; // @[el2_ifu_mem_ctl.scala 192:72]
  wire  _T_2490 = 2'h0 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2495 = 2'h1 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2515 = io_ifu_fetch_val == 2'h3; // @[el2_ifu_mem_ctl.scala 526:48]
  wire  two_byte_instr = io_ic_data_f[1:0] != 2'h3; // @[el2_ifu_mem_ctl.scala 390:42]
  wire  _T_2517 = io_ifu_fetch_val[0] & two_byte_instr; // @[el2_ifu_mem_ctl.scala 526:79]
  wire  _T_2518 = _T_2515 | _T_2517; // @[el2_ifu_mem_ctl.scala 526:56]
  wire  _T_2519 = io_exu_flush_final | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 526:122]
  wire  _T_2520 = ~_T_2519; // @[el2_ifu_mem_ctl.scala 526:101]
  wire  _T_2521 = _T_2518 & _T_2520; // @[el2_ifu_mem_ctl.scala 526:99]
  wire  _T_2522 = 2'h2 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _T_2536 = io_ifu_fetch_val[0] & _T_317; // @[el2_ifu_mem_ctl.scala 533:45]
  wire  _T_2537 = ~io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 533:69]
  wire  _T_2538 = _T_2536 & _T_2537; // @[el2_ifu_mem_ctl.scala 533:67]
  wire  _T_2539 = 2'h3 == err_stop_state; // @[Conditional.scala 37:30]
  wire  _GEN_55 = _T_2522 ? _T_2538 : _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_59 = _T_2495 ? _T_2521 : _GEN_55; // @[Conditional.scala 39:67]
  wire  err_stop_fetch = _T_2490 ? 1'h0 : _GEN_59; // @[Conditional.scala 40:58]
  wire  _T_11 = _T_10 | err_stop_fetch; // @[el2_ifu_mem_ctl.scala 192:112]
  wire  _T_13 = io_ifu_axi_rvalid & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 194:44]
  wire  _T_14 = _T_13 & io_ifu_axi_rready; // @[el2_ifu_mem_ctl.scala 194:65]
  wire  _T_227 = |io_ic_rd_hit; // @[el2_ifu_mem_ctl.scala 283:37]
  wire  _T_228 = ~_T_227; // @[el2_ifu_mem_ctl.scala 283:23]
  reg  reset_all_tags; // @[el2_ifu_mem_ctl.scala 700:53]
  wire  _T_229 = _T_228 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 283:41]
  wire  _T_207 = ~ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 274:48]
  wire  _T_208 = ifc_fetch_req_f & _T_207; // @[el2_ifu_mem_ctl.scala 274:46]
  reg  ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 324:42]
  wire  _T_209 = ~ifc_region_acc_fault_final_f; // @[el2_ifu_mem_ctl.scala 274:69]
  wire  fetch_req_icache_f = _T_208 & _T_209; // @[el2_ifu_mem_ctl.scala 274:67]
  wire  _T_230 = _T_229 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 283:59]
  wire  _T_231 = ~miss_pending; // @[el2_ifu_mem_ctl.scala 283:82]
  wire  _T_232 = _T_230 & _T_231; // @[el2_ifu_mem_ctl.scala 283:80]
  wire  _T_233 = _T_232 | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 283:97]
  wire  ic_act_miss_f = _T_233 & _T_209; // @[el2_ifu_mem_ctl.scala 283:114]
  reg  ifu_bus_rvalid_unq_ff; // @[Reg.scala 27:20]
  reg  bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 546:61]
  wire  ifu_bus_rvalid_ff = ifu_bus_rvalid_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 588:49]
  wire  bus_ifu_wr_en_ff = ifu_bus_rvalid_ff & miss_pending; // @[el2_ifu_mem_ctl.scala 615:41]
  reg  uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 310:33]
  reg [2:0] bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 596:56]
  wire  _T_2641 = bus_data_beat_count == 3'h1; // @[el2_ifu_mem_ctl.scala 613:69]
  wire  _T_2642 = &bus_data_beat_count; // @[el2_ifu_mem_ctl.scala 613:101]
  wire  bus_last_data_beat = uncacheable_miss_ff ? _T_2641 : _T_2642; // @[el2_ifu_mem_ctl.scala 613:28]
  wire  _T_2588 = bus_ifu_wr_en_ff & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 592:68]
  wire  _T_2589 = ic_act_miss_f | _T_2588; // @[el2_ifu_mem_ctl.scala 592:48]
  wire  bus_reset_data_beat_cnt = _T_2589 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 592:91]
  wire  _T_2585 = ~bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 591:50]
  wire  _T_2586 = bus_ifu_wr_en_ff & _T_2585; // @[el2_ifu_mem_ctl.scala 591:48]
  wire  _T_2587 = ~io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 591:72]
  wire  bus_inc_data_beat_cnt = _T_2586 & _T_2587; // @[el2_ifu_mem_ctl.scala 591:70]
  wire [2:0] _T_2593 = bus_data_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 595:115]
  wire [2:0] _T_2595 = bus_inc_data_beat_cnt ? _T_2593 : 3'h0; // @[Mux.scala 27:72]
  wire  _T_2590 = ~bus_inc_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 593:32]
  wire  _T_2591 = ~bus_reset_data_beat_cnt; // @[el2_ifu_mem_ctl.scala 593:57]
  wire  bus_hold_data_beat_cnt = _T_2590 & _T_2591; // @[el2_ifu_mem_ctl.scala 593:55]
  wire [2:0] _T_2596 = bus_hold_data_beat_cnt ? bus_data_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] bus_new_data_beat_count = _T_2595 | _T_2596; // @[Mux.scala 27:72]
  wire  _T_15 = &bus_new_data_beat_count; // @[el2_ifu_mem_ctl.scala 194:112]
  wire  _T_16 = _T_14 & _T_15; // @[el2_ifu_mem_ctl.scala 194:85]
  wire  _T_17 = ~uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 195:5]
  wire  _T_18 = _T_16 & _T_17; // @[el2_ifu_mem_ctl.scala 194:118]
  wire  _T_19 = miss_state == 3'h5; // @[el2_ifu_mem_ctl.scala 195:41]
  wire  _T_24 = 3'h0 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_26 = ic_act_miss_f & _T_317; // @[el2_ifu_mem_ctl.scala 201:43]
  wire [2:0] _T_28 = _T_26 ? 3'h1 : 3'h2; // @[el2_ifu_mem_ctl.scala 201:27]
  wire  _T_31 = 3'h1 == miss_state; // @[Conditional.scala 37:30]
  wire [4:0] byp_fetch_index = ifu_fetch_addr_int_f[4:0]; // @[el2_ifu_mem_ctl.scala 426:45]
  wire  _T_2120 = byp_fetch_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 447:127]
  reg [7:0] ic_miss_buff_data_valid; // @[el2_ifu_mem_ctl.scala 403:60]
  wire  _T_2151 = _T_2120 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2124 = byp_fetch_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2152 = _T_2124 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2159 = _T_2151 | _T_2152; // @[Mux.scala 27:72]
  wire  _T_2128 = byp_fetch_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2153 = _T_2128 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2160 = _T_2159 | _T_2153; // @[Mux.scala 27:72]
  wire  _T_2132 = byp_fetch_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2154 = _T_2132 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2161 = _T_2160 | _T_2154; // @[Mux.scala 27:72]
  wire  _T_2136 = byp_fetch_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2155 = _T_2136 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2162 = _T_2161 | _T_2155; // @[Mux.scala 27:72]
  wire  _T_2140 = byp_fetch_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2156 = _T_2140 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2163 = _T_2162 | _T_2156; // @[Mux.scala 27:72]
  wire  _T_2144 = byp_fetch_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2157 = _T_2144 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2164 = _T_2163 | _T_2157; // @[Mux.scala 27:72]
  wire  _T_2148 = byp_fetch_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 447:127]
  wire  _T_2158 = _T_2148 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_bypass_index = _T_2164 | _T_2158; // @[Mux.scala 27:72]
  wire  _T_2206 = ~byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 449:69]
  wire  _T_2207 = ic_miss_buff_data_valid_bypass_index & _T_2206; // @[el2_ifu_mem_ctl.scala 449:67]
  wire  _T_2209 = ~byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 449:91]
  wire  _T_2210 = _T_2207 & _T_2209; // @[el2_ifu_mem_ctl.scala 449:89]
  wire  _T_2215 = _T_2207 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 450:65]
  wire  _T_2216 = _T_2210 | _T_2215; // @[el2_ifu_mem_ctl.scala 449:112]
  wire  _T_2218 = ic_miss_buff_data_valid_bypass_index & byp_fetch_index[1]; // @[el2_ifu_mem_ctl.scala 451:43]
  wire  _T_2221 = _T_2218 & _T_2209; // @[el2_ifu_mem_ctl.scala 451:65]
  wire  _T_2222 = _T_2216 | _T_2221; // @[el2_ifu_mem_ctl.scala 450:88]
  wire  _T_2226 = _T_2218 & byp_fetch_index[0]; // @[el2_ifu_mem_ctl.scala 452:65]
  wire [2:0] byp_fetch_index_inc = ifu_fetch_addr_int_f[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 429:75]
  wire  _T_2166 = byp_fetch_index_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2190 = _T_2166 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2169 = byp_fetch_index_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2191 = _T_2169 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2198 = _T_2190 | _T_2191; // @[Mux.scala 27:72]
  wire  _T_2172 = byp_fetch_index_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2192 = _T_2172 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2199 = _T_2198 | _T_2192; // @[Mux.scala 27:72]
  wire  _T_2175 = byp_fetch_index_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2193 = _T_2175 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2200 = _T_2199 | _T_2193; // @[Mux.scala 27:72]
  wire  _T_2178 = byp_fetch_index_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2194 = _T_2178 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2201 = _T_2200 | _T_2194; // @[Mux.scala 27:72]
  wire  _T_2181 = byp_fetch_index_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2195 = _T_2181 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2202 = _T_2201 | _T_2195; // @[Mux.scala 27:72]
  wire  _T_2184 = byp_fetch_index_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2196 = _T_2184 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2203 = _T_2202 | _T_2196; // @[Mux.scala 27:72]
  wire  _T_2187 = byp_fetch_index_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 448:110]
  wire  _T_2197 = _T_2187 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_valid_inc_bypass_index = _T_2203 | _T_2197; // @[Mux.scala 27:72]
  wire  _T_2227 = _T_2226 & ic_miss_buff_data_valid_inc_bypass_index; // @[el2_ifu_mem_ctl.scala 452:87]
  wire  _T_2228 = _T_2222 | _T_2227; // @[el2_ifu_mem_ctl.scala 451:88]
  wire  _T_2232 = ic_miss_buff_data_valid_bypass_index & _T_2148; // @[el2_ifu_mem_ctl.scala 453:43]
  wire  miss_buff_hit_unq_f = _T_2228 | _T_2232; // @[el2_ifu_mem_ctl.scala 452:131]
  wire  _T_2248 = miss_state == 3'h4; // @[el2_ifu_mem_ctl.scala 458:55]
  wire  _T_2249 = miss_state == 3'h1; // @[el2_ifu_mem_ctl.scala 458:87]
  wire  _T_2250 = _T_2248 | _T_2249; // @[el2_ifu_mem_ctl.scala 458:74]
  wire  crit_byp_hit_f = miss_buff_hit_unq_f & _T_2250; // @[el2_ifu_mem_ctl.scala 458:41]
  wire  _T_2233 = miss_state == 3'h6; // @[el2_ifu_mem_ctl.scala 455:30]
  reg [30:0] imb_ff; // @[el2_ifu_mem_ctl.scala 311:20]
  wire  miss_wrap_f = imb_ff[5] != ifu_fetch_addr_int_f[5]; // @[el2_ifu_mem_ctl.scala 446:51]
  wire  _T_2234 = ~miss_wrap_f; // @[el2_ifu_mem_ctl.scala 455:68]
  wire  _T_2235 = miss_buff_hit_unq_f & _T_2234; // @[el2_ifu_mem_ctl.scala 455:66]
  wire  stream_hit_f = _T_2233 & _T_2235; // @[el2_ifu_mem_ctl.scala 455:43]
  wire  _T_215 = crit_byp_hit_f | stream_hit_f; // @[el2_ifu_mem_ctl.scala 278:35]
  wire  _T_216 = _T_215 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 278:52]
  wire  ic_byp_hit_f = _T_216 & miss_pending; // @[el2_ifu_mem_ctl.scala 278:73]
  reg  last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 598:58]
  wire  last_beat = bus_last_data_beat & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 625:35]
  wire  _T_32 = bus_ifu_wr_en_ff & last_beat; // @[el2_ifu_mem_ctl.scala 205:113]
  wire  _T_33 = last_data_recieved_ff | _T_32; // @[el2_ifu_mem_ctl.scala 205:93]
  wire  _T_34 = ic_byp_hit_f & _T_33; // @[el2_ifu_mem_ctl.scala 205:67]
  wire  _T_35 = _T_34 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 205:127]
  wire  _T_36 = io_dec_tlu_force_halt | _T_35; // @[el2_ifu_mem_ctl.scala 205:51]
  wire  _T_38 = ~last_data_recieved_ff; // @[el2_ifu_mem_ctl.scala 206:30]
  wire  _T_39 = ic_byp_hit_f & _T_38; // @[el2_ifu_mem_ctl.scala 206:27]
  wire  _T_40 = _T_39 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 206:53]
  wire  _T_42 = ~ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 207:16]
  wire  _T_44 = _T_42 & _T_317; // @[el2_ifu_mem_ctl.scala 207:30]
  wire  _T_46 = _T_44 & _T_32; // @[el2_ifu_mem_ctl.scala 207:52]
  wire  _T_47 = _T_46 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 207:85]
  wire  _T_51 = _T_32 & _T_17; // @[el2_ifu_mem_ctl.scala 208:49]
  wire  _T_54 = ic_byp_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 209:33]
  wire  _T_56 = ~_T_32; // @[el2_ifu_mem_ctl.scala 209:57]
  wire  _T_57 = _T_54 & _T_56; // @[el2_ifu_mem_ctl.scala 209:55]
  wire  ifu_bp_hit_taken_q_f = io_ifu_bp_hit_taken_f & io_ic_hit_f; // @[el2_ifu_mem_ctl.scala 197:52]
  wire  _T_58 = ~ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 209:91]
  wire  _T_59 = _T_57 & _T_58; // @[el2_ifu_mem_ctl.scala 209:89]
  wire  _T_61 = _T_59 & _T_17; // @[el2_ifu_mem_ctl.scala 209:113]
  wire  _T_64 = bus_ifu_wr_en_ff & _T_317; // @[el2_ifu_mem_ctl.scala 210:39]
  wire  _T_67 = _T_64 & _T_56; // @[el2_ifu_mem_ctl.scala 210:61]
  wire  _T_69 = _T_67 & _T_58; // @[el2_ifu_mem_ctl.scala 210:95]
  wire  _T_71 = _T_69 & _T_17; // @[el2_ifu_mem_ctl.scala 210:119]
  wire  _T_79 = _T_46 & _T_17; // @[el2_ifu_mem_ctl.scala 211:100]
  wire  _T_81 = io_exu_flush_final | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 212:44]
  wire  _T_84 = _T_81 & _T_56; // @[el2_ifu_mem_ctl.scala 212:68]
  wire [2:0] _T_86 = _T_84 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 212:22]
  wire [2:0] _T_87 = _T_79 ? 3'h0 : _T_86; // @[el2_ifu_mem_ctl.scala 211:20]
  wire [2:0] _T_88 = _T_71 ? 3'h6 : _T_87; // @[el2_ifu_mem_ctl.scala 210:20]
  wire [2:0] _T_89 = _T_61 ? 3'h6 : _T_88; // @[el2_ifu_mem_ctl.scala 209:18]
  wire [2:0] _T_90 = _T_51 ? 3'h0 : _T_89; // @[el2_ifu_mem_ctl.scala 208:16]
  wire [2:0] _T_91 = _T_47 ? 3'h4 : _T_90; // @[el2_ifu_mem_ctl.scala 207:14]
  wire [2:0] _T_92 = _T_40 ? 3'h3 : _T_91; // @[el2_ifu_mem_ctl.scala 206:12]
  wire [2:0] _T_93 = _T_36 ? 3'h0 : _T_92; // @[el2_ifu_mem_ctl.scala 205:27]
  wire  _T_102 = 3'h4 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_106 = 3'h6 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_2245 = byp_fetch_index[4:1] == 4'hf; // @[el2_ifu_mem_ctl.scala 457:60]
  wire  _T_2246 = _T_2245 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 457:94]
  wire  stream_eol_f = _T_2246 & stream_hit_f; // @[el2_ifu_mem_ctl.scala 457:112]
  wire  _T_108 = _T_81 | stream_eol_f; // @[el2_ifu_mem_ctl.scala 220:72]
  wire  _T_111 = _T_108 & _T_56; // @[el2_ifu_mem_ctl.scala 220:87]
  wire  _T_113 = _T_111 & _T_2587; // @[el2_ifu_mem_ctl.scala 220:122]
  wire [2:0] _T_115 = _T_113 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 220:27]
  wire  _T_121 = 3'h3 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_124 = io_exu_flush_final & _T_56; // @[el2_ifu_mem_ctl.scala 224:48]
  wire  _T_126 = _T_124 & _T_2587; // @[el2_ifu_mem_ctl.scala 224:82]
  wire [2:0] _T_128 = _T_126 ? 3'h2 : 3'h0; // @[el2_ifu_mem_ctl.scala 224:27]
  wire  _T_132 = 3'h2 == miss_state; // @[Conditional.scala 37:30]
  wire  _T_236 = io_ic_rd_hit == 2'h0; // @[el2_ifu_mem_ctl.scala 284:28]
  wire  _T_237 = _T_236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 284:42]
  wire  _T_238 = _T_237 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 284:60]
  wire  _T_239 = miss_state == 3'h2; // @[el2_ifu_mem_ctl.scala 284:94]
  wire  _T_240 = _T_238 & _T_239; // @[el2_ifu_mem_ctl.scala 284:81]
  wire  _T_243 = imb_ff[30:5] != ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 285:39]
  wire  _T_244 = _T_240 & _T_243; // @[el2_ifu_mem_ctl.scala 284:111]
  wire  _T_246 = _T_244 & _T_17; // @[el2_ifu_mem_ctl.scala 285:91]
  reg  sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 338:51]
  wire  _T_247 = ~sel_mb_addr_ff; // @[el2_ifu_mem_ctl.scala 285:116]
  wire  _T_248 = _T_246 & _T_247; // @[el2_ifu_mem_ctl.scala 285:114]
  wire  ic_miss_under_miss_f = _T_248 & _T_209; // @[el2_ifu_mem_ctl.scala 285:132]
  wire  _T_135 = ic_miss_under_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 228:50]
  wire  _T_137 = _T_135 & _T_2587; // @[el2_ifu_mem_ctl.scala 228:84]
  wire  _T_256 = _T_230 & _T_239; // @[el2_ifu_mem_ctl.scala 286:85]
  wire  _T_259 = imb_ff[30:5] == ifu_fetch_addr_int_f[30:5]; // @[el2_ifu_mem_ctl.scala 287:39]
  wire  _T_260 = _T_259 | uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 287:91]
  wire  ic_ignore_2nd_miss_f = _T_256 & _T_260; // @[el2_ifu_mem_ctl.scala 286:117]
  wire  _T_141 = ic_ignore_2nd_miss_f & _T_56; // @[el2_ifu_mem_ctl.scala 229:35]
  wire  _T_143 = _T_141 & _T_2587; // @[el2_ifu_mem_ctl.scala 229:69]
  wire [2:0] _T_145 = _T_143 ? 3'h7 : 3'h0; // @[el2_ifu_mem_ctl.scala 229:12]
  wire [2:0] _T_146 = _T_137 ? 3'h5 : _T_145; // @[el2_ifu_mem_ctl.scala 228:27]
  wire  _T_151 = 3'h5 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_154 = _T_32 ? 3'h0 : 3'h2; // @[el2_ifu_mem_ctl.scala 234:12]
  wire [2:0] _T_155 = io_exu_flush_final ? _T_154 : 3'h1; // @[el2_ifu_mem_ctl.scala 233:62]
  wire [2:0] _T_156 = io_dec_tlu_force_halt ? 3'h0 : _T_155; // @[el2_ifu_mem_ctl.scala 233:27]
  wire  _T_160 = 3'h7 == miss_state; // @[Conditional.scala 37:30]
  wire [2:0] _T_164 = io_exu_flush_final ? _T_154 : 3'h0; // @[el2_ifu_mem_ctl.scala 238:62]
  wire [2:0] _T_165 = io_dec_tlu_force_halt ? 3'h0 : _T_164; // @[el2_ifu_mem_ctl.scala 238:27]
  wire [2:0] _GEN_0 = _T_160 ? _T_165 : 3'h0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_2 = _T_151 ? _T_156 : _GEN_0; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_4 = _T_132 ? _T_146 : _GEN_2; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_6 = _T_121 ? _T_128 : _GEN_4; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_8 = _T_106 ? _T_115 : _GEN_6; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_10 = _T_102 ? 3'h0 : _GEN_8; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_12 = _T_31 ? _T_93 : _GEN_10; // @[Conditional.scala 39:67]
  wire [2:0] miss_nxtstate = _T_24 ? _T_28 : _GEN_12; // @[Conditional.scala 40:58]
  wire  _T_20 = miss_nxtstate == 3'h5; // @[el2_ifu_mem_ctl.scala 195:73]
  wire  _T_21 = _T_19 | _T_20; // @[el2_ifu_mem_ctl.scala 195:57]
  wire  _T_22 = _T_18 & _T_21; // @[el2_ifu_mem_ctl.scala 195:26]
  wire  scnd_miss_req_in = _T_22 & _T_317; // @[el2_ifu_mem_ctl.scala 195:91]
  wire  _T_30 = ic_act_miss_f & _T_2587; // @[el2_ifu_mem_ctl.scala 202:38]
  wire  _T_94 = io_dec_tlu_force_halt | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 213:46]
  wire  _T_95 = _T_94 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 213:67]
  wire  _T_96 = _T_95 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 213:82]
  wire  _T_98 = _T_96 | _T_32; // @[el2_ifu_mem_ctl.scala 213:105]
  wire  _T_100 = bus_ifu_wr_en_ff & _T_17; // @[el2_ifu_mem_ctl.scala 213:158]
  wire  _T_101 = _T_98 | _T_100; // @[el2_ifu_mem_ctl.scala 213:138]
  wire  _T_103 = io_exu_flush_final | flush_final_f; // @[el2_ifu_mem_ctl.scala 217:43]
  wire  _T_104 = _T_103 | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 217:59]
  wire  _T_105 = _T_104 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 217:74]
  wire  _T_119 = _T_108 | _T_32; // @[el2_ifu_mem_ctl.scala 221:84]
  wire  _T_120 = _T_119 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 221:118]
  wire  _T_130 = io_exu_flush_final | _T_32; // @[el2_ifu_mem_ctl.scala 225:43]
  wire  _T_131 = _T_130 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 225:76]
  wire  _T_148 = _T_32 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 230:55]
  wire  _T_149 = _T_148 | ic_ignore_2nd_miss_f; // @[el2_ifu_mem_ctl.scala 230:78]
  wire  _T_150 = _T_149 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 230:101]
  wire  _T_158 = _T_32 | io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 235:55]
  wire  _T_159 = _T_158 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 235:76]
  wire  _GEN_1 = _T_160 & _T_159; // @[Conditional.scala 39:67]
  wire  _GEN_3 = _T_151 ? _T_159 : _GEN_1; // @[Conditional.scala 39:67]
  wire  _GEN_5 = _T_132 ? _T_150 : _GEN_3; // @[Conditional.scala 39:67]
  wire  _GEN_7 = _T_121 ? _T_131 : _GEN_5; // @[Conditional.scala 39:67]
  wire  _GEN_9 = _T_106 ? _T_120 : _GEN_7; // @[Conditional.scala 39:67]
  wire  _GEN_11 = _T_102 ? _T_105 : _GEN_9; // @[Conditional.scala 39:67]
  wire  _GEN_13 = _T_31 ? _T_101 : _GEN_11; // @[Conditional.scala 39:67]
  wire  miss_state_en = _T_24 ? _T_30 : _GEN_13; // @[Conditional.scala 40:58]
  wire  _T_174 = ~flush_final_f; // @[el2_ifu_mem_ctl.scala 254:95]
  wire  _T_175 = _T_2248 & _T_174; // @[el2_ifu_mem_ctl.scala 254:93]
  wire  crit_wd_byp_ok_ff = _T_2249 | _T_175; // @[el2_ifu_mem_ctl.scala 254:58]
  wire  _T_178 = miss_pending & _T_56; // @[el2_ifu_mem_ctl.scala 255:36]
  wire  _T_180 = _T_2248 & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 255:106]
  wire  _T_181 = ~_T_180; // @[el2_ifu_mem_ctl.scala 255:72]
  wire  _T_182 = _T_178 & _T_181; // @[el2_ifu_mem_ctl.scala 255:70]
  wire  _T_184 = _T_2248 & crit_byp_hit_f; // @[el2_ifu_mem_ctl.scala 256:57]
  wire  _T_185 = ~_T_184; // @[el2_ifu_mem_ctl.scala 256:23]
  wire  _T_186 = _T_182 & _T_185; // @[el2_ifu_mem_ctl.scala 255:128]
  wire  _T_187 = _T_186 | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 256:77]
  wire  _T_188 = miss_nxtstate == 3'h4; // @[el2_ifu_mem_ctl.scala 257:36]
  wire  _T_189 = miss_pending & _T_188; // @[el2_ifu_mem_ctl.scala 257:19]
  wire  sel_hold_imb = _T_187 | _T_189; // @[el2_ifu_mem_ctl.scala 256:93]
  wire  _T_191 = _T_19 | ic_miss_under_miss_f; // @[el2_ifu_mem_ctl.scala 259:57]
  wire  sel_hold_imb_scnd = _T_191 & _T_174; // @[el2_ifu_mem_ctl.scala 259:81]
  reg  way_status_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 267:35]
  reg [6:0] ifu_ic_rw_int_addr_ff; // @[el2_ifu_mem_ctl.scala 734:14]
  wire  _T_4949 = ifu_ic_rw_int_addr_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_0; // @[Reg.scala 27:20]
  wire  _T_5077 = _T_4949 & way_status_out_0; // @[Mux.scala 27:72]
  wire  _T_4950 = ifu_ic_rw_int_addr_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_1; // @[Reg.scala 27:20]
  wire  _T_5078 = _T_4950 & way_status_out_1; // @[Mux.scala 27:72]
  wire  _T_5205 = _T_5077 | _T_5078; // @[Mux.scala 27:72]
  wire  _T_4951 = ifu_ic_rw_int_addr_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_2; // @[Reg.scala 27:20]
  wire  _T_5079 = _T_4951 & way_status_out_2; // @[Mux.scala 27:72]
  wire  _T_5206 = _T_5205 | _T_5079; // @[Mux.scala 27:72]
  wire  _T_4952 = ifu_ic_rw_int_addr_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_3; // @[Reg.scala 27:20]
  wire  _T_5080 = _T_4952 & way_status_out_3; // @[Mux.scala 27:72]
  wire  _T_5207 = _T_5206 | _T_5080; // @[Mux.scala 27:72]
  wire  _T_4953 = ifu_ic_rw_int_addr_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_4; // @[Reg.scala 27:20]
  wire  _T_5081 = _T_4953 & way_status_out_4; // @[Mux.scala 27:72]
  wire  _T_5208 = _T_5207 | _T_5081; // @[Mux.scala 27:72]
  wire  _T_4954 = ifu_ic_rw_int_addr_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_5; // @[Reg.scala 27:20]
  wire  _T_5082 = _T_4954 & way_status_out_5; // @[Mux.scala 27:72]
  wire  _T_5209 = _T_5208 | _T_5082; // @[Mux.scala 27:72]
  wire  _T_4955 = ifu_ic_rw_int_addr_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_6; // @[Reg.scala 27:20]
  wire  _T_5083 = _T_4955 & way_status_out_6; // @[Mux.scala 27:72]
  wire  _T_5210 = _T_5209 | _T_5083; // @[Mux.scala 27:72]
  wire  _T_4956 = ifu_ic_rw_int_addr_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_7; // @[Reg.scala 27:20]
  wire  _T_5084 = _T_4956 & way_status_out_7; // @[Mux.scala 27:72]
  wire  _T_5211 = _T_5210 | _T_5084; // @[Mux.scala 27:72]
  wire  _T_4957 = ifu_ic_rw_int_addr_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_8; // @[Reg.scala 27:20]
  wire  _T_5085 = _T_4957 & way_status_out_8; // @[Mux.scala 27:72]
  wire  _T_5212 = _T_5211 | _T_5085; // @[Mux.scala 27:72]
  wire  _T_4958 = ifu_ic_rw_int_addr_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_9; // @[Reg.scala 27:20]
  wire  _T_5086 = _T_4958 & way_status_out_9; // @[Mux.scala 27:72]
  wire  _T_5213 = _T_5212 | _T_5086; // @[Mux.scala 27:72]
  wire  _T_4959 = ifu_ic_rw_int_addr_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_10; // @[Reg.scala 27:20]
  wire  _T_5087 = _T_4959 & way_status_out_10; // @[Mux.scala 27:72]
  wire  _T_5214 = _T_5213 | _T_5087; // @[Mux.scala 27:72]
  wire  _T_4960 = ifu_ic_rw_int_addr_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_11; // @[Reg.scala 27:20]
  wire  _T_5088 = _T_4960 & way_status_out_11; // @[Mux.scala 27:72]
  wire  _T_5215 = _T_5214 | _T_5088; // @[Mux.scala 27:72]
  wire  _T_4961 = ifu_ic_rw_int_addr_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_12; // @[Reg.scala 27:20]
  wire  _T_5089 = _T_4961 & way_status_out_12; // @[Mux.scala 27:72]
  wire  _T_5216 = _T_5215 | _T_5089; // @[Mux.scala 27:72]
  wire  _T_4962 = ifu_ic_rw_int_addr_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_13; // @[Reg.scala 27:20]
  wire  _T_5090 = _T_4962 & way_status_out_13; // @[Mux.scala 27:72]
  wire  _T_5217 = _T_5216 | _T_5090; // @[Mux.scala 27:72]
  wire  _T_4963 = ifu_ic_rw_int_addr_ff == 7'he; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_14; // @[Reg.scala 27:20]
  wire  _T_5091 = _T_4963 & way_status_out_14; // @[Mux.scala 27:72]
  wire  _T_5218 = _T_5217 | _T_5091; // @[Mux.scala 27:72]
  wire  _T_4964 = ifu_ic_rw_int_addr_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_15; // @[Reg.scala 27:20]
  wire  _T_5092 = _T_4964 & way_status_out_15; // @[Mux.scala 27:72]
  wire  _T_5219 = _T_5218 | _T_5092; // @[Mux.scala 27:72]
  wire  _T_4965 = ifu_ic_rw_int_addr_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_16; // @[Reg.scala 27:20]
  wire  _T_5093 = _T_4965 & way_status_out_16; // @[Mux.scala 27:72]
  wire  _T_5220 = _T_5219 | _T_5093; // @[Mux.scala 27:72]
  wire  _T_4966 = ifu_ic_rw_int_addr_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_17; // @[Reg.scala 27:20]
  wire  _T_5094 = _T_4966 & way_status_out_17; // @[Mux.scala 27:72]
  wire  _T_5221 = _T_5220 | _T_5094; // @[Mux.scala 27:72]
  wire  _T_4967 = ifu_ic_rw_int_addr_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_18; // @[Reg.scala 27:20]
  wire  _T_5095 = _T_4967 & way_status_out_18; // @[Mux.scala 27:72]
  wire  _T_5222 = _T_5221 | _T_5095; // @[Mux.scala 27:72]
  wire  _T_4968 = ifu_ic_rw_int_addr_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_19; // @[Reg.scala 27:20]
  wire  _T_5096 = _T_4968 & way_status_out_19; // @[Mux.scala 27:72]
  wire  _T_5223 = _T_5222 | _T_5096; // @[Mux.scala 27:72]
  wire  _T_4969 = ifu_ic_rw_int_addr_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_20; // @[Reg.scala 27:20]
  wire  _T_5097 = _T_4969 & way_status_out_20; // @[Mux.scala 27:72]
  wire  _T_5224 = _T_5223 | _T_5097; // @[Mux.scala 27:72]
  wire  _T_4970 = ifu_ic_rw_int_addr_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_21; // @[Reg.scala 27:20]
  wire  _T_5098 = _T_4970 & way_status_out_21; // @[Mux.scala 27:72]
  wire  _T_5225 = _T_5224 | _T_5098; // @[Mux.scala 27:72]
  wire  _T_4971 = ifu_ic_rw_int_addr_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_22; // @[Reg.scala 27:20]
  wire  _T_5099 = _T_4971 & way_status_out_22; // @[Mux.scala 27:72]
  wire  _T_5226 = _T_5225 | _T_5099; // @[Mux.scala 27:72]
  wire  _T_4972 = ifu_ic_rw_int_addr_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_23; // @[Reg.scala 27:20]
  wire  _T_5100 = _T_4972 & way_status_out_23; // @[Mux.scala 27:72]
  wire  _T_5227 = _T_5226 | _T_5100; // @[Mux.scala 27:72]
  wire  _T_4973 = ifu_ic_rw_int_addr_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_24; // @[Reg.scala 27:20]
  wire  _T_5101 = _T_4973 & way_status_out_24; // @[Mux.scala 27:72]
  wire  _T_5228 = _T_5227 | _T_5101; // @[Mux.scala 27:72]
  wire  _T_4974 = ifu_ic_rw_int_addr_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_25; // @[Reg.scala 27:20]
  wire  _T_5102 = _T_4974 & way_status_out_25; // @[Mux.scala 27:72]
  wire  _T_5229 = _T_5228 | _T_5102; // @[Mux.scala 27:72]
  wire  _T_4975 = ifu_ic_rw_int_addr_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_26; // @[Reg.scala 27:20]
  wire  _T_5103 = _T_4975 & way_status_out_26; // @[Mux.scala 27:72]
  wire  _T_5230 = _T_5229 | _T_5103; // @[Mux.scala 27:72]
  wire  _T_4976 = ifu_ic_rw_int_addr_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_27; // @[Reg.scala 27:20]
  wire  _T_5104 = _T_4976 & way_status_out_27; // @[Mux.scala 27:72]
  wire  _T_5231 = _T_5230 | _T_5104; // @[Mux.scala 27:72]
  wire  _T_4977 = ifu_ic_rw_int_addr_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_28; // @[Reg.scala 27:20]
  wire  _T_5105 = _T_4977 & way_status_out_28; // @[Mux.scala 27:72]
  wire  _T_5232 = _T_5231 | _T_5105; // @[Mux.scala 27:72]
  wire  _T_4978 = ifu_ic_rw_int_addr_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_29; // @[Reg.scala 27:20]
  wire  _T_5106 = _T_4978 & way_status_out_29; // @[Mux.scala 27:72]
  wire  _T_5233 = _T_5232 | _T_5106; // @[Mux.scala 27:72]
  wire  _T_4979 = ifu_ic_rw_int_addr_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_30; // @[Reg.scala 27:20]
  wire  _T_5107 = _T_4979 & way_status_out_30; // @[Mux.scala 27:72]
  wire  _T_5234 = _T_5233 | _T_5107; // @[Mux.scala 27:72]
  wire  _T_4980 = ifu_ic_rw_int_addr_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_31; // @[Reg.scala 27:20]
  wire  _T_5108 = _T_4980 & way_status_out_31; // @[Mux.scala 27:72]
  wire  _T_5235 = _T_5234 | _T_5108; // @[Mux.scala 27:72]
  wire  _T_4981 = ifu_ic_rw_int_addr_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_32; // @[Reg.scala 27:20]
  wire  _T_5109 = _T_4981 & way_status_out_32; // @[Mux.scala 27:72]
  wire  _T_5236 = _T_5235 | _T_5109; // @[Mux.scala 27:72]
  wire  _T_4982 = ifu_ic_rw_int_addr_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_33; // @[Reg.scala 27:20]
  wire  _T_5110 = _T_4982 & way_status_out_33; // @[Mux.scala 27:72]
  wire  _T_5237 = _T_5236 | _T_5110; // @[Mux.scala 27:72]
  wire  _T_4983 = ifu_ic_rw_int_addr_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_34; // @[Reg.scala 27:20]
  wire  _T_5111 = _T_4983 & way_status_out_34; // @[Mux.scala 27:72]
  wire  _T_5238 = _T_5237 | _T_5111; // @[Mux.scala 27:72]
  wire  _T_4984 = ifu_ic_rw_int_addr_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_35; // @[Reg.scala 27:20]
  wire  _T_5112 = _T_4984 & way_status_out_35; // @[Mux.scala 27:72]
  wire  _T_5239 = _T_5238 | _T_5112; // @[Mux.scala 27:72]
  wire  _T_4985 = ifu_ic_rw_int_addr_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_36; // @[Reg.scala 27:20]
  wire  _T_5113 = _T_4985 & way_status_out_36; // @[Mux.scala 27:72]
  wire  _T_5240 = _T_5239 | _T_5113; // @[Mux.scala 27:72]
  wire  _T_4986 = ifu_ic_rw_int_addr_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_37; // @[Reg.scala 27:20]
  wire  _T_5114 = _T_4986 & way_status_out_37; // @[Mux.scala 27:72]
  wire  _T_5241 = _T_5240 | _T_5114; // @[Mux.scala 27:72]
  wire  _T_4987 = ifu_ic_rw_int_addr_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_38; // @[Reg.scala 27:20]
  wire  _T_5115 = _T_4987 & way_status_out_38; // @[Mux.scala 27:72]
  wire  _T_5242 = _T_5241 | _T_5115; // @[Mux.scala 27:72]
  wire  _T_4988 = ifu_ic_rw_int_addr_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_39; // @[Reg.scala 27:20]
  wire  _T_5116 = _T_4988 & way_status_out_39; // @[Mux.scala 27:72]
  wire  _T_5243 = _T_5242 | _T_5116; // @[Mux.scala 27:72]
  wire  _T_4989 = ifu_ic_rw_int_addr_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_40; // @[Reg.scala 27:20]
  wire  _T_5117 = _T_4989 & way_status_out_40; // @[Mux.scala 27:72]
  wire  _T_5244 = _T_5243 | _T_5117; // @[Mux.scala 27:72]
  wire  _T_4990 = ifu_ic_rw_int_addr_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_41; // @[Reg.scala 27:20]
  wire  _T_5118 = _T_4990 & way_status_out_41; // @[Mux.scala 27:72]
  wire  _T_5245 = _T_5244 | _T_5118; // @[Mux.scala 27:72]
  wire  _T_4991 = ifu_ic_rw_int_addr_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_42; // @[Reg.scala 27:20]
  wire  _T_5119 = _T_4991 & way_status_out_42; // @[Mux.scala 27:72]
  wire  _T_5246 = _T_5245 | _T_5119; // @[Mux.scala 27:72]
  wire  _T_4992 = ifu_ic_rw_int_addr_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_43; // @[Reg.scala 27:20]
  wire  _T_5120 = _T_4992 & way_status_out_43; // @[Mux.scala 27:72]
  wire  _T_5247 = _T_5246 | _T_5120; // @[Mux.scala 27:72]
  wire  _T_4993 = ifu_ic_rw_int_addr_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_44; // @[Reg.scala 27:20]
  wire  _T_5121 = _T_4993 & way_status_out_44; // @[Mux.scala 27:72]
  wire  _T_5248 = _T_5247 | _T_5121; // @[Mux.scala 27:72]
  wire  _T_4994 = ifu_ic_rw_int_addr_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_45; // @[Reg.scala 27:20]
  wire  _T_5122 = _T_4994 & way_status_out_45; // @[Mux.scala 27:72]
  wire  _T_5249 = _T_5248 | _T_5122; // @[Mux.scala 27:72]
  wire  _T_4995 = ifu_ic_rw_int_addr_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_46; // @[Reg.scala 27:20]
  wire  _T_5123 = _T_4995 & way_status_out_46; // @[Mux.scala 27:72]
  wire  _T_5250 = _T_5249 | _T_5123; // @[Mux.scala 27:72]
  wire  _T_4996 = ifu_ic_rw_int_addr_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_47; // @[Reg.scala 27:20]
  wire  _T_5124 = _T_4996 & way_status_out_47; // @[Mux.scala 27:72]
  wire  _T_5251 = _T_5250 | _T_5124; // @[Mux.scala 27:72]
  wire  _T_4997 = ifu_ic_rw_int_addr_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_48; // @[Reg.scala 27:20]
  wire  _T_5125 = _T_4997 & way_status_out_48; // @[Mux.scala 27:72]
  wire  _T_5252 = _T_5251 | _T_5125; // @[Mux.scala 27:72]
  wire  _T_4998 = ifu_ic_rw_int_addr_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_49; // @[Reg.scala 27:20]
  wire  _T_5126 = _T_4998 & way_status_out_49; // @[Mux.scala 27:72]
  wire  _T_5253 = _T_5252 | _T_5126; // @[Mux.scala 27:72]
  wire  _T_4999 = ifu_ic_rw_int_addr_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_50; // @[Reg.scala 27:20]
  wire  _T_5127 = _T_4999 & way_status_out_50; // @[Mux.scala 27:72]
  wire  _T_5254 = _T_5253 | _T_5127; // @[Mux.scala 27:72]
  wire  _T_5000 = ifu_ic_rw_int_addr_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_51; // @[Reg.scala 27:20]
  wire  _T_5128 = _T_5000 & way_status_out_51; // @[Mux.scala 27:72]
  wire  _T_5255 = _T_5254 | _T_5128; // @[Mux.scala 27:72]
  wire  _T_5001 = ifu_ic_rw_int_addr_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_52; // @[Reg.scala 27:20]
  wire  _T_5129 = _T_5001 & way_status_out_52; // @[Mux.scala 27:72]
  wire  _T_5256 = _T_5255 | _T_5129; // @[Mux.scala 27:72]
  wire  _T_5002 = ifu_ic_rw_int_addr_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_53; // @[Reg.scala 27:20]
  wire  _T_5130 = _T_5002 & way_status_out_53; // @[Mux.scala 27:72]
  wire  _T_5257 = _T_5256 | _T_5130; // @[Mux.scala 27:72]
  wire  _T_5003 = ifu_ic_rw_int_addr_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_54; // @[Reg.scala 27:20]
  wire  _T_5131 = _T_5003 & way_status_out_54; // @[Mux.scala 27:72]
  wire  _T_5258 = _T_5257 | _T_5131; // @[Mux.scala 27:72]
  wire  _T_5004 = ifu_ic_rw_int_addr_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_55; // @[Reg.scala 27:20]
  wire  _T_5132 = _T_5004 & way_status_out_55; // @[Mux.scala 27:72]
  wire  _T_5259 = _T_5258 | _T_5132; // @[Mux.scala 27:72]
  wire  _T_5005 = ifu_ic_rw_int_addr_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_56; // @[Reg.scala 27:20]
  wire  _T_5133 = _T_5005 & way_status_out_56; // @[Mux.scala 27:72]
  wire  _T_5260 = _T_5259 | _T_5133; // @[Mux.scala 27:72]
  wire  _T_5006 = ifu_ic_rw_int_addr_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_57; // @[Reg.scala 27:20]
  wire  _T_5134 = _T_5006 & way_status_out_57; // @[Mux.scala 27:72]
  wire  _T_5261 = _T_5260 | _T_5134; // @[Mux.scala 27:72]
  wire  _T_5007 = ifu_ic_rw_int_addr_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_58; // @[Reg.scala 27:20]
  wire  _T_5135 = _T_5007 & way_status_out_58; // @[Mux.scala 27:72]
  wire  _T_5262 = _T_5261 | _T_5135; // @[Mux.scala 27:72]
  wire  _T_5008 = ifu_ic_rw_int_addr_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_59; // @[Reg.scala 27:20]
  wire  _T_5136 = _T_5008 & way_status_out_59; // @[Mux.scala 27:72]
  wire  _T_5263 = _T_5262 | _T_5136; // @[Mux.scala 27:72]
  wire  _T_5009 = ifu_ic_rw_int_addr_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_60; // @[Reg.scala 27:20]
  wire  _T_5137 = _T_5009 & way_status_out_60; // @[Mux.scala 27:72]
  wire  _T_5264 = _T_5263 | _T_5137; // @[Mux.scala 27:72]
  wire  _T_5010 = ifu_ic_rw_int_addr_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_61; // @[Reg.scala 27:20]
  wire  _T_5138 = _T_5010 & way_status_out_61; // @[Mux.scala 27:72]
  wire  _T_5265 = _T_5264 | _T_5138; // @[Mux.scala 27:72]
  wire  _T_5011 = ifu_ic_rw_int_addr_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_62; // @[Reg.scala 27:20]
  wire  _T_5139 = _T_5011 & way_status_out_62; // @[Mux.scala 27:72]
  wire  _T_5266 = _T_5265 | _T_5139; // @[Mux.scala 27:72]
  wire  _T_5012 = ifu_ic_rw_int_addr_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_63; // @[Reg.scala 27:20]
  wire  _T_5140 = _T_5012 & way_status_out_63; // @[Mux.scala 27:72]
  wire  _T_5267 = _T_5266 | _T_5140; // @[Mux.scala 27:72]
  wire  _T_5013 = ifu_ic_rw_int_addr_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_64; // @[Reg.scala 27:20]
  wire  _T_5141 = _T_5013 & way_status_out_64; // @[Mux.scala 27:72]
  wire  _T_5268 = _T_5267 | _T_5141; // @[Mux.scala 27:72]
  wire  _T_5014 = ifu_ic_rw_int_addr_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_65; // @[Reg.scala 27:20]
  wire  _T_5142 = _T_5014 & way_status_out_65; // @[Mux.scala 27:72]
  wire  _T_5269 = _T_5268 | _T_5142; // @[Mux.scala 27:72]
  wire  _T_5015 = ifu_ic_rw_int_addr_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_66; // @[Reg.scala 27:20]
  wire  _T_5143 = _T_5015 & way_status_out_66; // @[Mux.scala 27:72]
  wire  _T_5270 = _T_5269 | _T_5143; // @[Mux.scala 27:72]
  wire  _T_5016 = ifu_ic_rw_int_addr_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_67; // @[Reg.scala 27:20]
  wire  _T_5144 = _T_5016 & way_status_out_67; // @[Mux.scala 27:72]
  wire  _T_5271 = _T_5270 | _T_5144; // @[Mux.scala 27:72]
  wire  _T_5017 = ifu_ic_rw_int_addr_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_68; // @[Reg.scala 27:20]
  wire  _T_5145 = _T_5017 & way_status_out_68; // @[Mux.scala 27:72]
  wire  _T_5272 = _T_5271 | _T_5145; // @[Mux.scala 27:72]
  wire  _T_5018 = ifu_ic_rw_int_addr_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_69; // @[Reg.scala 27:20]
  wire  _T_5146 = _T_5018 & way_status_out_69; // @[Mux.scala 27:72]
  wire  _T_5273 = _T_5272 | _T_5146; // @[Mux.scala 27:72]
  wire  _T_5019 = ifu_ic_rw_int_addr_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_70; // @[Reg.scala 27:20]
  wire  _T_5147 = _T_5019 & way_status_out_70; // @[Mux.scala 27:72]
  wire  _T_5274 = _T_5273 | _T_5147; // @[Mux.scala 27:72]
  wire  _T_5020 = ifu_ic_rw_int_addr_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_71; // @[Reg.scala 27:20]
  wire  _T_5148 = _T_5020 & way_status_out_71; // @[Mux.scala 27:72]
  wire  _T_5275 = _T_5274 | _T_5148; // @[Mux.scala 27:72]
  wire  _T_5021 = ifu_ic_rw_int_addr_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_72; // @[Reg.scala 27:20]
  wire  _T_5149 = _T_5021 & way_status_out_72; // @[Mux.scala 27:72]
  wire  _T_5276 = _T_5275 | _T_5149; // @[Mux.scala 27:72]
  wire  _T_5022 = ifu_ic_rw_int_addr_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_73; // @[Reg.scala 27:20]
  wire  _T_5150 = _T_5022 & way_status_out_73; // @[Mux.scala 27:72]
  wire  _T_5277 = _T_5276 | _T_5150; // @[Mux.scala 27:72]
  wire  _T_5023 = ifu_ic_rw_int_addr_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_74; // @[Reg.scala 27:20]
  wire  _T_5151 = _T_5023 & way_status_out_74; // @[Mux.scala 27:72]
  wire  _T_5278 = _T_5277 | _T_5151; // @[Mux.scala 27:72]
  wire  _T_5024 = ifu_ic_rw_int_addr_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_75; // @[Reg.scala 27:20]
  wire  _T_5152 = _T_5024 & way_status_out_75; // @[Mux.scala 27:72]
  wire  _T_5279 = _T_5278 | _T_5152; // @[Mux.scala 27:72]
  wire  _T_5025 = ifu_ic_rw_int_addr_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_76; // @[Reg.scala 27:20]
  wire  _T_5153 = _T_5025 & way_status_out_76; // @[Mux.scala 27:72]
  wire  _T_5280 = _T_5279 | _T_5153; // @[Mux.scala 27:72]
  wire  _T_5026 = ifu_ic_rw_int_addr_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_77; // @[Reg.scala 27:20]
  wire  _T_5154 = _T_5026 & way_status_out_77; // @[Mux.scala 27:72]
  wire  _T_5281 = _T_5280 | _T_5154; // @[Mux.scala 27:72]
  wire  _T_5027 = ifu_ic_rw_int_addr_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_78; // @[Reg.scala 27:20]
  wire  _T_5155 = _T_5027 & way_status_out_78; // @[Mux.scala 27:72]
  wire  _T_5282 = _T_5281 | _T_5155; // @[Mux.scala 27:72]
  wire  _T_5028 = ifu_ic_rw_int_addr_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_79; // @[Reg.scala 27:20]
  wire  _T_5156 = _T_5028 & way_status_out_79; // @[Mux.scala 27:72]
  wire  _T_5283 = _T_5282 | _T_5156; // @[Mux.scala 27:72]
  wire  _T_5029 = ifu_ic_rw_int_addr_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_80; // @[Reg.scala 27:20]
  wire  _T_5157 = _T_5029 & way_status_out_80; // @[Mux.scala 27:72]
  wire  _T_5284 = _T_5283 | _T_5157; // @[Mux.scala 27:72]
  wire  _T_5030 = ifu_ic_rw_int_addr_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_81; // @[Reg.scala 27:20]
  wire  _T_5158 = _T_5030 & way_status_out_81; // @[Mux.scala 27:72]
  wire  _T_5285 = _T_5284 | _T_5158; // @[Mux.scala 27:72]
  wire  _T_5031 = ifu_ic_rw_int_addr_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_82; // @[Reg.scala 27:20]
  wire  _T_5159 = _T_5031 & way_status_out_82; // @[Mux.scala 27:72]
  wire  _T_5286 = _T_5285 | _T_5159; // @[Mux.scala 27:72]
  wire  _T_5032 = ifu_ic_rw_int_addr_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_83; // @[Reg.scala 27:20]
  wire  _T_5160 = _T_5032 & way_status_out_83; // @[Mux.scala 27:72]
  wire  _T_5287 = _T_5286 | _T_5160; // @[Mux.scala 27:72]
  wire  _T_5033 = ifu_ic_rw_int_addr_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_84; // @[Reg.scala 27:20]
  wire  _T_5161 = _T_5033 & way_status_out_84; // @[Mux.scala 27:72]
  wire  _T_5288 = _T_5287 | _T_5161; // @[Mux.scala 27:72]
  wire  _T_5034 = ifu_ic_rw_int_addr_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_85; // @[Reg.scala 27:20]
  wire  _T_5162 = _T_5034 & way_status_out_85; // @[Mux.scala 27:72]
  wire  _T_5289 = _T_5288 | _T_5162; // @[Mux.scala 27:72]
  wire  _T_5035 = ifu_ic_rw_int_addr_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_86; // @[Reg.scala 27:20]
  wire  _T_5163 = _T_5035 & way_status_out_86; // @[Mux.scala 27:72]
  wire  _T_5290 = _T_5289 | _T_5163; // @[Mux.scala 27:72]
  wire  _T_5036 = ifu_ic_rw_int_addr_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_87; // @[Reg.scala 27:20]
  wire  _T_5164 = _T_5036 & way_status_out_87; // @[Mux.scala 27:72]
  wire  _T_5291 = _T_5290 | _T_5164; // @[Mux.scala 27:72]
  wire  _T_5037 = ifu_ic_rw_int_addr_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_88; // @[Reg.scala 27:20]
  wire  _T_5165 = _T_5037 & way_status_out_88; // @[Mux.scala 27:72]
  wire  _T_5292 = _T_5291 | _T_5165; // @[Mux.scala 27:72]
  wire  _T_5038 = ifu_ic_rw_int_addr_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_89; // @[Reg.scala 27:20]
  wire  _T_5166 = _T_5038 & way_status_out_89; // @[Mux.scala 27:72]
  wire  _T_5293 = _T_5292 | _T_5166; // @[Mux.scala 27:72]
  wire  _T_5039 = ifu_ic_rw_int_addr_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_90; // @[Reg.scala 27:20]
  wire  _T_5167 = _T_5039 & way_status_out_90; // @[Mux.scala 27:72]
  wire  _T_5294 = _T_5293 | _T_5167; // @[Mux.scala 27:72]
  wire  _T_5040 = ifu_ic_rw_int_addr_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_91; // @[Reg.scala 27:20]
  wire  _T_5168 = _T_5040 & way_status_out_91; // @[Mux.scala 27:72]
  wire  _T_5295 = _T_5294 | _T_5168; // @[Mux.scala 27:72]
  wire  _T_5041 = ifu_ic_rw_int_addr_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_92; // @[Reg.scala 27:20]
  wire  _T_5169 = _T_5041 & way_status_out_92; // @[Mux.scala 27:72]
  wire  _T_5296 = _T_5295 | _T_5169; // @[Mux.scala 27:72]
  wire  _T_5042 = ifu_ic_rw_int_addr_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_93; // @[Reg.scala 27:20]
  wire  _T_5170 = _T_5042 & way_status_out_93; // @[Mux.scala 27:72]
  wire  _T_5297 = _T_5296 | _T_5170; // @[Mux.scala 27:72]
  wire  _T_5043 = ifu_ic_rw_int_addr_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_94; // @[Reg.scala 27:20]
  wire  _T_5171 = _T_5043 & way_status_out_94; // @[Mux.scala 27:72]
  wire  _T_5298 = _T_5297 | _T_5171; // @[Mux.scala 27:72]
  wire  _T_5044 = ifu_ic_rw_int_addr_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_95; // @[Reg.scala 27:20]
  wire  _T_5172 = _T_5044 & way_status_out_95; // @[Mux.scala 27:72]
  wire  _T_5299 = _T_5298 | _T_5172; // @[Mux.scala 27:72]
  wire  _T_5045 = ifu_ic_rw_int_addr_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_96; // @[Reg.scala 27:20]
  wire  _T_5173 = _T_5045 & way_status_out_96; // @[Mux.scala 27:72]
  wire  _T_5300 = _T_5299 | _T_5173; // @[Mux.scala 27:72]
  wire  _T_5046 = ifu_ic_rw_int_addr_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_97; // @[Reg.scala 27:20]
  wire  _T_5174 = _T_5046 & way_status_out_97; // @[Mux.scala 27:72]
  wire  _T_5301 = _T_5300 | _T_5174; // @[Mux.scala 27:72]
  wire  _T_5047 = ifu_ic_rw_int_addr_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_98; // @[Reg.scala 27:20]
  wire  _T_5175 = _T_5047 & way_status_out_98; // @[Mux.scala 27:72]
  wire  _T_5302 = _T_5301 | _T_5175; // @[Mux.scala 27:72]
  wire  _T_5048 = ifu_ic_rw_int_addr_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_99; // @[Reg.scala 27:20]
  wire  _T_5176 = _T_5048 & way_status_out_99; // @[Mux.scala 27:72]
  wire  _T_5303 = _T_5302 | _T_5176; // @[Mux.scala 27:72]
  wire  _T_5049 = ifu_ic_rw_int_addr_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_100; // @[Reg.scala 27:20]
  wire  _T_5177 = _T_5049 & way_status_out_100; // @[Mux.scala 27:72]
  wire  _T_5304 = _T_5303 | _T_5177; // @[Mux.scala 27:72]
  wire  _T_5050 = ifu_ic_rw_int_addr_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_101; // @[Reg.scala 27:20]
  wire  _T_5178 = _T_5050 & way_status_out_101; // @[Mux.scala 27:72]
  wire  _T_5305 = _T_5304 | _T_5178; // @[Mux.scala 27:72]
  wire  _T_5051 = ifu_ic_rw_int_addr_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_102; // @[Reg.scala 27:20]
  wire  _T_5179 = _T_5051 & way_status_out_102; // @[Mux.scala 27:72]
  wire  _T_5306 = _T_5305 | _T_5179; // @[Mux.scala 27:72]
  wire  _T_5052 = ifu_ic_rw_int_addr_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_103; // @[Reg.scala 27:20]
  wire  _T_5180 = _T_5052 & way_status_out_103; // @[Mux.scala 27:72]
  wire  _T_5307 = _T_5306 | _T_5180; // @[Mux.scala 27:72]
  wire  _T_5053 = ifu_ic_rw_int_addr_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_104; // @[Reg.scala 27:20]
  wire  _T_5181 = _T_5053 & way_status_out_104; // @[Mux.scala 27:72]
  wire  _T_5308 = _T_5307 | _T_5181; // @[Mux.scala 27:72]
  wire  _T_5054 = ifu_ic_rw_int_addr_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_105; // @[Reg.scala 27:20]
  wire  _T_5182 = _T_5054 & way_status_out_105; // @[Mux.scala 27:72]
  wire  _T_5309 = _T_5308 | _T_5182; // @[Mux.scala 27:72]
  wire  _T_5055 = ifu_ic_rw_int_addr_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_106; // @[Reg.scala 27:20]
  wire  _T_5183 = _T_5055 & way_status_out_106; // @[Mux.scala 27:72]
  wire  _T_5310 = _T_5309 | _T_5183; // @[Mux.scala 27:72]
  wire  _T_5056 = ifu_ic_rw_int_addr_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_107; // @[Reg.scala 27:20]
  wire  _T_5184 = _T_5056 & way_status_out_107; // @[Mux.scala 27:72]
  wire  _T_5311 = _T_5310 | _T_5184; // @[Mux.scala 27:72]
  wire  _T_5057 = ifu_ic_rw_int_addr_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_108; // @[Reg.scala 27:20]
  wire  _T_5185 = _T_5057 & way_status_out_108; // @[Mux.scala 27:72]
  wire  _T_5312 = _T_5311 | _T_5185; // @[Mux.scala 27:72]
  wire  _T_5058 = ifu_ic_rw_int_addr_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_109; // @[Reg.scala 27:20]
  wire  _T_5186 = _T_5058 & way_status_out_109; // @[Mux.scala 27:72]
  wire  _T_5313 = _T_5312 | _T_5186; // @[Mux.scala 27:72]
  wire  _T_5059 = ifu_ic_rw_int_addr_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_110; // @[Reg.scala 27:20]
  wire  _T_5187 = _T_5059 & way_status_out_110; // @[Mux.scala 27:72]
  wire  _T_5314 = _T_5313 | _T_5187; // @[Mux.scala 27:72]
  wire  _T_5060 = ifu_ic_rw_int_addr_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_111; // @[Reg.scala 27:20]
  wire  _T_5188 = _T_5060 & way_status_out_111; // @[Mux.scala 27:72]
  wire  _T_5315 = _T_5314 | _T_5188; // @[Mux.scala 27:72]
  wire  _T_5061 = ifu_ic_rw_int_addr_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_112; // @[Reg.scala 27:20]
  wire  _T_5189 = _T_5061 & way_status_out_112; // @[Mux.scala 27:72]
  wire  _T_5316 = _T_5315 | _T_5189; // @[Mux.scala 27:72]
  wire  _T_5062 = ifu_ic_rw_int_addr_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_113; // @[Reg.scala 27:20]
  wire  _T_5190 = _T_5062 & way_status_out_113; // @[Mux.scala 27:72]
  wire  _T_5317 = _T_5316 | _T_5190; // @[Mux.scala 27:72]
  wire  _T_5063 = ifu_ic_rw_int_addr_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_114; // @[Reg.scala 27:20]
  wire  _T_5191 = _T_5063 & way_status_out_114; // @[Mux.scala 27:72]
  wire  _T_5318 = _T_5317 | _T_5191; // @[Mux.scala 27:72]
  wire  _T_5064 = ifu_ic_rw_int_addr_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_115; // @[Reg.scala 27:20]
  wire  _T_5192 = _T_5064 & way_status_out_115; // @[Mux.scala 27:72]
  wire  _T_5319 = _T_5318 | _T_5192; // @[Mux.scala 27:72]
  wire  _T_5065 = ifu_ic_rw_int_addr_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_116; // @[Reg.scala 27:20]
  wire  _T_5193 = _T_5065 & way_status_out_116; // @[Mux.scala 27:72]
  wire  _T_5320 = _T_5319 | _T_5193; // @[Mux.scala 27:72]
  wire  _T_5066 = ifu_ic_rw_int_addr_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_117; // @[Reg.scala 27:20]
  wire  _T_5194 = _T_5066 & way_status_out_117; // @[Mux.scala 27:72]
  wire  _T_5321 = _T_5320 | _T_5194; // @[Mux.scala 27:72]
  wire  _T_5067 = ifu_ic_rw_int_addr_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_118; // @[Reg.scala 27:20]
  wire  _T_5195 = _T_5067 & way_status_out_118; // @[Mux.scala 27:72]
  wire  _T_5322 = _T_5321 | _T_5195; // @[Mux.scala 27:72]
  wire  _T_5068 = ifu_ic_rw_int_addr_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_119; // @[Reg.scala 27:20]
  wire  _T_5196 = _T_5068 & way_status_out_119; // @[Mux.scala 27:72]
  wire  _T_5323 = _T_5322 | _T_5196; // @[Mux.scala 27:72]
  wire  _T_5069 = ifu_ic_rw_int_addr_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_120; // @[Reg.scala 27:20]
  wire  _T_5197 = _T_5069 & way_status_out_120; // @[Mux.scala 27:72]
  wire  _T_5324 = _T_5323 | _T_5197; // @[Mux.scala 27:72]
  wire  _T_5070 = ifu_ic_rw_int_addr_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_121; // @[Reg.scala 27:20]
  wire  _T_5198 = _T_5070 & way_status_out_121; // @[Mux.scala 27:72]
  wire  _T_5325 = _T_5324 | _T_5198; // @[Mux.scala 27:72]
  wire  _T_5071 = ifu_ic_rw_int_addr_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_122; // @[Reg.scala 27:20]
  wire  _T_5199 = _T_5071 & way_status_out_122; // @[Mux.scala 27:72]
  wire  _T_5326 = _T_5325 | _T_5199; // @[Mux.scala 27:72]
  wire  _T_5072 = ifu_ic_rw_int_addr_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_123; // @[Reg.scala 27:20]
  wire  _T_5200 = _T_5072 & way_status_out_123; // @[Mux.scala 27:72]
  wire  _T_5327 = _T_5326 | _T_5200; // @[Mux.scala 27:72]
  wire  _T_5073 = ifu_ic_rw_int_addr_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_124; // @[Reg.scala 27:20]
  wire  _T_5201 = _T_5073 & way_status_out_124; // @[Mux.scala 27:72]
  wire  _T_5328 = _T_5327 | _T_5201; // @[Mux.scala 27:72]
  wire  _T_5074 = ifu_ic_rw_int_addr_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_125; // @[Reg.scala 27:20]
  wire  _T_5202 = _T_5074 & way_status_out_125; // @[Mux.scala 27:72]
  wire  _T_5329 = _T_5328 | _T_5202; // @[Mux.scala 27:72]
  wire  _T_5075 = ifu_ic_rw_int_addr_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_126; // @[Reg.scala 27:20]
  wire  _T_5203 = _T_5075 & way_status_out_126; // @[Mux.scala 27:72]
  wire  _T_5330 = _T_5329 | _T_5203; // @[Mux.scala 27:72]
  wire  _T_5076 = ifu_ic_rw_int_addr_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 730:80]
  reg  way_status_out_127; // @[Reg.scala 27:20]
  wire  _T_5204 = _T_5076 & way_status_out_127; // @[Mux.scala 27:72]
  wire  way_status = _T_5330 | _T_5204; // @[Mux.scala 27:72]
  wire  _T_195 = ~reset_all_tags; // @[el2_ifu_mem_ctl.scala 262:96]
  wire [1:0] _T_197 = _T_195 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_198 = _T_197 & io_ic_tag_valid; // @[el2_ifu_mem_ctl.scala 262:113]
  reg [1:0] tagv_mb_scnd_ff; // @[el2_ifu_mem_ctl.scala 268:29]
  reg  uncacheable_miss_scnd_ff; // @[el2_ifu_mem_ctl.scala 264:38]
  reg [30:0] imb_scnd_ff; // @[el2_ifu_mem_ctl.scala 266:25]
  wire [2:0] _T_206 = bus_ifu_wr_en_ff ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  reg [2:0] ifu_bus_rid_ff; // @[Reg.scala 27:20]
  wire [2:0] ic_wr_addr_bits_hi_3 = ifu_bus_rid_ff & _T_206; // @[el2_ifu_mem_ctl.scala 271:45]
  wire  _T_212 = _T_231 | _T_239; // @[el2_ifu_mem_ctl.scala 276:59]
  wire  _T_214 = _T_212 | _T_2233; // @[el2_ifu_mem_ctl.scala 276:91]
  wire  ic_iccm_hit_f = fetch_req_iccm_f & _T_214; // @[el2_ifu_mem_ctl.scala 276:41]
  wire  _T_219 = _T_227 & fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 282:39]
  wire  _T_221 = _T_219 & _T_195; // @[el2_ifu_mem_ctl.scala 282:60]
  wire  _T_225 = _T_221 & _T_212; // @[el2_ifu_mem_ctl.scala 282:78]
  wire  ic_act_hit_f = _T_225 & _T_247; // @[el2_ifu_mem_ctl.scala 282:126]
  wire  _T_262 = ic_act_hit_f | ic_byp_hit_f; // @[el2_ifu_mem_ctl.scala 289:31]
  wire  _T_263 = _T_262 | ic_iccm_hit_f; // @[el2_ifu_mem_ctl.scala 289:46]
  wire  _T_264 = ifc_region_acc_fault_final_f & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 289:94]
  wire  _T_268 = sel_hold_imb ? uncacheable_miss_ff : io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 290:84]
  wire  uncacheable_miss_in = scnd_miss_req ? uncacheable_miss_scnd_ff : _T_268; // @[el2_ifu_mem_ctl.scala 290:32]
  wire  _T_274 = imb_ff[11:5] == imb_scnd_ff[11:5]; // @[el2_ifu_mem_ctl.scala 293:79]
  wire  _T_275 = _T_274 & scnd_miss_req; // @[el2_ifu_mem_ctl.scala 293:135]
  reg [1:0] ifu_bus_rresp_ff; // @[Reg.scala 27:20]
  wire  _T_2662 = |ifu_bus_rresp_ff; // @[el2_ifu_mem_ctl.scala 621:48]
  wire  _T_2663 = _T_2662 & ifu_bus_rvalid_ff; // @[el2_ifu_mem_ctl.scala 621:52]
  wire  bus_ifu_wr_data_error_ff = _T_2663 & miss_pending; // @[el2_ifu_mem_ctl.scala 621:73]
  reg  ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 366:61]
  wire  ifu_wr_cumulative_err_data = bus_ifu_wr_data_error_ff | ifu_wr_data_comb_err_ff; // @[el2_ifu_mem_ctl.scala 365:55]
  wire  _T_276 = ~ifu_wr_cumulative_err_data; // @[el2_ifu_mem_ctl.scala 293:153]
  wire  scnd_miss_index_match = _T_275 & _T_276; // @[el2_ifu_mem_ctl.scala 293:151]
  wire  _T_277 = ~scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 296:47]
  wire  _T_278 = scnd_miss_req & _T_277; // @[el2_ifu_mem_ctl.scala 296:45]
  wire  _T_280 = scnd_miss_req & scnd_miss_index_match; // @[el2_ifu_mem_ctl.scala 297:26]
  reg  way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 316:30]
  wire  _T_10538 = ~way_status_mb_ff; // @[el2_ifu_mem_ctl.scala 786:33]
  reg [1:0] tagv_mb_ff; // @[el2_ifu_mem_ctl.scala 317:24]
  wire  _T_10540 = _T_10538 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:51]
  wire  _T_10542 = _T_10540 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 786:67]
  wire  _T_10544 = ~tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 786:86]
  wire  replace_way_mb_any_0 = _T_10542 | _T_10544; // @[el2_ifu_mem_ctl.scala 786:84]
  wire [1:0] _T_287 = scnd_miss_index_match ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10547 = way_status_mb_ff & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 787:50]
  wire  _T_10549 = _T_10547 & tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 787:66]
  wire  _T_10551 = ~tagv_mb_ff[1]; // @[el2_ifu_mem_ctl.scala 787:85]
  wire  _T_10553 = _T_10551 & tagv_mb_ff[0]; // @[el2_ifu_mem_ctl.scala 787:100]
  wire  replace_way_mb_any_1 = _T_10549 | _T_10553; // @[el2_ifu_mem_ctl.scala 787:83]
  wire [1:0] _T_288 = {replace_way_mb_any_1,replace_way_mb_any_0}; // @[Cat.scala 29:58]
  wire [1:0] _T_289 = _T_287 & _T_288; // @[el2_ifu_mem_ctl.scala 301:110]
  wire [1:0] _T_290 = tagv_mb_scnd_ff | _T_289; // @[el2_ifu_mem_ctl.scala 301:62]
  wire [1:0] _T_295 = io_ic_tag_valid & _T_197; // @[el2_ifu_mem_ctl.scala 302:56]
  wire  _T_297 = ~scnd_miss_req_q; // @[el2_ifu_mem_ctl.scala 305:36]
  wire  _T_298 = miss_pending & _T_297; // @[el2_ifu_mem_ctl.scala 305:34]
  reg  reset_ic_ff; // @[el2_ifu_mem_ctl.scala 306:25]
  wire  _T_299 = reset_all_tags | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 305:72]
  wire  reset_ic_in = _T_298 & _T_299; // @[el2_ifu_mem_ctl.scala 305:53]
  reg  fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 307:37]
  reg [25:0] miss_addr; // @[el2_ifu_mem_ctl.scala 315:23]
  wire  _T_313 = _T_2248 & flush_final_f; // @[el2_ifu_mem_ctl.scala 319:87]
  wire  _T_314 = ~_T_313; // @[el2_ifu_mem_ctl.scala 319:55]
  wire  _T_315 = io_ifc_fetch_req_bf & _T_314; // @[el2_ifu_mem_ctl.scala 319:53]
  wire  _T_2240 = ~_T_2235; // @[el2_ifu_mem_ctl.scala 456:46]
  wire  _T_2241 = _T_2233 & _T_2240; // @[el2_ifu_mem_ctl.scala 456:44]
  wire  stream_miss_f = _T_2241 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 456:84]
  wire  _T_316 = ~stream_miss_f; // @[el2_ifu_mem_ctl.scala 319:106]
  wire  ifc_fetch_req_qual_bf = _T_315 & _T_316; // @[el2_ifu_mem_ctl.scala 319:104]
  reg  ifc_region_acc_fault_f; // @[el2_ifu_mem_ctl.scala 325:39]
  reg [2:0] bus_rd_addr_count; // @[Reg.scala 27:20]
  wire [28:0] ifu_ic_req_addr_f = {miss_addr,bus_rd_addr_count}; // @[Cat.scala 29:58]
  wire  _T_323 = _T_239 | _T_2233; // @[el2_ifu_mem_ctl.scala 327:55]
  wire  _T_326 = _T_323 & _T_56; // @[el2_ifu_mem_ctl.scala 327:82]
  wire  _T_2254 = ~ifu_bus_rid_ff[0]; // @[el2_ifu_mem_ctl.scala 461:55]
  wire [2:0] other_tag = {ifu_bus_rid_ff[2:1],_T_2254}; // @[Cat.scala 29:58]
  wire  _T_2255 = other_tag == 3'h0; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2279 = _T_2255 & ic_miss_buff_data_valid[0]; // @[Mux.scala 27:72]
  wire  _T_2258 = other_tag == 3'h1; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2280 = _T_2258 & ic_miss_buff_data_valid[1]; // @[Mux.scala 27:72]
  wire  _T_2287 = _T_2279 | _T_2280; // @[Mux.scala 27:72]
  wire  _T_2261 = other_tag == 3'h2; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2281 = _T_2261 & ic_miss_buff_data_valid[2]; // @[Mux.scala 27:72]
  wire  _T_2288 = _T_2287 | _T_2281; // @[Mux.scala 27:72]
  wire  _T_2264 = other_tag == 3'h3; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2282 = _T_2264 & ic_miss_buff_data_valid[3]; // @[Mux.scala 27:72]
  wire  _T_2289 = _T_2288 | _T_2282; // @[Mux.scala 27:72]
  wire  _T_2267 = other_tag == 3'h4; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2283 = _T_2267 & ic_miss_buff_data_valid[4]; // @[Mux.scala 27:72]
  wire  _T_2290 = _T_2289 | _T_2283; // @[Mux.scala 27:72]
  wire  _T_2270 = other_tag == 3'h5; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2284 = _T_2270 & ic_miss_buff_data_valid[5]; // @[Mux.scala 27:72]
  wire  _T_2291 = _T_2290 | _T_2284; // @[Mux.scala 27:72]
  wire  _T_2273 = other_tag == 3'h6; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2285 = _T_2273 & ic_miss_buff_data_valid[6]; // @[Mux.scala 27:72]
  wire  _T_2292 = _T_2291 | _T_2285; // @[Mux.scala 27:72]
  wire  _T_2276 = other_tag == 3'h7; // @[el2_ifu_mem_ctl.scala 462:81]
  wire  _T_2286 = _T_2276 & ic_miss_buff_data_valid[7]; // @[Mux.scala 27:72]
  wire  second_half_available = _T_2292 | _T_2286; // @[Mux.scala 27:72]
  wire  write_ic_16_bytes = second_half_available & bus_ifu_wr_en_ff; // @[el2_ifu_mem_ctl.scala 463:46]
  wire  _T_330 = miss_pending & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 331:35]
  wire  _T_332 = _T_330 & _T_17; // @[el2_ifu_mem_ctl.scala 331:55]
  reg  ic_act_miss_f_delayed; // @[el2_ifu_mem_ctl.scala 618:61]
  wire  _T_2656 = ic_act_miss_f_delayed & _T_2249; // @[el2_ifu_mem_ctl.scala 619:53]
  wire  reset_tag_valid_for_miss = _T_2656 & _T_17; // @[el2_ifu_mem_ctl.scala 619:84]
  wire  sel_mb_addr = _T_332 | reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 331:79]
  wire [30:0] _T_336 = {imb_ff[30:5],ic_wr_addr_bits_hi_3,imb_ff[1:0]}; // @[Cat.scala 29:58]
  wire  _T_337 = ~sel_mb_addr; // @[el2_ifu_mem_ctl.scala 333:37]
  wire [30:0] _T_338 = sel_mb_addr ? _T_336 : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] _T_339 = _T_337 ? io_ifc_fetch_addr_bf : 31'h0; // @[Mux.scala 27:72]
  wire [30:0] ifu_ic_rw_int_addr = _T_338 | _T_339; // @[Mux.scala 27:72]
  wire  _T_344 = _T_332 & last_beat; // @[el2_ifu_mem_ctl.scala 335:84]
  wire  _T_2650 = ~_T_2662; // @[el2_ifu_mem_ctl.scala 616:84]
  wire  _T_2651 = _T_100 & _T_2650; // @[el2_ifu_mem_ctl.scala 616:82]
  wire  bus_ifu_wr_en_ff_q = _T_2651 & write_ic_16_bytes; // @[el2_ifu_mem_ctl.scala 616:108]
  wire  sel_mb_status_addr = _T_344 & bus_ifu_wr_en_ff_q; // @[el2_ifu_mem_ctl.scala 335:96]
  wire [30:0] ifu_status_wr_addr = sel_mb_status_addr ? _T_336 : ifu_fetch_addr_int_f; // @[el2_ifu_mem_ctl.scala 336:31]
  reg [63:0] ifu_bus_rdata_ff; // @[Reg.scala 27:20]
  wire [6:0] _T_567 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[57]}; // @[el2_lib.scala 401:13]
  wire  _T_568 = ^_T_567; // @[el2_lib.scala 401:20]
  wire [6:0] _T_574 = {ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31],ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[26]}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_581 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33]}; // @[el2_lib.scala 401:30]
  wire [14:0] _T_582 = {ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[33],_T_574}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_589 = {ifu_bus_rdata_ff[48],ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[41]}; // @[el2_lib.scala 401:30]
  wire [30:0] _T_598 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_582}; // @[el2_lib.scala 401:30]
  wire  _T_599 = ^_T_598; // @[el2_lib.scala 401:37]
  wire [6:0] _T_605 = {ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[13],ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[11]}; // @[el2_lib.scala 401:47]
  wire [14:0] _T_613 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_605}; // @[el2_lib.scala 401:47]
  wire [30:0] _T_629 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_589,_T_613}; // @[el2_lib.scala 401:47]
  wire  _T_630 = ^_T_629; // @[el2_lib.scala 401:54]
  wire [6:0] _T_636 = {ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[4]}; // @[el2_lib.scala 401:64]
  wire [14:0] _T_644 = {ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[18],_T_636}; // @[el2_lib.scala 401:64]
  wire [30:0] _T_660 = {ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[49],_T_581,_T_644}; // @[el2_lib.scala 401:64]
  wire  _T_661 = ^_T_660; // @[el2_lib.scala 401:71]
  wire [7:0] _T_668 = {ifu_bus_rdata_ff[14],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[7],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[1]}; // @[el2_lib.scala 401:81]
  wire [16:0] _T_677 = {ifu_bus_rdata_ff[30],ifu_bus_rdata_ff[29],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[22],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[15],_T_668}; // @[el2_lib.scala 401:81]
  wire [8:0] _T_685 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[45],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[37],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 401:81]
  wire [17:0] _T_694 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[60],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[53],ifu_bus_rdata_ff[48],_T_685}; // @[el2_lib.scala 401:81]
  wire [34:0] _T_695 = {_T_694,_T_677}; // @[el2_lib.scala 401:81]
  wire  _T_696 = ^_T_695; // @[el2_lib.scala 401:88]
  wire [7:0] _T_703 = {ifu_bus_rdata_ff[12],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[9],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[5],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[2],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 401:98]
  wire [16:0] _T_712 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[27],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[24],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[20],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[16],ifu_bus_rdata_ff[13],_T_703}; // @[el2_lib.scala 401:98]
  wire [8:0] _T_720 = {ifu_bus_rdata_ff[47],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[43],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[39],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[35],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[31]}; // @[el2_lib.scala 401:98]
  wire [17:0] _T_729 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[62],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[58],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[55],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[51],ifu_bus_rdata_ff[48],_T_720}; // @[el2_lib.scala 401:98]
  wire [34:0] _T_730 = {_T_729,_T_712}; // @[el2_lib.scala 401:98]
  wire  _T_731 = ^_T_730; // @[el2_lib.scala 401:105]
  wire [7:0] _T_738 = {ifu_bus_rdata_ff[11],ifu_bus_rdata_ff[10],ifu_bus_rdata_ff[8],ifu_bus_rdata_ff[6],ifu_bus_rdata_ff[4],ifu_bus_rdata_ff[3],ifu_bus_rdata_ff[1],ifu_bus_rdata_ff[0]}; // @[el2_lib.scala 401:115]
  wire [16:0] _T_747 = {ifu_bus_rdata_ff[28],ifu_bus_rdata_ff[26],ifu_bus_rdata_ff[25],ifu_bus_rdata_ff[23],ifu_bus_rdata_ff[21],ifu_bus_rdata_ff[19],ifu_bus_rdata_ff[17],ifu_bus_rdata_ff[15],ifu_bus_rdata_ff[13],_T_738}; // @[el2_lib.scala 401:115]
  wire [8:0] _T_755 = {ifu_bus_rdata_ff[46],ifu_bus_rdata_ff[44],ifu_bus_rdata_ff[42],ifu_bus_rdata_ff[40],ifu_bus_rdata_ff[38],ifu_bus_rdata_ff[36],ifu_bus_rdata_ff[34],ifu_bus_rdata_ff[32],ifu_bus_rdata_ff[30]}; // @[el2_lib.scala 401:115]
  wire [17:0] _T_764 = {ifu_bus_rdata_ff[63],ifu_bus_rdata_ff[61],ifu_bus_rdata_ff[59],ifu_bus_rdata_ff[57],ifu_bus_rdata_ff[56],ifu_bus_rdata_ff[54],ifu_bus_rdata_ff[52],ifu_bus_rdata_ff[50],ifu_bus_rdata_ff[48],_T_755}; // @[el2_lib.scala 401:115]
  wire [34:0] _T_765 = {_T_764,_T_747}; // @[el2_lib.scala 401:115]
  wire  _T_766 = ^_T_765; // @[el2_lib.scala 401:122]
  wire [3:0] _T_2295 = {ifu_bus_rid_ff[2:1],_T_2254,1'h1}; // @[Cat.scala 29:58]
  wire  _T_2296 = _T_2295 == 4'h0; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_0; // @[Reg.scala 27:20]
  wire [31:0] _T_2343 = _T_2296 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2299 = _T_2295 == 4'h1; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_1; // @[Reg.scala 27:20]
  wire [31:0] _T_2344 = _T_2299 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2359 = _T_2343 | _T_2344; // @[Mux.scala 27:72]
  wire  _T_2302 = _T_2295 == 4'h2; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_2; // @[Reg.scala 27:20]
  wire [31:0] _T_2345 = _T_2302 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2360 = _T_2359 | _T_2345; // @[Mux.scala 27:72]
  wire  _T_2305 = _T_2295 == 4'h3; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_3; // @[Reg.scala 27:20]
  wire [31:0] _T_2346 = _T_2305 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2361 = _T_2360 | _T_2346; // @[Mux.scala 27:72]
  wire  _T_2308 = _T_2295 == 4'h4; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_4; // @[Reg.scala 27:20]
  wire [31:0] _T_2347 = _T_2308 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2362 = _T_2361 | _T_2347; // @[Mux.scala 27:72]
  wire  _T_2311 = _T_2295 == 4'h5; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_5; // @[Reg.scala 27:20]
  wire [31:0] _T_2348 = _T_2311 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2363 = _T_2362 | _T_2348; // @[Mux.scala 27:72]
  wire  _T_2314 = _T_2295 == 4'h6; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_6; // @[Reg.scala 27:20]
  wire [31:0] _T_2349 = _T_2314 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2364 = _T_2363 | _T_2349; // @[Mux.scala 27:72]
  wire  _T_2317 = _T_2295 == 4'h7; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_7; // @[Reg.scala 27:20]
  wire [31:0] _T_2350 = _T_2317 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2365 = _T_2364 | _T_2350; // @[Mux.scala 27:72]
  wire  _T_2320 = _T_2295 == 4'h8; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_8; // @[Reg.scala 27:20]
  wire [31:0] _T_2351 = _T_2320 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2366 = _T_2365 | _T_2351; // @[Mux.scala 27:72]
  wire  _T_2323 = _T_2295 == 4'h9; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_9; // @[Reg.scala 27:20]
  wire [31:0] _T_2352 = _T_2323 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2367 = _T_2366 | _T_2352; // @[Mux.scala 27:72]
  wire  _T_2326 = _T_2295 == 4'ha; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_10; // @[Reg.scala 27:20]
  wire [31:0] _T_2353 = _T_2326 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2368 = _T_2367 | _T_2353; // @[Mux.scala 27:72]
  wire  _T_2329 = _T_2295 == 4'hb; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_11; // @[Reg.scala 27:20]
  wire [31:0] _T_2354 = _T_2329 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2369 = _T_2368 | _T_2354; // @[Mux.scala 27:72]
  wire  _T_2332 = _T_2295 == 4'hc; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_12; // @[Reg.scala 27:20]
  wire [31:0] _T_2355 = _T_2332 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2370 = _T_2369 | _T_2355; // @[Mux.scala 27:72]
  wire  _T_2335 = _T_2295 == 4'hd; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_13; // @[Reg.scala 27:20]
  wire [31:0] _T_2356 = _T_2335 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2371 = _T_2370 | _T_2356; // @[Mux.scala 27:72]
  wire  _T_2338 = _T_2295 == 4'he; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_14; // @[Reg.scala 27:20]
  wire [31:0] _T_2357 = _T_2338 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2372 = _T_2371 | _T_2357; // @[Mux.scala 27:72]
  wire  _T_2341 = _T_2295 == 4'hf; // @[el2_ifu_mem_ctl.scala 464:89]
  reg [31:0] ic_miss_buff_data_15; // @[Reg.scala 27:20]
  wire [31:0] _T_2358 = _T_2341 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2373 = _T_2372 | _T_2358; // @[Mux.scala 27:72]
  wire [3:0] _T_2375 = {ifu_bus_rid_ff[2:1],_T_2254,1'h0}; // @[Cat.scala 29:58]
  wire  _T_2376 = _T_2375 == 4'h0; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2423 = _T_2376 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_2379 = _T_2375 == 4'h1; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2424 = _T_2379 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2439 = _T_2423 | _T_2424; // @[Mux.scala 27:72]
  wire  _T_2382 = _T_2375 == 4'h2; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2425 = _T_2382 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2440 = _T_2439 | _T_2425; // @[Mux.scala 27:72]
  wire  _T_2385 = _T_2375 == 4'h3; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2426 = _T_2385 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2441 = _T_2440 | _T_2426; // @[Mux.scala 27:72]
  wire  _T_2388 = _T_2375 == 4'h4; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2427 = _T_2388 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2442 = _T_2441 | _T_2427; // @[Mux.scala 27:72]
  wire  _T_2391 = _T_2375 == 4'h5; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2428 = _T_2391 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2443 = _T_2442 | _T_2428; // @[Mux.scala 27:72]
  wire  _T_2394 = _T_2375 == 4'h6; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2429 = _T_2394 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2444 = _T_2443 | _T_2429; // @[Mux.scala 27:72]
  wire  _T_2397 = _T_2375 == 4'h7; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2430 = _T_2397 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2445 = _T_2444 | _T_2430; // @[Mux.scala 27:72]
  wire  _T_2400 = _T_2375 == 4'h8; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2431 = _T_2400 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2446 = _T_2445 | _T_2431; // @[Mux.scala 27:72]
  wire  _T_2403 = _T_2375 == 4'h9; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2432 = _T_2403 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2447 = _T_2446 | _T_2432; // @[Mux.scala 27:72]
  wire  _T_2406 = _T_2375 == 4'ha; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2433 = _T_2406 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2448 = _T_2447 | _T_2433; // @[Mux.scala 27:72]
  wire  _T_2409 = _T_2375 == 4'hb; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2434 = _T_2409 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2449 = _T_2448 | _T_2434; // @[Mux.scala 27:72]
  wire  _T_2412 = _T_2375 == 4'hc; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2435 = _T_2412 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2450 = _T_2449 | _T_2435; // @[Mux.scala 27:72]
  wire  _T_2415 = _T_2375 == 4'hd; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2436 = _T_2415 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2451 = _T_2450 | _T_2436; // @[Mux.scala 27:72]
  wire  _T_2418 = _T_2375 == 4'he; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2437 = _T_2418 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2452 = _T_2451 | _T_2437; // @[Mux.scala 27:72]
  wire  _T_2421 = _T_2375 == 4'hf; // @[el2_ifu_mem_ctl.scala 465:66]
  wire [31:0] _T_2438 = _T_2421 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2453 = _T_2452 | _T_2438; // @[Mux.scala 27:72]
  wire [63:0] ic_miss_buff_half = {_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [6:0] _T_989 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[57]}; // @[el2_lib.scala 401:13]
  wire  _T_990 = ^_T_989; // @[el2_lib.scala 401:20]
  wire [6:0] _T_996 = {ic_miss_buff_half[32],ic_miss_buff_half[31],ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[26]}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_1003 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33]}; // @[el2_lib.scala 401:30]
  wire [14:0] _T_1004 = {ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[34],ic_miss_buff_half[33],_T_996}; // @[el2_lib.scala 401:30]
  wire [7:0] _T_1011 = {ic_miss_buff_half[48],ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[42],ic_miss_buff_half[41]}; // @[el2_lib.scala 401:30]
  wire [30:0] _T_1020 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1004}; // @[el2_lib.scala 401:30]
  wire  _T_1021 = ^_T_1020; // @[el2_lib.scala 401:37]
  wire [6:0] _T_1027 = {ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],ic_miss_buff_half[14],ic_miss_buff_half[13],ic_miss_buff_half[12],ic_miss_buff_half[11]}; // @[el2_lib.scala 401:47]
  wire [14:0] _T_1035 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1027}; // @[el2_lib.scala 401:47]
  wire [30:0] _T_1051 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1011,_T_1035}; // @[el2_lib.scala 401:47]
  wire  _T_1052 = ^_T_1051; // @[el2_lib.scala 401:54]
  wire [6:0] _T_1058 = {ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[4]}; // @[el2_lib.scala 401:64]
  wire [14:0] _T_1066 = {ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[19],ic_miss_buff_half[18],_T_1058}; // @[el2_lib.scala 401:64]
  wire [30:0] _T_1082 = {ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[50],ic_miss_buff_half[49],_T_1003,_T_1066}; // @[el2_lib.scala 401:64]
  wire  _T_1083 = ^_T_1082; // @[el2_lib.scala 401:71]
  wire [7:0] _T_1090 = {ic_miss_buff_half[14],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[8],ic_miss_buff_half[7],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[1]}; // @[el2_lib.scala 401:81]
  wire [16:0] _T_1099 = {ic_miss_buff_half[30],ic_miss_buff_half[29],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[23],ic_miss_buff_half[22],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[15],_T_1090}; // @[el2_lib.scala 401:81]
  wire [8:0] _T_1107 = {ic_miss_buff_half[47],ic_miss_buff_half[46],ic_miss_buff_half[45],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[38],ic_miss_buff_half[37],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 401:81]
  wire [17:0] _T_1116 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[61],ic_miss_buff_half[60],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[54],ic_miss_buff_half[53],ic_miss_buff_half[48],_T_1107}; // @[el2_lib.scala 401:81]
  wire [34:0] _T_1117 = {_T_1116,_T_1099}; // @[el2_lib.scala 401:81]
  wire  _T_1118 = ^_T_1117; // @[el2_lib.scala 401:88]
  wire [7:0] _T_1125 = {ic_miss_buff_half[12],ic_miss_buff_half[10],ic_miss_buff_half[9],ic_miss_buff_half[6],ic_miss_buff_half[5],ic_miss_buff_half[3],ic_miss_buff_half[2],ic_miss_buff_half[0]}; // @[el2_lib.scala 401:98]
  wire [16:0] _T_1134 = {ic_miss_buff_half[28],ic_miss_buff_half[27],ic_miss_buff_half[25],ic_miss_buff_half[24],ic_miss_buff_half[21],ic_miss_buff_half[20],ic_miss_buff_half[17],ic_miss_buff_half[16],ic_miss_buff_half[13],_T_1125}; // @[el2_lib.scala 401:98]
  wire [8:0] _T_1142 = {ic_miss_buff_half[47],ic_miss_buff_half[44],ic_miss_buff_half[43],ic_miss_buff_half[40],ic_miss_buff_half[39],ic_miss_buff_half[36],ic_miss_buff_half[35],ic_miss_buff_half[32],ic_miss_buff_half[31]}; // @[el2_lib.scala 401:98]
  wire [17:0] _T_1151 = {ic_miss_buff_half[63],ic_miss_buff_half[62],ic_miss_buff_half[59],ic_miss_buff_half[58],ic_miss_buff_half[56],ic_miss_buff_half[55],ic_miss_buff_half[52],ic_miss_buff_half[51],ic_miss_buff_half[48],_T_1142}; // @[el2_lib.scala 401:98]
  wire [34:0] _T_1152 = {_T_1151,_T_1134}; // @[el2_lib.scala 401:98]
  wire  _T_1153 = ^_T_1152; // @[el2_lib.scala 401:105]
  wire [7:0] _T_1160 = {ic_miss_buff_half[11],ic_miss_buff_half[10],ic_miss_buff_half[8],ic_miss_buff_half[6],ic_miss_buff_half[4],ic_miss_buff_half[3],ic_miss_buff_half[1],ic_miss_buff_half[0]}; // @[el2_lib.scala 401:115]
  wire [16:0] _T_1169 = {ic_miss_buff_half[28],ic_miss_buff_half[26],ic_miss_buff_half[25],ic_miss_buff_half[23],ic_miss_buff_half[21],ic_miss_buff_half[19],ic_miss_buff_half[17],ic_miss_buff_half[15],ic_miss_buff_half[13],_T_1160}; // @[el2_lib.scala 401:115]
  wire [8:0] _T_1177 = {ic_miss_buff_half[46],ic_miss_buff_half[44],ic_miss_buff_half[42],ic_miss_buff_half[40],ic_miss_buff_half[38],ic_miss_buff_half[36],ic_miss_buff_half[34],ic_miss_buff_half[32],ic_miss_buff_half[30]}; // @[el2_lib.scala 401:115]
  wire [17:0] _T_1186 = {ic_miss_buff_half[63],ic_miss_buff_half[61],ic_miss_buff_half[59],ic_miss_buff_half[57],ic_miss_buff_half[56],ic_miss_buff_half[54],ic_miss_buff_half[52],ic_miss_buff_half[50],ic_miss_buff_half[48],_T_1177}; // @[el2_lib.scala 401:115]
  wire [34:0] _T_1187 = {_T_1186,_T_1169}; // @[el2_lib.scala 401:115]
  wire  _T_1188 = ^_T_1187; // @[el2_lib.scala 401:122]
  wire [70:0] _T_1233 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff}; // @[Cat.scala 29:58]
  wire [70:0] _T_1232 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453}; // @[Cat.scala 29:58]
  wire [141:0] _T_1234 = {_T_568,_T_599,_T_630,_T_661,_T_696,_T_731,_T_766,ifu_bus_rdata_ff,_T_1232}; // @[Cat.scala 29:58]
  wire [141:0] _T_1237 = {_T_990,_T_1021,_T_1052,_T_1083,_T_1118,_T_1153,_T_1188,_T_2373,_T_2453,_T_1233}; // @[Cat.scala 29:58]
  wire [141:0] ic_wr_16bytes_data = ifu_bus_rid_ff[0] ? _T_1234 : _T_1237; // @[el2_ifu_mem_ctl.scala 357:28]
  wire  _T_1196 = |io_ic_eccerr; // @[el2_ifu_mem_ctl.scala 347:56]
  wire  _T_1197 = _T_1196 & ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 347:83]
  wire [4:0] bypass_index = imb_ff[4:0]; // @[el2_ifu_mem_ctl.scala 411:28]
  wire  _T_1413 = bypass_index[4:2] == 3'h0; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  bus_ifu_wr_en = _T_13 & miss_pending; // @[el2_ifu_mem_ctl.scala 614:35]
  wire  _T_1282 = io_ifu_axi_rid == 3'h0; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_0 = bus_ifu_wr_en & _T_1282; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1339 = ~ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 402:118]
  wire  _T_1340 = ic_miss_buff_data_valid[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_0 = write_fill_data_0 | _T_1340; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1436 = _T_1413 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1416 = bypass_index[4:2] == 3'h1; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1283 = io_ifu_axi_rid == 3'h1; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_1 = bus_ifu_wr_en & _T_1283; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1343 = ic_miss_buff_data_valid[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_1 = write_fill_data_1 | _T_1343; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1437 = _T_1416 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1444 = _T_1436 | _T_1437; // @[Mux.scala 27:72]
  wire  _T_1419 = bypass_index[4:2] == 3'h2; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1284 = io_ifu_axi_rid == 3'h2; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_2 = bus_ifu_wr_en & _T_1284; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1346 = ic_miss_buff_data_valid[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_2 = write_fill_data_2 | _T_1346; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1438 = _T_1419 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1445 = _T_1444 | _T_1438; // @[Mux.scala 27:72]
  wire  _T_1422 = bypass_index[4:2] == 3'h3; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1285 = io_ifu_axi_rid == 3'h3; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_3 = bus_ifu_wr_en & _T_1285; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1349 = ic_miss_buff_data_valid[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_3 = write_fill_data_3 | _T_1349; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1439 = _T_1422 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1446 = _T_1445 | _T_1439; // @[Mux.scala 27:72]
  wire  _T_1425 = bypass_index[4:2] == 3'h4; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1286 = io_ifu_axi_rid == 3'h4; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_4 = bus_ifu_wr_en & _T_1286; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1352 = ic_miss_buff_data_valid[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_4 = write_fill_data_4 | _T_1352; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1440 = _T_1425 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1447 = _T_1446 | _T_1440; // @[Mux.scala 27:72]
  wire  _T_1428 = bypass_index[4:2] == 3'h5; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1287 = io_ifu_axi_rid == 3'h5; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_5 = bus_ifu_wr_en & _T_1287; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1355 = ic_miss_buff_data_valid[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_5 = write_fill_data_5 | _T_1355; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1441 = _T_1428 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1448 = _T_1447 | _T_1441; // @[Mux.scala 27:72]
  wire  _T_1431 = bypass_index[4:2] == 3'h6; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1288 = io_ifu_axi_rid == 3'h6; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_6 = bus_ifu_wr_en & _T_1288; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1358 = ic_miss_buff_data_valid[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_6 = write_fill_data_6 | _T_1358; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1442 = _T_1431 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1449 = _T_1448 | _T_1442; // @[Mux.scala 27:72]
  wire  _T_1434 = bypass_index[4:2] == 3'h7; // @[el2_ifu_mem_ctl.scala 413:114]
  wire  _T_1289 = io_ifu_axi_rid == 3'h7; // @[el2_ifu_mem_ctl.scala 396:91]
  wire  write_fill_data_7 = bus_ifu_wr_en & _T_1289; // @[el2_ifu_mem_ctl.scala 396:73]
  wire  _T_1361 = ic_miss_buff_data_valid[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 402:116]
  wire  ic_miss_buff_data_valid_in_7 = write_fill_data_7 | _T_1361; // @[el2_ifu_mem_ctl.scala 402:88]
  wire  _T_1443 = _T_1434 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  bypass_valid_value_check = _T_1449 | _T_1443; // @[Mux.scala 27:72]
  wire  _T_1452 = ~bypass_index[1]; // @[el2_ifu_mem_ctl.scala 414:58]
  wire  _T_1453 = bypass_valid_value_check & _T_1452; // @[el2_ifu_mem_ctl.scala 414:56]
  wire  _T_1455 = ~bypass_index[0]; // @[el2_ifu_mem_ctl.scala 414:77]
  wire  _T_1456 = _T_1453 & _T_1455; // @[el2_ifu_mem_ctl.scala 414:75]
  wire  _T_1461 = _T_1453 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 415:75]
  wire  _T_1462 = _T_1456 | _T_1461; // @[el2_ifu_mem_ctl.scala 414:95]
  wire  _T_1464 = bypass_valid_value_check & bypass_index[1]; // @[el2_ifu_mem_ctl.scala 416:56]
  wire  _T_1467 = _T_1464 & _T_1455; // @[el2_ifu_mem_ctl.scala 416:74]
  wire  _T_1468 = _T_1462 | _T_1467; // @[el2_ifu_mem_ctl.scala 415:94]
  wire  _T_1472 = _T_1464 & bypass_index[0]; // @[el2_ifu_mem_ctl.scala 417:51]
  wire [2:0] bypass_index_5_3_inc = bypass_index[4:2] + 3'h1; // @[el2_ifu_mem_ctl.scala 412:70]
  wire  _T_1473 = bypass_index_5_3_inc == 3'h0; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1489 = _T_1473 & ic_miss_buff_data_valid_in_0; // @[Mux.scala 27:72]
  wire  _T_1475 = bypass_index_5_3_inc == 3'h1; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1490 = _T_1475 & ic_miss_buff_data_valid_in_1; // @[Mux.scala 27:72]
  wire  _T_1497 = _T_1489 | _T_1490; // @[Mux.scala 27:72]
  wire  _T_1477 = bypass_index_5_3_inc == 3'h2; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1491 = _T_1477 & ic_miss_buff_data_valid_in_2; // @[Mux.scala 27:72]
  wire  _T_1498 = _T_1497 | _T_1491; // @[Mux.scala 27:72]
  wire  _T_1479 = bypass_index_5_3_inc == 3'h3; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1492 = _T_1479 & ic_miss_buff_data_valid_in_3; // @[Mux.scala 27:72]
  wire  _T_1499 = _T_1498 | _T_1492; // @[Mux.scala 27:72]
  wire  _T_1481 = bypass_index_5_3_inc == 3'h4; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1493 = _T_1481 & ic_miss_buff_data_valid_in_4; // @[Mux.scala 27:72]
  wire  _T_1500 = _T_1499 | _T_1493; // @[Mux.scala 27:72]
  wire  _T_1483 = bypass_index_5_3_inc == 3'h5; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1494 = _T_1483 & ic_miss_buff_data_valid_in_5; // @[Mux.scala 27:72]
  wire  _T_1501 = _T_1500 | _T_1494; // @[Mux.scala 27:72]
  wire  _T_1485 = bypass_index_5_3_inc == 3'h6; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1495 = _T_1485 & ic_miss_buff_data_valid_in_6; // @[Mux.scala 27:72]
  wire  _T_1502 = _T_1501 | _T_1495; // @[Mux.scala 27:72]
  wire  _T_1487 = bypass_index_5_3_inc == 3'h7; // @[el2_ifu_mem_ctl.scala 417:132]
  wire  _T_1496 = _T_1487 & ic_miss_buff_data_valid_in_7; // @[Mux.scala 27:72]
  wire  _T_1503 = _T_1502 | _T_1496; // @[Mux.scala 27:72]
  wire  _T_1505 = _T_1472 & _T_1503; // @[el2_ifu_mem_ctl.scala 417:69]
  wire  _T_1506 = _T_1468 | _T_1505; // @[el2_ifu_mem_ctl.scala 416:94]
  wire [4:0] _GEN_473 = {{2'd0}, bypass_index[4:2]}; // @[el2_ifu_mem_ctl.scala 418:95]
  wire  _T_1509 = _GEN_473 == 5'h1f; // @[el2_ifu_mem_ctl.scala 418:95]
  wire  _T_1510 = bypass_valid_value_check & _T_1509; // @[el2_ifu_mem_ctl.scala 418:56]
  wire  bypass_data_ready_in = _T_1506 | _T_1510; // @[el2_ifu_mem_ctl.scala 417:181]
  wire  _T_1511 = bypass_data_ready_in & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 422:53]
  wire  _T_1512 = _T_1511 & uncacheable_miss_ff; // @[el2_ifu_mem_ctl.scala 422:73]
  wire  _T_1514 = _T_1512 & _T_317; // @[el2_ifu_mem_ctl.scala 422:96]
  wire  _T_1516 = _T_1514 & _T_58; // @[el2_ifu_mem_ctl.scala 422:118]
  wire  _T_1518 = crit_wd_byp_ok_ff & _T_17; // @[el2_ifu_mem_ctl.scala 423:73]
  wire  _T_1520 = _T_1518 & _T_317; // @[el2_ifu_mem_ctl.scala 423:96]
  wire  _T_1522 = _T_1520 & _T_58; // @[el2_ifu_mem_ctl.scala 423:118]
  wire  _T_1523 = _T_1516 | _T_1522; // @[el2_ifu_mem_ctl.scala 422:143]
  reg  ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 425:58]
  wire  _T_1524 = ic_crit_wd_rdy_new_ff & crit_wd_byp_ok_ff; // @[el2_ifu_mem_ctl.scala 424:54]
  wire  _T_1525 = ~fetch_req_icache_f; // @[el2_ifu_mem_ctl.scala 424:76]
  wire  _T_1526 = _T_1524 & _T_1525; // @[el2_ifu_mem_ctl.scala 424:74]
  wire  _T_1528 = _T_1526 & _T_317; // @[el2_ifu_mem_ctl.scala 424:96]
  wire  ic_crit_wd_rdy_new_in = _T_1523 | _T_1528; // @[el2_ifu_mem_ctl.scala 423:143]
  wire  ic_crit_wd_rdy = ic_crit_wd_rdy_new_in | ic_crit_wd_rdy_new_ff; // @[el2_ifu_mem_ctl.scala 624:43]
  wire  _T_1249 = ic_crit_wd_rdy | _T_2233; // @[el2_ifu_mem_ctl.scala 370:38]
  wire  _T_1251 = _T_1249 | _T_2249; // @[el2_ifu_mem_ctl.scala 370:64]
  wire  _T_1252 = ~_T_1251; // @[el2_ifu_mem_ctl.scala 370:21]
  wire  _T_1253 = ~fetch_req_iccm_f; // @[el2_ifu_mem_ctl.scala 370:98]
  wire  sel_ic_data = _T_1252 & _T_1253; // @[el2_ifu_mem_ctl.scala 370:96]
  wire  _T_2456 = io_ic_tag_perr & sel_ic_data; // @[el2_ifu_mem_ctl.scala 469:44]
  wire  _T_1622 = ifu_fetch_addr_int_f[1] & ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 436:31]
  reg [7:0] ic_miss_buff_data_error; // @[el2_ifu_mem_ctl.scala 408:60]
  wire  _T_1566 = _T_1413 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1567 = _T_1416 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1574 = _T_1566 | _T_1567; // @[Mux.scala 27:72]
  wire  _T_1568 = _T_1419 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1575 = _T_1574 | _T_1568; // @[Mux.scala 27:72]
  wire  _T_1569 = _T_1422 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1576 = _T_1575 | _T_1569; // @[Mux.scala 27:72]
  wire  _T_1570 = _T_1425 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1577 = _T_1576 | _T_1570; // @[Mux.scala 27:72]
  wire  _T_1571 = _T_1428 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1578 = _T_1577 | _T_1571; // @[Mux.scala 27:72]
  wire  _T_1572 = _T_1431 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1579 = _T_1578 | _T_1572; // @[Mux.scala 27:72]
  wire  _T_1573 = _T_1434 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass = _T_1579 | _T_1573; // @[Mux.scala 27:72]
  wire  _T_1605 = _T_2166 & ic_miss_buff_data_error[0]; // @[Mux.scala 27:72]
  wire  _T_1606 = _T_2169 & ic_miss_buff_data_error[1]; // @[Mux.scala 27:72]
  wire  _T_1613 = _T_1605 | _T_1606; // @[Mux.scala 27:72]
  wire  _T_1607 = _T_2172 & ic_miss_buff_data_error[2]; // @[Mux.scala 27:72]
  wire  _T_1614 = _T_1613 | _T_1607; // @[Mux.scala 27:72]
  wire  _T_1608 = _T_2175 & ic_miss_buff_data_error[3]; // @[Mux.scala 27:72]
  wire  _T_1615 = _T_1614 | _T_1608; // @[Mux.scala 27:72]
  wire  _T_1609 = _T_2178 & ic_miss_buff_data_error[4]; // @[Mux.scala 27:72]
  wire  _T_1616 = _T_1615 | _T_1609; // @[Mux.scala 27:72]
  wire  _T_1610 = _T_2181 & ic_miss_buff_data_error[5]; // @[Mux.scala 27:72]
  wire  _T_1617 = _T_1616 | _T_1610; // @[Mux.scala 27:72]
  wire  _T_1611 = _T_2184 & ic_miss_buff_data_error[6]; // @[Mux.scala 27:72]
  wire  _T_1618 = _T_1617 | _T_1611; // @[Mux.scala 27:72]
  wire  _T_1612 = _T_2187 & ic_miss_buff_data_error[7]; // @[Mux.scala 27:72]
  wire  ic_miss_buff_data_error_bypass_inc = _T_1618 | _T_1612; // @[Mux.scala 27:72]
  wire  _T_1623 = ic_miss_buff_data_error_bypass | ic_miss_buff_data_error_bypass_inc; // @[el2_ifu_mem_ctl.scala 438:70]
  wire  ifu_byp_data_err_new = _T_1622 ? ic_miss_buff_data_error_bypass : _T_1623; // @[el2_ifu_mem_ctl.scala 436:56]
  wire  ifc_bus_acc_fault_f = ic_byp_hit_f & ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 381:42]
  wire  _T_2457 = ifc_region_acc_fault_final_f | ifc_bus_acc_fault_f; // @[el2_ifu_mem_ctl.scala 469:91]
  wire  _T_2458 = ~_T_2457; // @[el2_ifu_mem_ctl.scala 469:60]
  wire  ic_rd_parity_final_err = _T_2456 & _T_2458; // @[el2_ifu_mem_ctl.scala 469:58]
  reg  ic_debug_ict_array_sel_ff; // @[Reg.scala 27:20]
  reg  ic_tag_valid_out_1_0; // @[Reg.scala 27:20]
  wire  _T_10156 = _T_4949 & ic_tag_valid_out_1_0; // @[el2_ifu_mem_ctl.scala 761:10]
  reg  ic_tag_valid_out_1_1; // @[Reg.scala 27:20]
  wire  _T_10158 = _T_4950 & ic_tag_valid_out_1_1; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10411 = _T_10156 | _T_10158; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_2; // @[Reg.scala 27:20]
  wire  _T_10160 = _T_4951 & ic_tag_valid_out_1_2; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10412 = _T_10411 | _T_10160; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_3; // @[Reg.scala 27:20]
  wire  _T_10162 = _T_4952 & ic_tag_valid_out_1_3; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10413 = _T_10412 | _T_10162; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_4; // @[Reg.scala 27:20]
  wire  _T_10164 = _T_4953 & ic_tag_valid_out_1_4; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10414 = _T_10413 | _T_10164; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_5; // @[Reg.scala 27:20]
  wire  _T_10166 = _T_4954 & ic_tag_valid_out_1_5; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10415 = _T_10414 | _T_10166; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_6; // @[Reg.scala 27:20]
  wire  _T_10168 = _T_4955 & ic_tag_valid_out_1_6; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10416 = _T_10415 | _T_10168; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_7; // @[Reg.scala 27:20]
  wire  _T_10170 = _T_4956 & ic_tag_valid_out_1_7; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10417 = _T_10416 | _T_10170; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_8; // @[Reg.scala 27:20]
  wire  _T_10172 = _T_4957 & ic_tag_valid_out_1_8; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10418 = _T_10417 | _T_10172; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_9; // @[Reg.scala 27:20]
  wire  _T_10174 = _T_4958 & ic_tag_valid_out_1_9; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10419 = _T_10418 | _T_10174; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_10; // @[Reg.scala 27:20]
  wire  _T_10176 = _T_4959 & ic_tag_valid_out_1_10; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10420 = _T_10419 | _T_10176; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_11; // @[Reg.scala 27:20]
  wire  _T_10178 = _T_4960 & ic_tag_valid_out_1_11; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10421 = _T_10420 | _T_10178; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_12; // @[Reg.scala 27:20]
  wire  _T_10180 = _T_4961 & ic_tag_valid_out_1_12; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10422 = _T_10421 | _T_10180; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_13; // @[Reg.scala 27:20]
  wire  _T_10182 = _T_4962 & ic_tag_valid_out_1_13; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10423 = _T_10422 | _T_10182; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_14; // @[Reg.scala 27:20]
  wire  _T_10184 = _T_4963 & ic_tag_valid_out_1_14; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10424 = _T_10423 | _T_10184; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_15; // @[Reg.scala 27:20]
  wire  _T_10186 = _T_4964 & ic_tag_valid_out_1_15; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10425 = _T_10424 | _T_10186; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_16; // @[Reg.scala 27:20]
  wire  _T_10188 = _T_4965 & ic_tag_valid_out_1_16; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10426 = _T_10425 | _T_10188; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_17; // @[Reg.scala 27:20]
  wire  _T_10190 = _T_4966 & ic_tag_valid_out_1_17; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10427 = _T_10426 | _T_10190; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_18; // @[Reg.scala 27:20]
  wire  _T_10192 = _T_4967 & ic_tag_valid_out_1_18; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10428 = _T_10427 | _T_10192; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_19; // @[Reg.scala 27:20]
  wire  _T_10194 = _T_4968 & ic_tag_valid_out_1_19; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10429 = _T_10428 | _T_10194; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_20; // @[Reg.scala 27:20]
  wire  _T_10196 = _T_4969 & ic_tag_valid_out_1_20; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10430 = _T_10429 | _T_10196; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_21; // @[Reg.scala 27:20]
  wire  _T_10198 = _T_4970 & ic_tag_valid_out_1_21; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10431 = _T_10430 | _T_10198; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_22; // @[Reg.scala 27:20]
  wire  _T_10200 = _T_4971 & ic_tag_valid_out_1_22; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10432 = _T_10431 | _T_10200; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_23; // @[Reg.scala 27:20]
  wire  _T_10202 = _T_4972 & ic_tag_valid_out_1_23; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10433 = _T_10432 | _T_10202; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_24; // @[Reg.scala 27:20]
  wire  _T_10204 = _T_4973 & ic_tag_valid_out_1_24; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10434 = _T_10433 | _T_10204; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_25; // @[Reg.scala 27:20]
  wire  _T_10206 = _T_4974 & ic_tag_valid_out_1_25; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10435 = _T_10434 | _T_10206; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_26; // @[Reg.scala 27:20]
  wire  _T_10208 = _T_4975 & ic_tag_valid_out_1_26; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10436 = _T_10435 | _T_10208; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_27; // @[Reg.scala 27:20]
  wire  _T_10210 = _T_4976 & ic_tag_valid_out_1_27; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10437 = _T_10436 | _T_10210; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_28; // @[Reg.scala 27:20]
  wire  _T_10212 = _T_4977 & ic_tag_valid_out_1_28; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10438 = _T_10437 | _T_10212; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_29; // @[Reg.scala 27:20]
  wire  _T_10214 = _T_4978 & ic_tag_valid_out_1_29; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10439 = _T_10438 | _T_10214; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_30; // @[Reg.scala 27:20]
  wire  _T_10216 = _T_4979 & ic_tag_valid_out_1_30; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10440 = _T_10439 | _T_10216; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_31; // @[Reg.scala 27:20]
  wire  _T_10218 = _T_4980 & ic_tag_valid_out_1_31; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10441 = _T_10440 | _T_10218; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_32; // @[Reg.scala 27:20]
  wire  _T_10220 = _T_4981 & ic_tag_valid_out_1_32; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10442 = _T_10441 | _T_10220; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_33; // @[Reg.scala 27:20]
  wire  _T_10222 = _T_4982 & ic_tag_valid_out_1_33; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10443 = _T_10442 | _T_10222; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_34; // @[Reg.scala 27:20]
  wire  _T_10224 = _T_4983 & ic_tag_valid_out_1_34; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10444 = _T_10443 | _T_10224; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_35; // @[Reg.scala 27:20]
  wire  _T_10226 = _T_4984 & ic_tag_valid_out_1_35; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10445 = _T_10444 | _T_10226; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_36; // @[Reg.scala 27:20]
  wire  _T_10228 = _T_4985 & ic_tag_valid_out_1_36; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10446 = _T_10445 | _T_10228; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_37; // @[Reg.scala 27:20]
  wire  _T_10230 = _T_4986 & ic_tag_valid_out_1_37; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10447 = _T_10446 | _T_10230; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_38; // @[Reg.scala 27:20]
  wire  _T_10232 = _T_4987 & ic_tag_valid_out_1_38; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10448 = _T_10447 | _T_10232; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_39; // @[Reg.scala 27:20]
  wire  _T_10234 = _T_4988 & ic_tag_valid_out_1_39; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10449 = _T_10448 | _T_10234; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_40; // @[Reg.scala 27:20]
  wire  _T_10236 = _T_4989 & ic_tag_valid_out_1_40; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10450 = _T_10449 | _T_10236; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_41; // @[Reg.scala 27:20]
  wire  _T_10238 = _T_4990 & ic_tag_valid_out_1_41; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10451 = _T_10450 | _T_10238; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_42; // @[Reg.scala 27:20]
  wire  _T_10240 = _T_4991 & ic_tag_valid_out_1_42; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10452 = _T_10451 | _T_10240; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_43; // @[Reg.scala 27:20]
  wire  _T_10242 = _T_4992 & ic_tag_valid_out_1_43; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10453 = _T_10452 | _T_10242; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_44; // @[Reg.scala 27:20]
  wire  _T_10244 = _T_4993 & ic_tag_valid_out_1_44; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10454 = _T_10453 | _T_10244; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_45; // @[Reg.scala 27:20]
  wire  _T_10246 = _T_4994 & ic_tag_valid_out_1_45; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10455 = _T_10454 | _T_10246; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_46; // @[Reg.scala 27:20]
  wire  _T_10248 = _T_4995 & ic_tag_valid_out_1_46; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10456 = _T_10455 | _T_10248; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_47; // @[Reg.scala 27:20]
  wire  _T_10250 = _T_4996 & ic_tag_valid_out_1_47; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10457 = _T_10456 | _T_10250; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_48; // @[Reg.scala 27:20]
  wire  _T_10252 = _T_4997 & ic_tag_valid_out_1_48; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10458 = _T_10457 | _T_10252; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_49; // @[Reg.scala 27:20]
  wire  _T_10254 = _T_4998 & ic_tag_valid_out_1_49; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10459 = _T_10458 | _T_10254; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_50; // @[Reg.scala 27:20]
  wire  _T_10256 = _T_4999 & ic_tag_valid_out_1_50; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10460 = _T_10459 | _T_10256; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_51; // @[Reg.scala 27:20]
  wire  _T_10258 = _T_5000 & ic_tag_valid_out_1_51; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10461 = _T_10460 | _T_10258; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_52; // @[Reg.scala 27:20]
  wire  _T_10260 = _T_5001 & ic_tag_valid_out_1_52; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10462 = _T_10461 | _T_10260; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_53; // @[Reg.scala 27:20]
  wire  _T_10262 = _T_5002 & ic_tag_valid_out_1_53; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10463 = _T_10462 | _T_10262; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_54; // @[Reg.scala 27:20]
  wire  _T_10264 = _T_5003 & ic_tag_valid_out_1_54; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10464 = _T_10463 | _T_10264; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_55; // @[Reg.scala 27:20]
  wire  _T_10266 = _T_5004 & ic_tag_valid_out_1_55; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10465 = _T_10464 | _T_10266; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_56; // @[Reg.scala 27:20]
  wire  _T_10268 = _T_5005 & ic_tag_valid_out_1_56; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10466 = _T_10465 | _T_10268; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_57; // @[Reg.scala 27:20]
  wire  _T_10270 = _T_5006 & ic_tag_valid_out_1_57; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10467 = _T_10466 | _T_10270; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_58; // @[Reg.scala 27:20]
  wire  _T_10272 = _T_5007 & ic_tag_valid_out_1_58; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10468 = _T_10467 | _T_10272; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_59; // @[Reg.scala 27:20]
  wire  _T_10274 = _T_5008 & ic_tag_valid_out_1_59; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10469 = _T_10468 | _T_10274; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_60; // @[Reg.scala 27:20]
  wire  _T_10276 = _T_5009 & ic_tag_valid_out_1_60; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10470 = _T_10469 | _T_10276; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_61; // @[Reg.scala 27:20]
  wire  _T_10278 = _T_5010 & ic_tag_valid_out_1_61; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10471 = _T_10470 | _T_10278; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_62; // @[Reg.scala 27:20]
  wire  _T_10280 = _T_5011 & ic_tag_valid_out_1_62; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10472 = _T_10471 | _T_10280; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_63; // @[Reg.scala 27:20]
  wire  _T_10282 = _T_5012 & ic_tag_valid_out_1_63; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10473 = _T_10472 | _T_10282; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_64; // @[Reg.scala 27:20]
  wire  _T_10284 = _T_5013 & ic_tag_valid_out_1_64; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10474 = _T_10473 | _T_10284; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_65; // @[Reg.scala 27:20]
  wire  _T_10286 = _T_5014 & ic_tag_valid_out_1_65; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10475 = _T_10474 | _T_10286; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_66; // @[Reg.scala 27:20]
  wire  _T_10288 = _T_5015 & ic_tag_valid_out_1_66; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10476 = _T_10475 | _T_10288; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_67; // @[Reg.scala 27:20]
  wire  _T_10290 = _T_5016 & ic_tag_valid_out_1_67; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10477 = _T_10476 | _T_10290; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_68; // @[Reg.scala 27:20]
  wire  _T_10292 = _T_5017 & ic_tag_valid_out_1_68; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10478 = _T_10477 | _T_10292; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_69; // @[Reg.scala 27:20]
  wire  _T_10294 = _T_5018 & ic_tag_valid_out_1_69; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10479 = _T_10478 | _T_10294; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_70; // @[Reg.scala 27:20]
  wire  _T_10296 = _T_5019 & ic_tag_valid_out_1_70; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10480 = _T_10479 | _T_10296; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_71; // @[Reg.scala 27:20]
  wire  _T_10298 = _T_5020 & ic_tag_valid_out_1_71; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10481 = _T_10480 | _T_10298; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_72; // @[Reg.scala 27:20]
  wire  _T_10300 = _T_5021 & ic_tag_valid_out_1_72; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10482 = _T_10481 | _T_10300; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_73; // @[Reg.scala 27:20]
  wire  _T_10302 = _T_5022 & ic_tag_valid_out_1_73; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10483 = _T_10482 | _T_10302; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_74; // @[Reg.scala 27:20]
  wire  _T_10304 = _T_5023 & ic_tag_valid_out_1_74; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10484 = _T_10483 | _T_10304; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_75; // @[Reg.scala 27:20]
  wire  _T_10306 = _T_5024 & ic_tag_valid_out_1_75; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10485 = _T_10484 | _T_10306; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_76; // @[Reg.scala 27:20]
  wire  _T_10308 = _T_5025 & ic_tag_valid_out_1_76; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10486 = _T_10485 | _T_10308; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_77; // @[Reg.scala 27:20]
  wire  _T_10310 = _T_5026 & ic_tag_valid_out_1_77; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10487 = _T_10486 | _T_10310; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_78; // @[Reg.scala 27:20]
  wire  _T_10312 = _T_5027 & ic_tag_valid_out_1_78; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10488 = _T_10487 | _T_10312; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_79; // @[Reg.scala 27:20]
  wire  _T_10314 = _T_5028 & ic_tag_valid_out_1_79; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10489 = _T_10488 | _T_10314; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_80; // @[Reg.scala 27:20]
  wire  _T_10316 = _T_5029 & ic_tag_valid_out_1_80; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10490 = _T_10489 | _T_10316; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_81; // @[Reg.scala 27:20]
  wire  _T_10318 = _T_5030 & ic_tag_valid_out_1_81; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10491 = _T_10490 | _T_10318; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_82; // @[Reg.scala 27:20]
  wire  _T_10320 = _T_5031 & ic_tag_valid_out_1_82; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10492 = _T_10491 | _T_10320; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_83; // @[Reg.scala 27:20]
  wire  _T_10322 = _T_5032 & ic_tag_valid_out_1_83; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10493 = _T_10492 | _T_10322; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_84; // @[Reg.scala 27:20]
  wire  _T_10324 = _T_5033 & ic_tag_valid_out_1_84; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10494 = _T_10493 | _T_10324; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_85; // @[Reg.scala 27:20]
  wire  _T_10326 = _T_5034 & ic_tag_valid_out_1_85; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10495 = _T_10494 | _T_10326; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_86; // @[Reg.scala 27:20]
  wire  _T_10328 = _T_5035 & ic_tag_valid_out_1_86; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10496 = _T_10495 | _T_10328; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_87; // @[Reg.scala 27:20]
  wire  _T_10330 = _T_5036 & ic_tag_valid_out_1_87; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10497 = _T_10496 | _T_10330; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_88; // @[Reg.scala 27:20]
  wire  _T_10332 = _T_5037 & ic_tag_valid_out_1_88; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10498 = _T_10497 | _T_10332; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_89; // @[Reg.scala 27:20]
  wire  _T_10334 = _T_5038 & ic_tag_valid_out_1_89; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10499 = _T_10498 | _T_10334; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_90; // @[Reg.scala 27:20]
  wire  _T_10336 = _T_5039 & ic_tag_valid_out_1_90; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10500 = _T_10499 | _T_10336; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_91; // @[Reg.scala 27:20]
  wire  _T_10338 = _T_5040 & ic_tag_valid_out_1_91; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10501 = _T_10500 | _T_10338; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_92; // @[Reg.scala 27:20]
  wire  _T_10340 = _T_5041 & ic_tag_valid_out_1_92; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10502 = _T_10501 | _T_10340; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_93; // @[Reg.scala 27:20]
  wire  _T_10342 = _T_5042 & ic_tag_valid_out_1_93; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10503 = _T_10502 | _T_10342; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_94; // @[Reg.scala 27:20]
  wire  _T_10344 = _T_5043 & ic_tag_valid_out_1_94; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10504 = _T_10503 | _T_10344; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_95; // @[Reg.scala 27:20]
  wire  _T_10346 = _T_5044 & ic_tag_valid_out_1_95; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10505 = _T_10504 | _T_10346; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_96; // @[Reg.scala 27:20]
  wire  _T_10348 = _T_5045 & ic_tag_valid_out_1_96; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10506 = _T_10505 | _T_10348; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_97; // @[Reg.scala 27:20]
  wire  _T_10350 = _T_5046 & ic_tag_valid_out_1_97; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10507 = _T_10506 | _T_10350; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_98; // @[Reg.scala 27:20]
  wire  _T_10352 = _T_5047 & ic_tag_valid_out_1_98; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10508 = _T_10507 | _T_10352; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_99; // @[Reg.scala 27:20]
  wire  _T_10354 = _T_5048 & ic_tag_valid_out_1_99; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10509 = _T_10508 | _T_10354; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_100; // @[Reg.scala 27:20]
  wire  _T_10356 = _T_5049 & ic_tag_valid_out_1_100; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10510 = _T_10509 | _T_10356; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_101; // @[Reg.scala 27:20]
  wire  _T_10358 = _T_5050 & ic_tag_valid_out_1_101; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10511 = _T_10510 | _T_10358; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_102; // @[Reg.scala 27:20]
  wire  _T_10360 = _T_5051 & ic_tag_valid_out_1_102; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10512 = _T_10511 | _T_10360; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_103; // @[Reg.scala 27:20]
  wire  _T_10362 = _T_5052 & ic_tag_valid_out_1_103; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10513 = _T_10512 | _T_10362; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_104; // @[Reg.scala 27:20]
  wire  _T_10364 = _T_5053 & ic_tag_valid_out_1_104; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10514 = _T_10513 | _T_10364; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_105; // @[Reg.scala 27:20]
  wire  _T_10366 = _T_5054 & ic_tag_valid_out_1_105; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10515 = _T_10514 | _T_10366; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_106; // @[Reg.scala 27:20]
  wire  _T_10368 = _T_5055 & ic_tag_valid_out_1_106; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10516 = _T_10515 | _T_10368; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_107; // @[Reg.scala 27:20]
  wire  _T_10370 = _T_5056 & ic_tag_valid_out_1_107; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10517 = _T_10516 | _T_10370; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_108; // @[Reg.scala 27:20]
  wire  _T_10372 = _T_5057 & ic_tag_valid_out_1_108; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10518 = _T_10517 | _T_10372; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_109; // @[Reg.scala 27:20]
  wire  _T_10374 = _T_5058 & ic_tag_valid_out_1_109; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10519 = _T_10518 | _T_10374; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_110; // @[Reg.scala 27:20]
  wire  _T_10376 = _T_5059 & ic_tag_valid_out_1_110; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10520 = _T_10519 | _T_10376; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_111; // @[Reg.scala 27:20]
  wire  _T_10378 = _T_5060 & ic_tag_valid_out_1_111; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10521 = _T_10520 | _T_10378; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_112; // @[Reg.scala 27:20]
  wire  _T_10380 = _T_5061 & ic_tag_valid_out_1_112; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10522 = _T_10521 | _T_10380; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_113; // @[Reg.scala 27:20]
  wire  _T_10382 = _T_5062 & ic_tag_valid_out_1_113; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10523 = _T_10522 | _T_10382; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_114; // @[Reg.scala 27:20]
  wire  _T_10384 = _T_5063 & ic_tag_valid_out_1_114; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10524 = _T_10523 | _T_10384; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_115; // @[Reg.scala 27:20]
  wire  _T_10386 = _T_5064 & ic_tag_valid_out_1_115; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10525 = _T_10524 | _T_10386; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_116; // @[Reg.scala 27:20]
  wire  _T_10388 = _T_5065 & ic_tag_valid_out_1_116; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10526 = _T_10525 | _T_10388; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_117; // @[Reg.scala 27:20]
  wire  _T_10390 = _T_5066 & ic_tag_valid_out_1_117; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10527 = _T_10526 | _T_10390; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_118; // @[Reg.scala 27:20]
  wire  _T_10392 = _T_5067 & ic_tag_valid_out_1_118; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10528 = _T_10527 | _T_10392; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_119; // @[Reg.scala 27:20]
  wire  _T_10394 = _T_5068 & ic_tag_valid_out_1_119; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10529 = _T_10528 | _T_10394; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_120; // @[Reg.scala 27:20]
  wire  _T_10396 = _T_5069 & ic_tag_valid_out_1_120; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10530 = _T_10529 | _T_10396; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_121; // @[Reg.scala 27:20]
  wire  _T_10398 = _T_5070 & ic_tag_valid_out_1_121; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10531 = _T_10530 | _T_10398; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_122; // @[Reg.scala 27:20]
  wire  _T_10400 = _T_5071 & ic_tag_valid_out_1_122; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10532 = _T_10531 | _T_10400; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_123; // @[Reg.scala 27:20]
  wire  _T_10402 = _T_5072 & ic_tag_valid_out_1_123; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10533 = _T_10532 | _T_10402; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_124; // @[Reg.scala 27:20]
  wire  _T_10404 = _T_5073 & ic_tag_valid_out_1_124; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10534 = _T_10533 | _T_10404; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_125; // @[Reg.scala 27:20]
  wire  _T_10406 = _T_5074 & ic_tag_valid_out_1_125; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10535 = _T_10534 | _T_10406; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_126; // @[Reg.scala 27:20]
  wire  _T_10408 = _T_5075 & ic_tag_valid_out_1_126; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10536 = _T_10535 | _T_10408; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_1_127; // @[Reg.scala 27:20]
  wire  _T_10410 = _T_5076 & ic_tag_valid_out_1_127; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10537 = _T_10536 | _T_10410; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_0; // @[Reg.scala 27:20]
  wire  _T_9773 = _T_4949 & ic_tag_valid_out_0_0; // @[el2_ifu_mem_ctl.scala 761:10]
  reg  ic_tag_valid_out_0_1; // @[Reg.scala 27:20]
  wire  _T_9775 = _T_4950 & ic_tag_valid_out_0_1; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10028 = _T_9773 | _T_9775; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_2; // @[Reg.scala 27:20]
  wire  _T_9777 = _T_4951 & ic_tag_valid_out_0_2; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10029 = _T_10028 | _T_9777; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_3; // @[Reg.scala 27:20]
  wire  _T_9779 = _T_4952 & ic_tag_valid_out_0_3; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10030 = _T_10029 | _T_9779; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_4; // @[Reg.scala 27:20]
  wire  _T_9781 = _T_4953 & ic_tag_valid_out_0_4; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10031 = _T_10030 | _T_9781; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_5; // @[Reg.scala 27:20]
  wire  _T_9783 = _T_4954 & ic_tag_valid_out_0_5; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10032 = _T_10031 | _T_9783; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_6; // @[Reg.scala 27:20]
  wire  _T_9785 = _T_4955 & ic_tag_valid_out_0_6; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10033 = _T_10032 | _T_9785; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_7; // @[Reg.scala 27:20]
  wire  _T_9787 = _T_4956 & ic_tag_valid_out_0_7; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10034 = _T_10033 | _T_9787; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_8; // @[Reg.scala 27:20]
  wire  _T_9789 = _T_4957 & ic_tag_valid_out_0_8; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10035 = _T_10034 | _T_9789; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_9; // @[Reg.scala 27:20]
  wire  _T_9791 = _T_4958 & ic_tag_valid_out_0_9; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10036 = _T_10035 | _T_9791; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_10; // @[Reg.scala 27:20]
  wire  _T_9793 = _T_4959 & ic_tag_valid_out_0_10; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10037 = _T_10036 | _T_9793; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_11; // @[Reg.scala 27:20]
  wire  _T_9795 = _T_4960 & ic_tag_valid_out_0_11; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10038 = _T_10037 | _T_9795; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_12; // @[Reg.scala 27:20]
  wire  _T_9797 = _T_4961 & ic_tag_valid_out_0_12; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10039 = _T_10038 | _T_9797; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_13; // @[Reg.scala 27:20]
  wire  _T_9799 = _T_4962 & ic_tag_valid_out_0_13; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10040 = _T_10039 | _T_9799; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_14; // @[Reg.scala 27:20]
  wire  _T_9801 = _T_4963 & ic_tag_valid_out_0_14; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10041 = _T_10040 | _T_9801; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_15; // @[Reg.scala 27:20]
  wire  _T_9803 = _T_4964 & ic_tag_valid_out_0_15; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10042 = _T_10041 | _T_9803; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_16; // @[Reg.scala 27:20]
  wire  _T_9805 = _T_4965 & ic_tag_valid_out_0_16; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10043 = _T_10042 | _T_9805; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_17; // @[Reg.scala 27:20]
  wire  _T_9807 = _T_4966 & ic_tag_valid_out_0_17; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10044 = _T_10043 | _T_9807; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_18; // @[Reg.scala 27:20]
  wire  _T_9809 = _T_4967 & ic_tag_valid_out_0_18; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10045 = _T_10044 | _T_9809; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_19; // @[Reg.scala 27:20]
  wire  _T_9811 = _T_4968 & ic_tag_valid_out_0_19; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10046 = _T_10045 | _T_9811; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_20; // @[Reg.scala 27:20]
  wire  _T_9813 = _T_4969 & ic_tag_valid_out_0_20; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10047 = _T_10046 | _T_9813; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_21; // @[Reg.scala 27:20]
  wire  _T_9815 = _T_4970 & ic_tag_valid_out_0_21; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10048 = _T_10047 | _T_9815; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_22; // @[Reg.scala 27:20]
  wire  _T_9817 = _T_4971 & ic_tag_valid_out_0_22; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10049 = _T_10048 | _T_9817; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_23; // @[Reg.scala 27:20]
  wire  _T_9819 = _T_4972 & ic_tag_valid_out_0_23; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10050 = _T_10049 | _T_9819; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_24; // @[Reg.scala 27:20]
  wire  _T_9821 = _T_4973 & ic_tag_valid_out_0_24; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10051 = _T_10050 | _T_9821; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_25; // @[Reg.scala 27:20]
  wire  _T_9823 = _T_4974 & ic_tag_valid_out_0_25; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10052 = _T_10051 | _T_9823; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_26; // @[Reg.scala 27:20]
  wire  _T_9825 = _T_4975 & ic_tag_valid_out_0_26; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10053 = _T_10052 | _T_9825; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_27; // @[Reg.scala 27:20]
  wire  _T_9827 = _T_4976 & ic_tag_valid_out_0_27; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10054 = _T_10053 | _T_9827; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_28; // @[Reg.scala 27:20]
  wire  _T_9829 = _T_4977 & ic_tag_valid_out_0_28; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10055 = _T_10054 | _T_9829; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_29; // @[Reg.scala 27:20]
  wire  _T_9831 = _T_4978 & ic_tag_valid_out_0_29; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10056 = _T_10055 | _T_9831; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_30; // @[Reg.scala 27:20]
  wire  _T_9833 = _T_4979 & ic_tag_valid_out_0_30; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10057 = _T_10056 | _T_9833; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_31; // @[Reg.scala 27:20]
  wire  _T_9835 = _T_4980 & ic_tag_valid_out_0_31; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10058 = _T_10057 | _T_9835; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_32; // @[Reg.scala 27:20]
  wire  _T_9837 = _T_4981 & ic_tag_valid_out_0_32; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10059 = _T_10058 | _T_9837; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_33; // @[Reg.scala 27:20]
  wire  _T_9839 = _T_4982 & ic_tag_valid_out_0_33; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10060 = _T_10059 | _T_9839; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_34; // @[Reg.scala 27:20]
  wire  _T_9841 = _T_4983 & ic_tag_valid_out_0_34; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10061 = _T_10060 | _T_9841; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_35; // @[Reg.scala 27:20]
  wire  _T_9843 = _T_4984 & ic_tag_valid_out_0_35; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10062 = _T_10061 | _T_9843; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_36; // @[Reg.scala 27:20]
  wire  _T_9845 = _T_4985 & ic_tag_valid_out_0_36; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10063 = _T_10062 | _T_9845; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_37; // @[Reg.scala 27:20]
  wire  _T_9847 = _T_4986 & ic_tag_valid_out_0_37; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10064 = _T_10063 | _T_9847; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_38; // @[Reg.scala 27:20]
  wire  _T_9849 = _T_4987 & ic_tag_valid_out_0_38; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10065 = _T_10064 | _T_9849; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_39; // @[Reg.scala 27:20]
  wire  _T_9851 = _T_4988 & ic_tag_valid_out_0_39; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10066 = _T_10065 | _T_9851; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_40; // @[Reg.scala 27:20]
  wire  _T_9853 = _T_4989 & ic_tag_valid_out_0_40; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10067 = _T_10066 | _T_9853; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_41; // @[Reg.scala 27:20]
  wire  _T_9855 = _T_4990 & ic_tag_valid_out_0_41; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10068 = _T_10067 | _T_9855; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_42; // @[Reg.scala 27:20]
  wire  _T_9857 = _T_4991 & ic_tag_valid_out_0_42; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10069 = _T_10068 | _T_9857; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_43; // @[Reg.scala 27:20]
  wire  _T_9859 = _T_4992 & ic_tag_valid_out_0_43; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10070 = _T_10069 | _T_9859; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_44; // @[Reg.scala 27:20]
  wire  _T_9861 = _T_4993 & ic_tag_valid_out_0_44; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10071 = _T_10070 | _T_9861; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_45; // @[Reg.scala 27:20]
  wire  _T_9863 = _T_4994 & ic_tag_valid_out_0_45; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10072 = _T_10071 | _T_9863; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_46; // @[Reg.scala 27:20]
  wire  _T_9865 = _T_4995 & ic_tag_valid_out_0_46; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10073 = _T_10072 | _T_9865; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_47; // @[Reg.scala 27:20]
  wire  _T_9867 = _T_4996 & ic_tag_valid_out_0_47; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10074 = _T_10073 | _T_9867; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_48; // @[Reg.scala 27:20]
  wire  _T_9869 = _T_4997 & ic_tag_valid_out_0_48; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10075 = _T_10074 | _T_9869; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_49; // @[Reg.scala 27:20]
  wire  _T_9871 = _T_4998 & ic_tag_valid_out_0_49; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10076 = _T_10075 | _T_9871; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_50; // @[Reg.scala 27:20]
  wire  _T_9873 = _T_4999 & ic_tag_valid_out_0_50; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10077 = _T_10076 | _T_9873; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_51; // @[Reg.scala 27:20]
  wire  _T_9875 = _T_5000 & ic_tag_valid_out_0_51; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10078 = _T_10077 | _T_9875; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_52; // @[Reg.scala 27:20]
  wire  _T_9877 = _T_5001 & ic_tag_valid_out_0_52; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10079 = _T_10078 | _T_9877; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_53; // @[Reg.scala 27:20]
  wire  _T_9879 = _T_5002 & ic_tag_valid_out_0_53; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10080 = _T_10079 | _T_9879; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_54; // @[Reg.scala 27:20]
  wire  _T_9881 = _T_5003 & ic_tag_valid_out_0_54; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10081 = _T_10080 | _T_9881; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_55; // @[Reg.scala 27:20]
  wire  _T_9883 = _T_5004 & ic_tag_valid_out_0_55; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10082 = _T_10081 | _T_9883; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_56; // @[Reg.scala 27:20]
  wire  _T_9885 = _T_5005 & ic_tag_valid_out_0_56; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10083 = _T_10082 | _T_9885; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_57; // @[Reg.scala 27:20]
  wire  _T_9887 = _T_5006 & ic_tag_valid_out_0_57; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10084 = _T_10083 | _T_9887; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_58; // @[Reg.scala 27:20]
  wire  _T_9889 = _T_5007 & ic_tag_valid_out_0_58; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10085 = _T_10084 | _T_9889; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_59; // @[Reg.scala 27:20]
  wire  _T_9891 = _T_5008 & ic_tag_valid_out_0_59; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10086 = _T_10085 | _T_9891; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_60; // @[Reg.scala 27:20]
  wire  _T_9893 = _T_5009 & ic_tag_valid_out_0_60; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10087 = _T_10086 | _T_9893; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_61; // @[Reg.scala 27:20]
  wire  _T_9895 = _T_5010 & ic_tag_valid_out_0_61; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10088 = _T_10087 | _T_9895; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_62; // @[Reg.scala 27:20]
  wire  _T_9897 = _T_5011 & ic_tag_valid_out_0_62; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10089 = _T_10088 | _T_9897; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_63; // @[Reg.scala 27:20]
  wire  _T_9899 = _T_5012 & ic_tag_valid_out_0_63; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10090 = _T_10089 | _T_9899; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_64; // @[Reg.scala 27:20]
  wire  _T_9901 = _T_5013 & ic_tag_valid_out_0_64; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10091 = _T_10090 | _T_9901; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_65; // @[Reg.scala 27:20]
  wire  _T_9903 = _T_5014 & ic_tag_valid_out_0_65; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10092 = _T_10091 | _T_9903; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_66; // @[Reg.scala 27:20]
  wire  _T_9905 = _T_5015 & ic_tag_valid_out_0_66; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10093 = _T_10092 | _T_9905; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_67; // @[Reg.scala 27:20]
  wire  _T_9907 = _T_5016 & ic_tag_valid_out_0_67; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10094 = _T_10093 | _T_9907; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_68; // @[Reg.scala 27:20]
  wire  _T_9909 = _T_5017 & ic_tag_valid_out_0_68; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10095 = _T_10094 | _T_9909; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_69; // @[Reg.scala 27:20]
  wire  _T_9911 = _T_5018 & ic_tag_valid_out_0_69; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10096 = _T_10095 | _T_9911; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_70; // @[Reg.scala 27:20]
  wire  _T_9913 = _T_5019 & ic_tag_valid_out_0_70; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10097 = _T_10096 | _T_9913; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_71; // @[Reg.scala 27:20]
  wire  _T_9915 = _T_5020 & ic_tag_valid_out_0_71; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10098 = _T_10097 | _T_9915; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_72; // @[Reg.scala 27:20]
  wire  _T_9917 = _T_5021 & ic_tag_valid_out_0_72; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10099 = _T_10098 | _T_9917; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_73; // @[Reg.scala 27:20]
  wire  _T_9919 = _T_5022 & ic_tag_valid_out_0_73; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10100 = _T_10099 | _T_9919; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_74; // @[Reg.scala 27:20]
  wire  _T_9921 = _T_5023 & ic_tag_valid_out_0_74; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10101 = _T_10100 | _T_9921; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_75; // @[Reg.scala 27:20]
  wire  _T_9923 = _T_5024 & ic_tag_valid_out_0_75; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10102 = _T_10101 | _T_9923; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_76; // @[Reg.scala 27:20]
  wire  _T_9925 = _T_5025 & ic_tag_valid_out_0_76; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10103 = _T_10102 | _T_9925; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_77; // @[Reg.scala 27:20]
  wire  _T_9927 = _T_5026 & ic_tag_valid_out_0_77; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10104 = _T_10103 | _T_9927; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_78; // @[Reg.scala 27:20]
  wire  _T_9929 = _T_5027 & ic_tag_valid_out_0_78; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10105 = _T_10104 | _T_9929; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_79; // @[Reg.scala 27:20]
  wire  _T_9931 = _T_5028 & ic_tag_valid_out_0_79; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10106 = _T_10105 | _T_9931; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_80; // @[Reg.scala 27:20]
  wire  _T_9933 = _T_5029 & ic_tag_valid_out_0_80; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10107 = _T_10106 | _T_9933; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_81; // @[Reg.scala 27:20]
  wire  _T_9935 = _T_5030 & ic_tag_valid_out_0_81; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10108 = _T_10107 | _T_9935; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_82; // @[Reg.scala 27:20]
  wire  _T_9937 = _T_5031 & ic_tag_valid_out_0_82; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10109 = _T_10108 | _T_9937; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_83; // @[Reg.scala 27:20]
  wire  _T_9939 = _T_5032 & ic_tag_valid_out_0_83; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10110 = _T_10109 | _T_9939; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_84; // @[Reg.scala 27:20]
  wire  _T_9941 = _T_5033 & ic_tag_valid_out_0_84; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10111 = _T_10110 | _T_9941; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_85; // @[Reg.scala 27:20]
  wire  _T_9943 = _T_5034 & ic_tag_valid_out_0_85; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10112 = _T_10111 | _T_9943; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_86; // @[Reg.scala 27:20]
  wire  _T_9945 = _T_5035 & ic_tag_valid_out_0_86; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10113 = _T_10112 | _T_9945; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_87; // @[Reg.scala 27:20]
  wire  _T_9947 = _T_5036 & ic_tag_valid_out_0_87; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10114 = _T_10113 | _T_9947; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_88; // @[Reg.scala 27:20]
  wire  _T_9949 = _T_5037 & ic_tag_valid_out_0_88; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10115 = _T_10114 | _T_9949; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_89; // @[Reg.scala 27:20]
  wire  _T_9951 = _T_5038 & ic_tag_valid_out_0_89; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10116 = _T_10115 | _T_9951; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_90; // @[Reg.scala 27:20]
  wire  _T_9953 = _T_5039 & ic_tag_valid_out_0_90; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10117 = _T_10116 | _T_9953; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_91; // @[Reg.scala 27:20]
  wire  _T_9955 = _T_5040 & ic_tag_valid_out_0_91; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10118 = _T_10117 | _T_9955; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_92; // @[Reg.scala 27:20]
  wire  _T_9957 = _T_5041 & ic_tag_valid_out_0_92; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10119 = _T_10118 | _T_9957; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_93; // @[Reg.scala 27:20]
  wire  _T_9959 = _T_5042 & ic_tag_valid_out_0_93; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10120 = _T_10119 | _T_9959; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_94; // @[Reg.scala 27:20]
  wire  _T_9961 = _T_5043 & ic_tag_valid_out_0_94; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10121 = _T_10120 | _T_9961; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_95; // @[Reg.scala 27:20]
  wire  _T_9963 = _T_5044 & ic_tag_valid_out_0_95; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10122 = _T_10121 | _T_9963; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_96; // @[Reg.scala 27:20]
  wire  _T_9965 = _T_5045 & ic_tag_valid_out_0_96; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10123 = _T_10122 | _T_9965; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_97; // @[Reg.scala 27:20]
  wire  _T_9967 = _T_5046 & ic_tag_valid_out_0_97; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10124 = _T_10123 | _T_9967; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_98; // @[Reg.scala 27:20]
  wire  _T_9969 = _T_5047 & ic_tag_valid_out_0_98; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10125 = _T_10124 | _T_9969; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_99; // @[Reg.scala 27:20]
  wire  _T_9971 = _T_5048 & ic_tag_valid_out_0_99; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10126 = _T_10125 | _T_9971; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_100; // @[Reg.scala 27:20]
  wire  _T_9973 = _T_5049 & ic_tag_valid_out_0_100; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10127 = _T_10126 | _T_9973; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_101; // @[Reg.scala 27:20]
  wire  _T_9975 = _T_5050 & ic_tag_valid_out_0_101; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10128 = _T_10127 | _T_9975; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_102; // @[Reg.scala 27:20]
  wire  _T_9977 = _T_5051 & ic_tag_valid_out_0_102; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10129 = _T_10128 | _T_9977; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_103; // @[Reg.scala 27:20]
  wire  _T_9979 = _T_5052 & ic_tag_valid_out_0_103; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10130 = _T_10129 | _T_9979; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_104; // @[Reg.scala 27:20]
  wire  _T_9981 = _T_5053 & ic_tag_valid_out_0_104; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10131 = _T_10130 | _T_9981; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_105; // @[Reg.scala 27:20]
  wire  _T_9983 = _T_5054 & ic_tag_valid_out_0_105; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10132 = _T_10131 | _T_9983; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_106; // @[Reg.scala 27:20]
  wire  _T_9985 = _T_5055 & ic_tag_valid_out_0_106; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10133 = _T_10132 | _T_9985; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_107; // @[Reg.scala 27:20]
  wire  _T_9987 = _T_5056 & ic_tag_valid_out_0_107; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10134 = _T_10133 | _T_9987; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_108; // @[Reg.scala 27:20]
  wire  _T_9989 = _T_5057 & ic_tag_valid_out_0_108; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10135 = _T_10134 | _T_9989; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_109; // @[Reg.scala 27:20]
  wire  _T_9991 = _T_5058 & ic_tag_valid_out_0_109; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10136 = _T_10135 | _T_9991; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_110; // @[Reg.scala 27:20]
  wire  _T_9993 = _T_5059 & ic_tag_valid_out_0_110; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10137 = _T_10136 | _T_9993; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_111; // @[Reg.scala 27:20]
  wire  _T_9995 = _T_5060 & ic_tag_valid_out_0_111; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10138 = _T_10137 | _T_9995; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_112; // @[Reg.scala 27:20]
  wire  _T_9997 = _T_5061 & ic_tag_valid_out_0_112; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10139 = _T_10138 | _T_9997; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_113; // @[Reg.scala 27:20]
  wire  _T_9999 = _T_5062 & ic_tag_valid_out_0_113; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10140 = _T_10139 | _T_9999; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_114; // @[Reg.scala 27:20]
  wire  _T_10001 = _T_5063 & ic_tag_valid_out_0_114; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10141 = _T_10140 | _T_10001; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_115; // @[Reg.scala 27:20]
  wire  _T_10003 = _T_5064 & ic_tag_valid_out_0_115; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10142 = _T_10141 | _T_10003; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_116; // @[Reg.scala 27:20]
  wire  _T_10005 = _T_5065 & ic_tag_valid_out_0_116; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10143 = _T_10142 | _T_10005; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_117; // @[Reg.scala 27:20]
  wire  _T_10007 = _T_5066 & ic_tag_valid_out_0_117; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10144 = _T_10143 | _T_10007; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_118; // @[Reg.scala 27:20]
  wire  _T_10009 = _T_5067 & ic_tag_valid_out_0_118; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10145 = _T_10144 | _T_10009; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_119; // @[Reg.scala 27:20]
  wire  _T_10011 = _T_5068 & ic_tag_valid_out_0_119; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10146 = _T_10145 | _T_10011; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_120; // @[Reg.scala 27:20]
  wire  _T_10013 = _T_5069 & ic_tag_valid_out_0_120; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10147 = _T_10146 | _T_10013; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_121; // @[Reg.scala 27:20]
  wire  _T_10015 = _T_5070 & ic_tag_valid_out_0_121; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10148 = _T_10147 | _T_10015; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_122; // @[Reg.scala 27:20]
  wire  _T_10017 = _T_5071 & ic_tag_valid_out_0_122; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10149 = _T_10148 | _T_10017; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_123; // @[Reg.scala 27:20]
  wire  _T_10019 = _T_5072 & ic_tag_valid_out_0_123; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10150 = _T_10149 | _T_10019; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_124; // @[Reg.scala 27:20]
  wire  _T_10021 = _T_5073 & ic_tag_valid_out_0_124; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10151 = _T_10150 | _T_10021; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_125; // @[Reg.scala 27:20]
  wire  _T_10023 = _T_5074 & ic_tag_valid_out_0_125; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10152 = _T_10151 | _T_10023; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_126; // @[Reg.scala 27:20]
  wire  _T_10025 = _T_5075 & ic_tag_valid_out_0_126; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10153 = _T_10152 | _T_10025; // @[el2_ifu_mem_ctl.scala 761:91]
  reg  ic_tag_valid_out_0_127; // @[Reg.scala 27:20]
  wire  _T_10027 = _T_5076 & ic_tag_valid_out_0_127; // @[el2_ifu_mem_ctl.scala 761:10]
  wire  _T_10154 = _T_10153 | _T_10027; // @[el2_ifu_mem_ctl.scala 761:91]
  wire [1:0] ic_tag_valid_unq = {_T_10537,_T_10154}; // @[Cat.scala 29:58]
  reg [1:0] ic_debug_way_ff; // @[Reg.scala 27:20]
  reg  ic_debug_rd_en_ff; // @[el2_ifu_mem_ctl.scala 835:54]
  wire [1:0] _T_10577 = ic_debug_rd_en_ff ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] _T_10578 = ic_debug_way_ff & _T_10577; // @[el2_ifu_mem_ctl.scala 816:67]
  wire [1:0] _T_10579 = ic_tag_valid_unq & _T_10578; // @[el2_ifu_mem_ctl.scala 816:48]
  wire  ic_debug_tag_val_rd_out = |_T_10579; // @[el2_ifu_mem_ctl.scala 816:115]
  wire [65:0] _T_1208 = {2'h0,io_ictag_debug_rd_data[25:21],32'h0,io_ictag_debug_rd_data[20:0],1'h0,way_status,3'h0,ic_debug_tag_val_rd_out}; // @[Cat.scala 29:58]
  reg [70:0] _T_1209; // @[Reg.scala 27:20]
  wire  ifu_wr_cumulative_err = ifu_wr_cumulative_err_data & _T_2591; // @[el2_ifu_mem_ctl.scala 364:80]
  wire  _T_1247 = ~ifu_byp_data_err_new; // @[el2_ifu_mem_ctl.scala 369:98]
  wire  sel_byp_data = _T_1251 & _T_1247; // @[el2_ifu_mem_ctl.scala 369:96]
  wire [63:0] _T_1258 = fetch_req_iccm_f ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1259 = _T_1258 & io_iccm_rd_data; // @[el2_ifu_mem_ctl.scala 376:69]
  wire [63:0] _T_1261 = sel_byp_data ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire  _T_2113 = ~ifu_fetch_addr_int_f[0]; // @[el2_ifu_mem_ctl.scala 444:31]
  wire  _T_1626 = ~ifu_fetch_addr_int_f[1]; // @[el2_ifu_mem_ctl.scala 440:38]
  wire [3:0] byp_fetch_index_inc_0 = {byp_fetch_index_inc,1'h0}; // @[Cat.scala 29:58]
  wire  _T_1627 = byp_fetch_index_inc_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1675 = _T_1627 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1630 = byp_fetch_index_inc_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1676 = _T_1630 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1691 = _T_1675 | _T_1676; // @[Mux.scala 27:72]
  wire  _T_1633 = byp_fetch_index_inc_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1677 = _T_1633 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1692 = _T_1691 | _T_1677; // @[Mux.scala 27:72]
  wire  _T_1636 = byp_fetch_index_inc_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1678 = _T_1636 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1693 = _T_1692 | _T_1678; // @[Mux.scala 27:72]
  wire  _T_1639 = byp_fetch_index_inc_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1679 = _T_1639 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1694 = _T_1693 | _T_1679; // @[Mux.scala 27:72]
  wire  _T_1642 = byp_fetch_index_inc_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1680 = _T_1642 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1695 = _T_1694 | _T_1680; // @[Mux.scala 27:72]
  wire  _T_1645 = byp_fetch_index_inc_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1681 = _T_1645 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1696 = _T_1695 | _T_1681; // @[Mux.scala 27:72]
  wire  _T_1648 = byp_fetch_index_inc_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1682 = _T_1648 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1697 = _T_1696 | _T_1682; // @[Mux.scala 27:72]
  wire  _T_1651 = byp_fetch_index_inc_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1683 = _T_1651 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1698 = _T_1697 | _T_1683; // @[Mux.scala 27:72]
  wire  _T_1654 = byp_fetch_index_inc_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1684 = _T_1654 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1699 = _T_1698 | _T_1684; // @[Mux.scala 27:72]
  wire  _T_1657 = byp_fetch_index_inc_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1685 = _T_1657 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1700 = _T_1699 | _T_1685; // @[Mux.scala 27:72]
  wire  _T_1660 = byp_fetch_index_inc_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1686 = _T_1660 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1701 = _T_1700 | _T_1686; // @[Mux.scala 27:72]
  wire  _T_1663 = byp_fetch_index_inc_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1687 = _T_1663 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1702 = _T_1701 | _T_1687; // @[Mux.scala 27:72]
  wire  _T_1666 = byp_fetch_index_inc_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1688 = _T_1666 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1703 = _T_1702 | _T_1688; // @[Mux.scala 27:72]
  wire  _T_1669 = byp_fetch_index_inc_0 == 4'he; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1689 = _T_1669 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1704 = _T_1703 | _T_1689; // @[Mux.scala 27:72]
  wire  _T_1672 = byp_fetch_index_inc_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 441:73]
  wire [15:0] _T_1690 = _T_1672 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1705 = _T_1704 | _T_1690; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_1 = {ifu_fetch_addr_int_f[4:2],1'h1}; // @[Cat.scala 29:58]
  wire  _T_1707 = byp_fetch_index_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1755 = _T_1707 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1710 = byp_fetch_index_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1756 = _T_1710 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1771 = _T_1755 | _T_1756; // @[Mux.scala 27:72]
  wire  _T_1713 = byp_fetch_index_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1757 = _T_1713 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1772 = _T_1771 | _T_1757; // @[Mux.scala 27:72]
  wire  _T_1716 = byp_fetch_index_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1758 = _T_1716 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1773 = _T_1772 | _T_1758; // @[Mux.scala 27:72]
  wire  _T_1719 = byp_fetch_index_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1759 = _T_1719 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1774 = _T_1773 | _T_1759; // @[Mux.scala 27:72]
  wire  _T_1722 = byp_fetch_index_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1760 = _T_1722 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1775 = _T_1774 | _T_1760; // @[Mux.scala 27:72]
  wire  _T_1725 = byp_fetch_index_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1761 = _T_1725 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1776 = _T_1775 | _T_1761; // @[Mux.scala 27:72]
  wire  _T_1728 = byp_fetch_index_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1762 = _T_1728 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1777 = _T_1776 | _T_1762; // @[Mux.scala 27:72]
  wire  _T_1731 = byp_fetch_index_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1763 = _T_1731 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1778 = _T_1777 | _T_1763; // @[Mux.scala 27:72]
  wire  _T_1734 = byp_fetch_index_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1764 = _T_1734 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1779 = _T_1778 | _T_1764; // @[Mux.scala 27:72]
  wire  _T_1737 = byp_fetch_index_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1765 = _T_1737 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1780 = _T_1779 | _T_1765; // @[Mux.scala 27:72]
  wire  _T_1740 = byp_fetch_index_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1766 = _T_1740 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1781 = _T_1780 | _T_1766; // @[Mux.scala 27:72]
  wire  _T_1743 = byp_fetch_index_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1767 = _T_1743 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1782 = _T_1781 | _T_1767; // @[Mux.scala 27:72]
  wire  _T_1746 = byp_fetch_index_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1768 = _T_1746 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1783 = _T_1782 | _T_1768; // @[Mux.scala 27:72]
  wire  _T_1749 = byp_fetch_index_1 == 4'he; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1769 = _T_1749 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1784 = _T_1783 | _T_1769; // @[Mux.scala 27:72]
  wire  _T_1752 = byp_fetch_index_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 441:179]
  wire [31:0] _T_1770 = _T_1752 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1785 = _T_1784 | _T_1770; // @[Mux.scala 27:72]
  wire [3:0] byp_fetch_index_0 = {ifu_fetch_addr_int_f[4:2],1'h0}; // @[Cat.scala 29:58]
  wire  _T_1787 = byp_fetch_index_0 == 4'h0; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1835 = _T_1787 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire  _T_1790 = byp_fetch_index_0 == 4'h1; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1836 = _T_1790 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1851 = _T_1835 | _T_1836; // @[Mux.scala 27:72]
  wire  _T_1793 = byp_fetch_index_0 == 4'h2; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1837 = _T_1793 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1852 = _T_1851 | _T_1837; // @[Mux.scala 27:72]
  wire  _T_1796 = byp_fetch_index_0 == 4'h3; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1838 = _T_1796 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1853 = _T_1852 | _T_1838; // @[Mux.scala 27:72]
  wire  _T_1799 = byp_fetch_index_0 == 4'h4; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1839 = _T_1799 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1854 = _T_1853 | _T_1839; // @[Mux.scala 27:72]
  wire  _T_1802 = byp_fetch_index_0 == 4'h5; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1840 = _T_1802 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1855 = _T_1854 | _T_1840; // @[Mux.scala 27:72]
  wire  _T_1805 = byp_fetch_index_0 == 4'h6; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1841 = _T_1805 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1856 = _T_1855 | _T_1841; // @[Mux.scala 27:72]
  wire  _T_1808 = byp_fetch_index_0 == 4'h7; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1842 = _T_1808 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1857 = _T_1856 | _T_1842; // @[Mux.scala 27:72]
  wire  _T_1811 = byp_fetch_index_0 == 4'h8; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1843 = _T_1811 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1858 = _T_1857 | _T_1843; // @[Mux.scala 27:72]
  wire  _T_1814 = byp_fetch_index_0 == 4'h9; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1844 = _T_1814 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1859 = _T_1858 | _T_1844; // @[Mux.scala 27:72]
  wire  _T_1817 = byp_fetch_index_0 == 4'ha; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1845 = _T_1817 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1860 = _T_1859 | _T_1845; // @[Mux.scala 27:72]
  wire  _T_1820 = byp_fetch_index_0 == 4'hb; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1846 = _T_1820 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1861 = _T_1860 | _T_1846; // @[Mux.scala 27:72]
  wire  _T_1823 = byp_fetch_index_0 == 4'hc; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1847 = _T_1823 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1862 = _T_1861 | _T_1847; // @[Mux.scala 27:72]
  wire  _T_1826 = byp_fetch_index_0 == 4'hd; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1848 = _T_1826 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1863 = _T_1862 | _T_1848; // @[Mux.scala 27:72]
  wire  _T_1829 = byp_fetch_index_0 == 4'he; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1849 = _T_1829 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1864 = _T_1863 | _T_1849; // @[Mux.scala 27:72]
  wire  _T_1832 = byp_fetch_index_0 == 4'hf; // @[el2_ifu_mem_ctl.scala 441:285]
  wire [31:0] _T_1850 = _T_1832 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1865 = _T_1864 | _T_1850; // @[Mux.scala 27:72]
  wire [79:0] _T_1868 = {_T_1705,_T_1785,_T_1865}; // @[Cat.scala 29:58]
  wire [3:0] byp_fetch_index_inc_1 = {byp_fetch_index_inc,1'h1}; // @[Cat.scala 29:58]
  wire  _T_1869 = byp_fetch_index_inc_1 == 4'h0; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1917 = _T_1869 ? ic_miss_buff_data_0[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire  _T_1872 = byp_fetch_index_inc_1 == 4'h1; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1918 = _T_1872 ? ic_miss_buff_data_1[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1933 = _T_1917 | _T_1918; // @[Mux.scala 27:72]
  wire  _T_1875 = byp_fetch_index_inc_1 == 4'h2; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1919 = _T_1875 ? ic_miss_buff_data_2[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1934 = _T_1933 | _T_1919; // @[Mux.scala 27:72]
  wire  _T_1878 = byp_fetch_index_inc_1 == 4'h3; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1920 = _T_1878 ? ic_miss_buff_data_3[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1935 = _T_1934 | _T_1920; // @[Mux.scala 27:72]
  wire  _T_1881 = byp_fetch_index_inc_1 == 4'h4; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1921 = _T_1881 ? ic_miss_buff_data_4[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1936 = _T_1935 | _T_1921; // @[Mux.scala 27:72]
  wire  _T_1884 = byp_fetch_index_inc_1 == 4'h5; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1922 = _T_1884 ? ic_miss_buff_data_5[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1937 = _T_1936 | _T_1922; // @[Mux.scala 27:72]
  wire  _T_1887 = byp_fetch_index_inc_1 == 4'h6; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1923 = _T_1887 ? ic_miss_buff_data_6[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1938 = _T_1937 | _T_1923; // @[Mux.scala 27:72]
  wire  _T_1890 = byp_fetch_index_inc_1 == 4'h7; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1924 = _T_1890 ? ic_miss_buff_data_7[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1939 = _T_1938 | _T_1924; // @[Mux.scala 27:72]
  wire  _T_1893 = byp_fetch_index_inc_1 == 4'h8; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1925 = _T_1893 ? ic_miss_buff_data_8[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1940 = _T_1939 | _T_1925; // @[Mux.scala 27:72]
  wire  _T_1896 = byp_fetch_index_inc_1 == 4'h9; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1926 = _T_1896 ? ic_miss_buff_data_9[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1941 = _T_1940 | _T_1926; // @[Mux.scala 27:72]
  wire  _T_1899 = byp_fetch_index_inc_1 == 4'ha; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1927 = _T_1899 ? ic_miss_buff_data_10[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1942 = _T_1941 | _T_1927; // @[Mux.scala 27:72]
  wire  _T_1902 = byp_fetch_index_inc_1 == 4'hb; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1928 = _T_1902 ? ic_miss_buff_data_11[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1943 = _T_1942 | _T_1928; // @[Mux.scala 27:72]
  wire  _T_1905 = byp_fetch_index_inc_1 == 4'hc; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1929 = _T_1905 ? ic_miss_buff_data_12[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1944 = _T_1943 | _T_1929; // @[Mux.scala 27:72]
  wire  _T_1908 = byp_fetch_index_inc_1 == 4'hd; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1930 = _T_1908 ? ic_miss_buff_data_13[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1945 = _T_1944 | _T_1930; // @[Mux.scala 27:72]
  wire  _T_1911 = byp_fetch_index_inc_1 == 4'he; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1931 = _T_1911 ? ic_miss_buff_data_14[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1946 = _T_1945 | _T_1931; // @[Mux.scala 27:72]
  wire  _T_1914 = byp_fetch_index_inc_1 == 4'hf; // @[el2_ifu_mem_ctl.scala 442:73]
  wire [15:0] _T_1932 = _T_1914 ? ic_miss_buff_data_15[15:0] : 16'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_1947 = _T_1946 | _T_1932; // @[Mux.scala 27:72]
  wire [31:0] _T_1997 = _T_1627 ? ic_miss_buff_data_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_1998 = _T_1630 ? ic_miss_buff_data_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2013 = _T_1997 | _T_1998; // @[Mux.scala 27:72]
  wire [31:0] _T_1999 = _T_1633 ? ic_miss_buff_data_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2014 = _T_2013 | _T_1999; // @[Mux.scala 27:72]
  wire [31:0] _T_2000 = _T_1636 ? ic_miss_buff_data_3 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2015 = _T_2014 | _T_2000; // @[Mux.scala 27:72]
  wire [31:0] _T_2001 = _T_1639 ? ic_miss_buff_data_4 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2016 = _T_2015 | _T_2001; // @[Mux.scala 27:72]
  wire [31:0] _T_2002 = _T_1642 ? ic_miss_buff_data_5 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2017 = _T_2016 | _T_2002; // @[Mux.scala 27:72]
  wire [31:0] _T_2003 = _T_1645 ? ic_miss_buff_data_6 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2018 = _T_2017 | _T_2003; // @[Mux.scala 27:72]
  wire [31:0] _T_2004 = _T_1648 ? ic_miss_buff_data_7 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2019 = _T_2018 | _T_2004; // @[Mux.scala 27:72]
  wire [31:0] _T_2005 = _T_1651 ? ic_miss_buff_data_8 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2020 = _T_2019 | _T_2005; // @[Mux.scala 27:72]
  wire [31:0] _T_2006 = _T_1654 ? ic_miss_buff_data_9 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2021 = _T_2020 | _T_2006; // @[Mux.scala 27:72]
  wire [31:0] _T_2007 = _T_1657 ? ic_miss_buff_data_10 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2022 = _T_2021 | _T_2007; // @[Mux.scala 27:72]
  wire [31:0] _T_2008 = _T_1660 ? ic_miss_buff_data_11 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2023 = _T_2022 | _T_2008; // @[Mux.scala 27:72]
  wire [31:0] _T_2009 = _T_1663 ? ic_miss_buff_data_12 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2024 = _T_2023 | _T_2009; // @[Mux.scala 27:72]
  wire [31:0] _T_2010 = _T_1666 ? ic_miss_buff_data_13 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2025 = _T_2024 | _T_2010; // @[Mux.scala 27:72]
  wire [31:0] _T_2011 = _T_1669 ? ic_miss_buff_data_14 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2026 = _T_2025 | _T_2011; // @[Mux.scala 27:72]
  wire [31:0] _T_2012 = _T_1672 ? ic_miss_buff_data_15 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_2027 = _T_2026 | _T_2012; // @[Mux.scala 27:72]
  wire [79:0] _T_2110 = {_T_1947,_T_2027,_T_1785}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_pre_new = _T_1626 ? _T_1868 : _T_2110; // @[el2_ifu_mem_ctl.scala 440:37]
  wire [79:0] _T_2115 = {16'h0,ic_byp_data_only_pre_new[79:16]}; // @[Cat.scala 29:58]
  wire [79:0] ic_byp_data_only_new = _T_2113 ? ic_byp_data_only_pre_new : _T_2115; // @[el2_ifu_mem_ctl.scala 444:30]
  wire [79:0] _GEN_474 = {{16'd0}, _T_1261}; // @[el2_ifu_mem_ctl.scala 376:114]
  wire [79:0] _T_1262 = _GEN_474 & ic_byp_data_only_new; // @[el2_ifu_mem_ctl.scala 376:114]
  wire [79:0] _GEN_475 = {{16'd0}, _T_1259}; // @[el2_ifu_mem_ctl.scala 376:88]
  wire [79:0] ic_premux_data_temp = _GEN_475 | _T_1262; // @[el2_ifu_mem_ctl.scala 376:88]
  wire  fetch_req_f_qual = io_ic_hit_f & _T_317; // @[el2_ifu_mem_ctl.scala 383:38]
  wire [1:0] _T_1271 = ifc_region_acc_fault_f ? 2'h2 : 2'h0; // @[el2_ifu_mem_ctl.scala 387:8]
  wire  _T_1273 = fetch_req_f_qual & io_ifu_bp_inst_mask_f; // @[el2_ifu_mem_ctl.scala 389:45]
  wire  _T_1275 = byp_fetch_index == 5'h1f; // @[el2_ifu_mem_ctl.scala 389:80]
  wire  _T_1276 = ~_T_1275; // @[el2_ifu_mem_ctl.scala 389:71]
  wire  _T_1277 = _T_1273 & _T_1276; // @[el2_ifu_mem_ctl.scala 389:69]
  wire  _T_1278 = err_stop_state != 2'h2; // @[el2_ifu_mem_ctl.scala 389:131]
  wire  _T_1279 = _T_1277 & _T_1278; // @[el2_ifu_mem_ctl.scala 389:114]
  wire [7:0] _T_1368 = {ic_miss_buff_data_valid_in_7,ic_miss_buff_data_valid_in_6,ic_miss_buff_data_valid_in_5,ic_miss_buff_data_valid_in_4,ic_miss_buff_data_valid_in_3,ic_miss_buff_data_valid_in_2,ic_miss_buff_data_valid_in_1,ic_miss_buff_data_valid_in_0}; // @[Cat.scala 29:58]
  wire  _T_1373 = ic_miss_buff_data_error[0] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  _T_2659 = |io_ifu_axi_rresp; // @[el2_ifu_mem_ctl.scala 620:47]
  wire  _T_2660 = _T_2659 & _T_13; // @[el2_ifu_mem_ctl.scala 620:50]
  wire  bus_ifu_wr_data_error = _T_2660 & miss_pending; // @[el2_ifu_mem_ctl.scala 620:68]
  wire  ic_miss_buff_data_error_in_0 = write_fill_data_0 ? bus_ifu_wr_data_error : _T_1373; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1377 = ic_miss_buff_data_error[1] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_1 = write_fill_data_1 ? bus_ifu_wr_data_error : _T_1377; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1381 = ic_miss_buff_data_error[2] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_2 = write_fill_data_2 ? bus_ifu_wr_data_error : _T_1381; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1385 = ic_miss_buff_data_error[3] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_3 = write_fill_data_3 ? bus_ifu_wr_data_error : _T_1385; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1389 = ic_miss_buff_data_error[4] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_4 = write_fill_data_4 ? bus_ifu_wr_data_error : _T_1389; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1393 = ic_miss_buff_data_error[5] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_5 = write_fill_data_5 ? bus_ifu_wr_data_error : _T_1393; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1397 = ic_miss_buff_data_error[6] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_6 = write_fill_data_6 ? bus_ifu_wr_data_error : _T_1397; // @[el2_ifu_mem_ctl.scala 406:72]
  wire  _T_1401 = ic_miss_buff_data_error[7] & _T_1339; // @[el2_ifu_mem_ctl.scala 407:32]
  wire  ic_miss_buff_data_error_in_7 = write_fill_data_7 ? bus_ifu_wr_data_error : _T_1401; // @[el2_ifu_mem_ctl.scala 406:72]
  wire [7:0] _T_1408 = {ic_miss_buff_data_error_in_7,ic_miss_buff_data_error_in_6,ic_miss_buff_data_error_in_5,ic_miss_buff_data_error_in_4,ic_miss_buff_data_error_in_3,ic_miss_buff_data_error_in_2,ic_miss_buff_data_error_in_1,ic_miss_buff_data_error_in_0}; // @[Cat.scala 29:58]
  reg [6:0] perr_ic_index_ff; // @[Reg.scala 27:20]
  wire  _T_2465 = 3'h0 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2473 = _T_6 & _T_317; // @[el2_ifu_mem_ctl.scala 489:65]
  wire  _T_2474 = _T_2473 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 489:88]
  wire  _T_2476 = _T_2474 & _T_2587; // @[el2_ifu_mem_ctl.scala 489:112]
  wire  _T_2477 = 3'h1 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2478 = io_dec_tlu_flush_lower_wb | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 494:50]
  wire  _T_2480 = 3'h2 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2486 = 3'h4 == perr_state; // @[Conditional.scala 37:30]
  wire  _T_2488 = 3'h3 == perr_state; // @[Conditional.scala 37:30]
  wire  _GEN_39 = _T_2486 | _T_2488; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_2480 ? _T_2478 : _GEN_39; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_2477 ? _T_2478 : _GEN_41; // @[Conditional.scala 39:67]
  wire  perr_state_en = _T_2465 ? _T_2476 : _GEN_43; // @[Conditional.scala 40:58]
  wire  perr_sb_write_status = _T_2465 & perr_state_en; // @[Conditional.scala 40:58]
  wire  _T_2479 = io_dec_tlu_flush_lower_wb & io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 495:56]
  wire  _GEN_44 = _T_2477 & _T_2479; // @[Conditional.scala 39:67]
  wire  perr_sel_invalidate = _T_2465 ? 1'h0 : _GEN_44; // @[Conditional.scala 40:58]
  wire [1:0] perr_err_inv_way = perr_sel_invalidate ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 480:58]
  wire  _T_2462 = ~dma_sb_err_state_ff; // @[el2_ifu_mem_ctl.scala 479:49]
  wire  _T_2467 = io_ic_error_start & _T_317; // @[el2_ifu_mem_ctl.scala 488:87]
  wire  _T_2481 = io_dec_tlu_flush_err_wb & io_dec_tlu_flush_lower_wb; // @[el2_ifu_mem_ctl.scala 498:54]
  wire  _T_2482 = _T_2481 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 498:84]
  wire  _T_2491 = perr_state == 3'h2; // @[el2_ifu_mem_ctl.scala 519:66]
  wire  _T_2492 = io_dec_tlu_flush_err_wb & _T_2491; // @[el2_ifu_mem_ctl.scala 519:52]
  wire  _T_2494 = _T_2492 & _T_2587; // @[el2_ifu_mem_ctl.scala 519:81]
  wire  _T_2496 = io_dec_tlu_flush_lower_wb | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 522:59]
  wire  _T_2497 = _T_2496 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 522:86]
  wire  _T_2511 = _T_2496 | io_ifu_fetch_val[0]; // @[el2_ifu_mem_ctl.scala 525:81]
  wire  _T_2512 = _T_2511 | ifu_bp_hit_taken_q_f; // @[el2_ifu_mem_ctl.scala 525:103]
  wire  _T_2513 = _T_2512 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 525:126]
  wire  _T_2533 = _T_2511 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 532:103]
  wire  _T_2540 = ~io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 537:62]
  wire  _T_2541 = io_dec_tlu_flush_lower_wb & _T_2540; // @[el2_ifu_mem_ctl.scala 537:60]
  wire  _T_2542 = _T_2541 | io_dec_tlu_i0_commit_cmt; // @[el2_ifu_mem_ctl.scala 537:88]
  wire  _T_2543 = _T_2542 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 537:115]
  wire  _GEN_51 = _T_2539 & _T_2497; // @[Conditional.scala 39:67]
  wire  _GEN_54 = _T_2522 ? _T_2533 : _GEN_51; // @[Conditional.scala 39:67]
  wire  _GEN_56 = _T_2522 | _T_2539; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_2495 ? _T_2513 : _GEN_54; // @[Conditional.scala 39:67]
  wire  _GEN_60 = _T_2495 | _GEN_56; // @[Conditional.scala 39:67]
  wire  err_stop_state_en = _T_2490 ? _T_2494 : _GEN_58; // @[Conditional.scala 40:58]
  reg  ifu_bus_cmd_valid; // @[Reg.scala 27:20]
  wire  _T_2555 = ic_act_miss_f | ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 554:64]
  wire  _T_2557 = _T_2555 & _T_2587; // @[el2_ifu_mem_ctl.scala 554:85]
  reg [2:0] bus_cmd_beat_count; // @[Reg.scala 27:20]
  wire  _T_2559 = bus_cmd_beat_count == 3'h7; // @[el2_ifu_mem_ctl.scala 554:133]
  wire  _T_2560 = _T_2559 & ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 554:164]
  wire  _T_2561 = _T_2560 & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 554:184]
  wire  _T_2562 = _T_2561 & miss_pending; // @[el2_ifu_mem_ctl.scala 554:204]
  wire  _T_2563 = ~_T_2562; // @[el2_ifu_mem_ctl.scala 554:112]
  wire  ifc_bus_ic_req_ff_in = _T_2557 & _T_2563; // @[el2_ifu_mem_ctl.scala 554:110]
  wire  _T_2564 = io_ifu_bus_clk_en | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 555:80]
  wire  ifu_bus_arready = io_ifu_axi_arready & io_ifu_bus_clk_en; // @[el2_ifu_mem_ctl.scala 586:45]
  wire  _T_2581 = io_ifu_axi_arvalid & ifu_bus_arready; // @[el2_ifu_mem_ctl.scala 589:35]
  wire  _T_2582 = _T_2581 & miss_pending; // @[el2_ifu_mem_ctl.scala 589:53]
  wire  bus_cmd_sent = _T_2582 & _T_2587; // @[el2_ifu_mem_ctl.scala 589:68]
  wire [2:0] _T_2572 = ifu_bus_cmd_valid ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _T_2574 = {miss_addr,bus_rd_addr_count,3'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_2576 = ifu_bus_cmd_valid ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  reg  ifu_bus_arready_unq_ff; // @[Reg.scala 27:20]
  reg  ifu_bus_arvalid_ff; // @[Reg.scala 27:20]
  wire  ifu_bus_arready_ff = ifu_bus_arready_unq_ff & bus_ifu_bus_clk_en_ff; // @[el2_ifu_mem_ctl.scala 587:51]
  wire  _T_2602 = ~scnd_miss_req; // @[el2_ifu_mem_ctl.scala 597:73]
  wire  _T_2603 = _T_2588 & _T_2602; // @[el2_ifu_mem_ctl.scala 597:71]
  wire  _T_2605 = last_data_recieved_ff & _T_1339; // @[el2_ifu_mem_ctl.scala 597:114]
  wire  last_data_recieved_in = _T_2603 | _T_2605; // @[el2_ifu_mem_ctl.scala 597:89]
  wire [2:0] _T_2611 = bus_rd_addr_count + 3'h1; // @[el2_ifu_mem_ctl.scala 602:45]
  wire  _T_2614 = io_ifu_bus_clk_en | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 603:81]
  wire  _T_2615 = _T_2614 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 603:97]
  wire  _T_2617 = ifu_bus_cmd_valid & io_ifu_axi_arready; // @[el2_ifu_mem_ctl.scala 605:48]
  wire  _T_2618 = _T_2617 & miss_pending; // @[el2_ifu_mem_ctl.scala 605:68]
  wire  bus_inc_cmd_beat_cnt = _T_2618 & _T_2587; // @[el2_ifu_mem_ctl.scala 605:83]
  wire  bus_reset_cmd_beat_cnt_secondlast = ic_act_miss_f & uncacheable_miss_in; // @[el2_ifu_mem_ctl.scala 607:57]
  wire  _T_2622 = ~bus_inc_cmd_beat_cnt; // @[el2_ifu_mem_ctl.scala 608:31]
  wire  _T_2623 = ic_act_miss_f | scnd_miss_req; // @[el2_ifu_mem_ctl.scala 608:71]
  wire  _T_2624 = _T_2623 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 608:87]
  wire  _T_2625 = ~_T_2624; // @[el2_ifu_mem_ctl.scala 608:55]
  wire  bus_hold_cmd_beat_cnt = _T_2622 & _T_2625; // @[el2_ifu_mem_ctl.scala 608:53]
  wire  _T_2626 = bus_inc_cmd_beat_cnt | ic_act_miss_f; // @[el2_ifu_mem_ctl.scala 609:46]
  wire  bus_cmd_beat_en = _T_2626 | io_dec_tlu_force_halt; // @[el2_ifu_mem_ctl.scala 609:62]
  wire [2:0] _T_2629 = bus_cmd_beat_count + 3'h1; // @[el2_ifu_mem_ctl.scala 611:46]
  wire [2:0] _T_2631 = bus_reset_cmd_beat_cnt_secondlast ? 3'h6 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2632 = bus_inc_cmd_beat_cnt ? _T_2629 : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2633 = bus_hold_cmd_beat_cnt ? bus_cmd_beat_count : 3'h0; // @[Mux.scala 27:72]
  wire [2:0] _T_2635 = _T_2631 | _T_2632; // @[Mux.scala 27:72]
  wire [2:0] bus_new_cmd_beat_count = _T_2635 | _T_2633; // @[Mux.scala 27:72]
  wire  _T_2639 = _T_2615 & bus_cmd_beat_en; // @[el2_ifu_mem_ctl.scala 612:125]
  reg  ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 623:62]
  wire  _T_2667 = ~iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 628:50]
  wire  _T_2668 = io_ifc_dma_access_ok & _T_2667; // @[el2_ifu_mem_ctl.scala 628:47]
  wire  _T_2669 = ~io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 628:70]
  wire  ifc_dma_access_ok_d = _T_2668 & _T_2669; // @[el2_ifu_mem_ctl.scala 628:68]
  wire  _T_2673 = _T_2668 & ifc_dma_access_ok_prev; // @[el2_ifu_mem_ctl.scala 629:72]
  wire  _T_2674 = perr_state == 3'h0; // @[el2_ifu_mem_ctl.scala 629:111]
  wire  _T_2675 = _T_2673 & _T_2674; // @[el2_ifu_mem_ctl.scala 629:97]
  wire  ifc_dma_access_q_ok = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 629:127]
  wire  _T_2678 = ifc_dma_access_q_ok & io_dma_iccm_req; // @[el2_ifu_mem_ctl.scala 632:40]
  wire  _T_2679 = _T_2678 & io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 632:58]
  wire  _T_2682 = ~io_dma_mem_write; // @[el2_ifu_mem_ctl.scala 633:60]
  wire  _T_2683 = _T_2678 & _T_2682; // @[el2_ifu_mem_ctl.scala 633:58]
  wire  _T_2684 = io_ifc_iccm_access_bf & io_ifc_fetch_req_bf; // @[el2_ifu_mem_ctl.scala 633:104]
  wire [2:0] _T_2689 = io_dma_iccm_req ? 3'h7 : 3'h0; // @[Bitwise.scala 72:12]
  wire  _T_2710 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[1]; // @[el2_lib.scala 244:74]
  wire  _T_2711 = _T_2710 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 244:74]
  wire  _T_2712 = _T_2711 ^ io_dma_mem_wdata[4]; // @[el2_lib.scala 244:74]
  wire  _T_2713 = _T_2712 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 244:74]
  wire  _T_2714 = _T_2713 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 244:74]
  wire  _T_2715 = _T_2714 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2716 = _T_2715 ^ io_dma_mem_wdata[11]; // @[el2_lib.scala 244:74]
  wire  _T_2717 = _T_2716 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 244:74]
  wire  _T_2718 = _T_2717 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 244:74]
  wire  _T_2719 = _T_2718 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2720 = _T_2719 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 244:74]
  wire  _T_2721 = _T_2720 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2722 = _T_2721 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2723 = _T_2722 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2724 = _T_2723 ^ io_dma_mem_wdata[26]; // @[el2_lib.scala 244:74]
  wire  _T_2725 = _T_2724 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 244:74]
  wire  _T_2726 = _T_2725 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 244:74]
  wire  _T_2745 = io_dma_mem_wdata[0] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 244:74]
  wire  _T_2746 = _T_2745 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 244:74]
  wire  _T_2747 = _T_2746 ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 244:74]
  wire  _T_2748 = _T_2747 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 244:74]
  wire  _T_2749 = _T_2748 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 244:74]
  wire  _T_2750 = _T_2749 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2751 = _T_2750 ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 244:74]
  wire  _T_2752 = _T_2751 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 244:74]
  wire  _T_2753 = _T_2752 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 244:74]
  wire  _T_2754 = _T_2753 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2755 = _T_2754 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 244:74]
  wire  _T_2756 = _T_2755 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2757 = _T_2756 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2758 = _T_2757 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2759 = _T_2758 ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 244:74]
  wire  _T_2760 = _T_2759 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 244:74]
  wire  _T_2761 = _T_2760 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 244:74]
  wire  _T_2780 = io_dma_mem_wdata[1] ^ io_dma_mem_wdata[2]; // @[el2_lib.scala 244:74]
  wire  _T_2781 = _T_2780 ^ io_dma_mem_wdata[3]; // @[el2_lib.scala 244:74]
  wire  _T_2782 = _T_2781 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 244:74]
  wire  _T_2783 = _T_2782 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 244:74]
  wire  _T_2784 = _T_2783 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 244:74]
  wire  _T_2785 = _T_2784 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2786 = _T_2785 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 244:74]
  wire  _T_2787 = _T_2786 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 244:74]
  wire  _T_2788 = _T_2787 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 244:74]
  wire  _T_2789 = _T_2788 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2790 = _T_2789 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 244:74]
  wire  _T_2791 = _T_2790 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2792 = _T_2791 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2793 = _T_2792 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2794 = _T_2793 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 244:74]
  wire  _T_2795 = _T_2794 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 244:74]
  wire  _T_2796 = _T_2795 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 244:74]
  wire  _T_2812 = io_dma_mem_wdata[4] ^ io_dma_mem_wdata[5]; // @[el2_lib.scala 244:74]
  wire  _T_2813 = _T_2812 ^ io_dma_mem_wdata[6]; // @[el2_lib.scala 244:74]
  wire  _T_2814 = _T_2813 ^ io_dma_mem_wdata[7]; // @[el2_lib.scala 244:74]
  wire  _T_2815 = _T_2814 ^ io_dma_mem_wdata[8]; // @[el2_lib.scala 244:74]
  wire  _T_2816 = _T_2815 ^ io_dma_mem_wdata[9]; // @[el2_lib.scala 244:74]
  wire  _T_2817 = _T_2816 ^ io_dma_mem_wdata[10]; // @[el2_lib.scala 244:74]
  wire  _T_2818 = _T_2817 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 244:74]
  wire  _T_2819 = _T_2818 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 244:74]
  wire  _T_2820 = _T_2819 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 244:74]
  wire  _T_2821 = _T_2820 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2822 = _T_2821 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 244:74]
  wire  _T_2823 = _T_2822 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2824 = _T_2823 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2825 = _T_2824 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2841 = io_dma_mem_wdata[11] ^ io_dma_mem_wdata[12]; // @[el2_lib.scala 244:74]
  wire  _T_2842 = _T_2841 ^ io_dma_mem_wdata[13]; // @[el2_lib.scala 244:74]
  wire  _T_2843 = _T_2842 ^ io_dma_mem_wdata[14]; // @[el2_lib.scala 244:74]
  wire  _T_2844 = _T_2843 ^ io_dma_mem_wdata[15]; // @[el2_lib.scala 244:74]
  wire  _T_2845 = _T_2844 ^ io_dma_mem_wdata[16]; // @[el2_lib.scala 244:74]
  wire  _T_2846 = _T_2845 ^ io_dma_mem_wdata[17]; // @[el2_lib.scala 244:74]
  wire  _T_2847 = _T_2846 ^ io_dma_mem_wdata[18]; // @[el2_lib.scala 244:74]
  wire  _T_2848 = _T_2847 ^ io_dma_mem_wdata[19]; // @[el2_lib.scala 244:74]
  wire  _T_2849 = _T_2848 ^ io_dma_mem_wdata[20]; // @[el2_lib.scala 244:74]
  wire  _T_2850 = _T_2849 ^ io_dma_mem_wdata[21]; // @[el2_lib.scala 244:74]
  wire  _T_2851 = _T_2850 ^ io_dma_mem_wdata[22]; // @[el2_lib.scala 244:74]
  wire  _T_2852 = _T_2851 ^ io_dma_mem_wdata[23]; // @[el2_lib.scala 244:74]
  wire  _T_2853 = _T_2852 ^ io_dma_mem_wdata[24]; // @[el2_lib.scala 244:74]
  wire  _T_2854 = _T_2853 ^ io_dma_mem_wdata[25]; // @[el2_lib.scala 244:74]
  wire  _T_2861 = io_dma_mem_wdata[26] ^ io_dma_mem_wdata[27]; // @[el2_lib.scala 244:74]
  wire  _T_2862 = _T_2861 ^ io_dma_mem_wdata[28]; // @[el2_lib.scala 244:74]
  wire  _T_2863 = _T_2862 ^ io_dma_mem_wdata[29]; // @[el2_lib.scala 244:74]
  wire  _T_2864 = _T_2863 ^ io_dma_mem_wdata[30]; // @[el2_lib.scala 244:74]
  wire  _T_2865 = _T_2864 ^ io_dma_mem_wdata[31]; // @[el2_lib.scala 244:74]
  wire [5:0] _T_2870 = {_T_2865,_T_2854,_T_2825,_T_2796,_T_2761,_T_2726}; // @[Cat.scala 29:58]
  wire  _T_2871 = ^io_dma_mem_wdata[31:0]; // @[el2_lib.scala 252:13]
  wire  _T_2872 = ^_T_2870; // @[el2_lib.scala 252:23]
  wire  _T_2873 = _T_2871 ^ _T_2872; // @[el2_lib.scala 252:18]
  wire [6:0] _T_2874 = {_T_2873,_T_2865,_T_2854,_T_2825,_T_2796,_T_2761,_T_2726}; // @[Cat.scala 29:58]
  wire  _T_2894 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[33]; // @[el2_lib.scala 244:74]
  wire  _T_2895 = _T_2894 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 244:74]
  wire  _T_2896 = _T_2895 ^ io_dma_mem_wdata[36]; // @[el2_lib.scala 244:74]
  wire  _T_2897 = _T_2896 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 244:74]
  wire  _T_2898 = _T_2897 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 244:74]
  wire  _T_2899 = _T_2898 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_2900 = _T_2899 ^ io_dma_mem_wdata[43]; // @[el2_lib.scala 244:74]
  wire  _T_2901 = _T_2900 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 244:74]
  wire  _T_2902 = _T_2901 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 244:74]
  wire  _T_2903 = _T_2902 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_2904 = _T_2903 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 244:74]
  wire  _T_2905 = _T_2904 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_2906 = _T_2905 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_2907 = _T_2906 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_2908 = _T_2907 ^ io_dma_mem_wdata[58]; // @[el2_lib.scala 244:74]
  wire  _T_2909 = _T_2908 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 244:74]
  wire  _T_2910 = _T_2909 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 244:74]
  wire  _T_2929 = io_dma_mem_wdata[32] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 244:74]
  wire  _T_2930 = _T_2929 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 244:74]
  wire  _T_2931 = _T_2930 ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 244:74]
  wire  _T_2932 = _T_2931 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 244:74]
  wire  _T_2933 = _T_2932 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 244:74]
  wire  _T_2934 = _T_2933 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_2935 = _T_2934 ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 244:74]
  wire  _T_2936 = _T_2935 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 244:74]
  wire  _T_2937 = _T_2936 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 244:74]
  wire  _T_2938 = _T_2937 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_2939 = _T_2938 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 244:74]
  wire  _T_2940 = _T_2939 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_2941 = _T_2940 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_2942 = _T_2941 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_2943 = _T_2942 ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 244:74]
  wire  _T_2944 = _T_2943 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 244:74]
  wire  _T_2945 = _T_2944 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 244:74]
  wire  _T_2964 = io_dma_mem_wdata[33] ^ io_dma_mem_wdata[34]; // @[el2_lib.scala 244:74]
  wire  _T_2965 = _T_2964 ^ io_dma_mem_wdata[35]; // @[el2_lib.scala 244:74]
  wire  _T_2966 = _T_2965 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 244:74]
  wire  _T_2967 = _T_2966 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 244:74]
  wire  _T_2968 = _T_2967 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 244:74]
  wire  _T_2969 = _T_2968 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_2970 = _T_2969 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 244:74]
  wire  _T_2971 = _T_2970 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 244:74]
  wire  _T_2972 = _T_2971 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 244:74]
  wire  _T_2973 = _T_2972 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_2974 = _T_2973 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 244:74]
  wire  _T_2975 = _T_2974 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_2976 = _T_2975 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_2977 = _T_2976 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_2978 = _T_2977 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 244:74]
  wire  _T_2979 = _T_2978 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 244:74]
  wire  _T_2980 = _T_2979 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 244:74]
  wire  _T_2996 = io_dma_mem_wdata[36] ^ io_dma_mem_wdata[37]; // @[el2_lib.scala 244:74]
  wire  _T_2997 = _T_2996 ^ io_dma_mem_wdata[38]; // @[el2_lib.scala 244:74]
  wire  _T_2998 = _T_2997 ^ io_dma_mem_wdata[39]; // @[el2_lib.scala 244:74]
  wire  _T_2999 = _T_2998 ^ io_dma_mem_wdata[40]; // @[el2_lib.scala 244:74]
  wire  _T_3000 = _T_2999 ^ io_dma_mem_wdata[41]; // @[el2_lib.scala 244:74]
  wire  _T_3001 = _T_3000 ^ io_dma_mem_wdata[42]; // @[el2_lib.scala 244:74]
  wire  _T_3002 = _T_3001 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 244:74]
  wire  _T_3003 = _T_3002 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 244:74]
  wire  _T_3004 = _T_3003 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 244:74]
  wire  _T_3005 = _T_3004 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_3006 = _T_3005 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 244:74]
  wire  _T_3007 = _T_3006 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_3008 = _T_3007 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_3009 = _T_3008 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_3025 = io_dma_mem_wdata[43] ^ io_dma_mem_wdata[44]; // @[el2_lib.scala 244:74]
  wire  _T_3026 = _T_3025 ^ io_dma_mem_wdata[45]; // @[el2_lib.scala 244:74]
  wire  _T_3027 = _T_3026 ^ io_dma_mem_wdata[46]; // @[el2_lib.scala 244:74]
  wire  _T_3028 = _T_3027 ^ io_dma_mem_wdata[47]; // @[el2_lib.scala 244:74]
  wire  _T_3029 = _T_3028 ^ io_dma_mem_wdata[48]; // @[el2_lib.scala 244:74]
  wire  _T_3030 = _T_3029 ^ io_dma_mem_wdata[49]; // @[el2_lib.scala 244:74]
  wire  _T_3031 = _T_3030 ^ io_dma_mem_wdata[50]; // @[el2_lib.scala 244:74]
  wire  _T_3032 = _T_3031 ^ io_dma_mem_wdata[51]; // @[el2_lib.scala 244:74]
  wire  _T_3033 = _T_3032 ^ io_dma_mem_wdata[52]; // @[el2_lib.scala 244:74]
  wire  _T_3034 = _T_3033 ^ io_dma_mem_wdata[53]; // @[el2_lib.scala 244:74]
  wire  _T_3035 = _T_3034 ^ io_dma_mem_wdata[54]; // @[el2_lib.scala 244:74]
  wire  _T_3036 = _T_3035 ^ io_dma_mem_wdata[55]; // @[el2_lib.scala 244:74]
  wire  _T_3037 = _T_3036 ^ io_dma_mem_wdata[56]; // @[el2_lib.scala 244:74]
  wire  _T_3038 = _T_3037 ^ io_dma_mem_wdata[57]; // @[el2_lib.scala 244:74]
  wire  _T_3045 = io_dma_mem_wdata[58] ^ io_dma_mem_wdata[59]; // @[el2_lib.scala 244:74]
  wire  _T_3046 = _T_3045 ^ io_dma_mem_wdata[60]; // @[el2_lib.scala 244:74]
  wire  _T_3047 = _T_3046 ^ io_dma_mem_wdata[61]; // @[el2_lib.scala 244:74]
  wire  _T_3048 = _T_3047 ^ io_dma_mem_wdata[62]; // @[el2_lib.scala 244:74]
  wire  _T_3049 = _T_3048 ^ io_dma_mem_wdata[63]; // @[el2_lib.scala 244:74]
  wire [5:0] _T_3054 = {_T_3049,_T_3038,_T_3009,_T_2980,_T_2945,_T_2910}; // @[Cat.scala 29:58]
  wire  _T_3055 = ^io_dma_mem_wdata[63:32]; // @[el2_lib.scala 252:13]
  wire  _T_3056 = ^_T_3054; // @[el2_lib.scala 252:23]
  wire  _T_3057 = _T_3055 ^ _T_3056; // @[el2_lib.scala 252:18]
  wire [13:0] dma_mem_ecc = {_T_3057,_T_3049,_T_3038,_T_3009,_T_2980,_T_2945,_T_2910,_T_2874}; // @[Cat.scala 29:58]
  wire  _T_3244 = ~_T_2678; // @[el2_ifu_mem_ctl.scala 639:45]
  wire  _T_3245 = iccm_correct_ecc & _T_3244; // @[el2_ifu_mem_ctl.scala 639:43]
  reg [38:0] iccm_ecc_corr_data_ff; // @[Reg.scala 27:20]
  wire [77:0] _T_3246 = {iccm_ecc_corr_data_ff,iccm_ecc_corr_data_ff}; // @[Cat.scala 29:58]
  wire [77:0] _T_3253 = {dma_mem_ecc[13:7],io_dma_mem_wdata[63:32],dma_mem_ecc[6:0],io_dma_mem_wdata[31:0]}; // @[Cat.scala 29:58]
  reg [1:0] dma_mem_addr_ff; // @[el2_ifu_mem_ctl.scala 653:53]
  wire  _T_3585 = _T_3497[5:0] == 6'h27; // @[el2_lib.scala 324:41]
  wire  _T_3583 = _T_3497[5:0] == 6'h26; // @[el2_lib.scala 324:41]
  wire  _T_3581 = _T_3497[5:0] == 6'h25; // @[el2_lib.scala 324:41]
  wire  _T_3579 = _T_3497[5:0] == 6'h24; // @[el2_lib.scala 324:41]
  wire  _T_3577 = _T_3497[5:0] == 6'h23; // @[el2_lib.scala 324:41]
  wire  _T_3575 = _T_3497[5:0] == 6'h22; // @[el2_lib.scala 324:41]
  wire  _T_3573 = _T_3497[5:0] == 6'h21; // @[el2_lib.scala 324:41]
  wire  _T_3571 = _T_3497[5:0] == 6'h20; // @[el2_lib.scala 324:41]
  wire  _T_3569 = _T_3497[5:0] == 6'h1f; // @[el2_lib.scala 324:41]
  wire  _T_3567 = _T_3497[5:0] == 6'h1e; // @[el2_lib.scala 324:41]
  wire [9:0] _T_3643 = {_T_3585,_T_3583,_T_3581,_T_3579,_T_3577,_T_3575,_T_3573,_T_3571,_T_3569,_T_3567}; // @[el2_lib.scala 327:69]
  wire  _T_3565 = _T_3497[5:0] == 6'h1d; // @[el2_lib.scala 324:41]
  wire  _T_3563 = _T_3497[5:0] == 6'h1c; // @[el2_lib.scala 324:41]
  wire  _T_3561 = _T_3497[5:0] == 6'h1b; // @[el2_lib.scala 324:41]
  wire  _T_3559 = _T_3497[5:0] == 6'h1a; // @[el2_lib.scala 324:41]
  wire  _T_3557 = _T_3497[5:0] == 6'h19; // @[el2_lib.scala 324:41]
  wire  _T_3555 = _T_3497[5:0] == 6'h18; // @[el2_lib.scala 324:41]
  wire  _T_3553 = _T_3497[5:0] == 6'h17; // @[el2_lib.scala 324:41]
  wire  _T_3551 = _T_3497[5:0] == 6'h16; // @[el2_lib.scala 324:41]
  wire  _T_3549 = _T_3497[5:0] == 6'h15; // @[el2_lib.scala 324:41]
  wire  _T_3547 = _T_3497[5:0] == 6'h14; // @[el2_lib.scala 324:41]
  wire [9:0] _T_3634 = {_T_3565,_T_3563,_T_3561,_T_3559,_T_3557,_T_3555,_T_3553,_T_3551,_T_3549,_T_3547}; // @[el2_lib.scala 327:69]
  wire  _T_3545 = _T_3497[5:0] == 6'h13; // @[el2_lib.scala 324:41]
  wire  _T_3543 = _T_3497[5:0] == 6'h12; // @[el2_lib.scala 324:41]
  wire  _T_3541 = _T_3497[5:0] == 6'h11; // @[el2_lib.scala 324:41]
  wire  _T_3539 = _T_3497[5:0] == 6'h10; // @[el2_lib.scala 324:41]
  wire  _T_3537 = _T_3497[5:0] == 6'hf; // @[el2_lib.scala 324:41]
  wire  _T_3535 = _T_3497[5:0] == 6'he; // @[el2_lib.scala 324:41]
  wire  _T_3533 = _T_3497[5:0] == 6'hd; // @[el2_lib.scala 324:41]
  wire  _T_3531 = _T_3497[5:0] == 6'hc; // @[el2_lib.scala 324:41]
  wire  _T_3529 = _T_3497[5:0] == 6'hb; // @[el2_lib.scala 324:41]
  wire  _T_3527 = _T_3497[5:0] == 6'ha; // @[el2_lib.scala 324:41]
  wire [9:0] _T_3624 = {_T_3545,_T_3543,_T_3541,_T_3539,_T_3537,_T_3535,_T_3533,_T_3531,_T_3529,_T_3527}; // @[el2_lib.scala 327:69]
  wire  _T_3525 = _T_3497[5:0] == 6'h9; // @[el2_lib.scala 324:41]
  wire  _T_3523 = _T_3497[5:0] == 6'h8; // @[el2_lib.scala 324:41]
  wire  _T_3521 = _T_3497[5:0] == 6'h7; // @[el2_lib.scala 324:41]
  wire  _T_3519 = _T_3497[5:0] == 6'h6; // @[el2_lib.scala 324:41]
  wire  _T_3517 = _T_3497[5:0] == 6'h5; // @[el2_lib.scala 324:41]
  wire  _T_3515 = _T_3497[5:0] == 6'h4; // @[el2_lib.scala 324:41]
  wire  _T_3513 = _T_3497[5:0] == 6'h3; // @[el2_lib.scala 324:41]
  wire  _T_3511 = _T_3497[5:0] == 6'h2; // @[el2_lib.scala 324:41]
  wire  _T_3509 = _T_3497[5:0] == 6'h1; // @[el2_lib.scala 324:41]
  wire [18:0] _T_3625 = {_T_3624,_T_3525,_T_3523,_T_3521,_T_3519,_T_3517,_T_3515,_T_3513,_T_3511,_T_3509}; // @[el2_lib.scala 327:69]
  wire [38:0] _T_3645 = {_T_3643,_T_3634,_T_3625}; // @[el2_lib.scala 327:69]
  wire [7:0] _T_3600 = {io_iccm_rd_data_ecc[35],io_iccm_rd_data_ecc[3:1],io_iccm_rd_data_ecc[34],io_iccm_rd_data_ecc[0],io_iccm_rd_data_ecc[33:32]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3606 = {io_iccm_rd_data_ecc[38],io_iccm_rd_data_ecc[31:26],io_iccm_rd_data_ecc[37],io_iccm_rd_data_ecc[25:11],io_iccm_rd_data_ecc[36],io_iccm_rd_data_ecc[10:4],_T_3600}; // @[Cat.scala 29:58]
  wire [38:0] _T_3646 = _T_3645 ^ _T_3606; // @[el2_lib.scala 327:76]
  wire [38:0] _T_3647 = _T_3501 ? _T_3646 : _T_3606; // @[el2_lib.scala 327:31]
  wire [31:0] iccm_corrected_data_0 = {_T_3647[37:32],_T_3647[30:16],_T_3647[14:8],_T_3647[6:4],_T_3647[2]}; // @[Cat.scala 29:58]
  wire  _T_3970 = _T_3882[5:0] == 6'h27; // @[el2_lib.scala 324:41]
  wire  _T_3968 = _T_3882[5:0] == 6'h26; // @[el2_lib.scala 324:41]
  wire  _T_3966 = _T_3882[5:0] == 6'h25; // @[el2_lib.scala 324:41]
  wire  _T_3964 = _T_3882[5:0] == 6'h24; // @[el2_lib.scala 324:41]
  wire  _T_3962 = _T_3882[5:0] == 6'h23; // @[el2_lib.scala 324:41]
  wire  _T_3960 = _T_3882[5:0] == 6'h22; // @[el2_lib.scala 324:41]
  wire  _T_3958 = _T_3882[5:0] == 6'h21; // @[el2_lib.scala 324:41]
  wire  _T_3956 = _T_3882[5:0] == 6'h20; // @[el2_lib.scala 324:41]
  wire  _T_3954 = _T_3882[5:0] == 6'h1f; // @[el2_lib.scala 324:41]
  wire  _T_3952 = _T_3882[5:0] == 6'h1e; // @[el2_lib.scala 324:41]
  wire [9:0] _T_4028 = {_T_3970,_T_3968,_T_3966,_T_3964,_T_3962,_T_3960,_T_3958,_T_3956,_T_3954,_T_3952}; // @[el2_lib.scala 327:69]
  wire  _T_3950 = _T_3882[5:0] == 6'h1d; // @[el2_lib.scala 324:41]
  wire  _T_3948 = _T_3882[5:0] == 6'h1c; // @[el2_lib.scala 324:41]
  wire  _T_3946 = _T_3882[5:0] == 6'h1b; // @[el2_lib.scala 324:41]
  wire  _T_3944 = _T_3882[5:0] == 6'h1a; // @[el2_lib.scala 324:41]
  wire  _T_3942 = _T_3882[5:0] == 6'h19; // @[el2_lib.scala 324:41]
  wire  _T_3940 = _T_3882[5:0] == 6'h18; // @[el2_lib.scala 324:41]
  wire  _T_3938 = _T_3882[5:0] == 6'h17; // @[el2_lib.scala 324:41]
  wire  _T_3936 = _T_3882[5:0] == 6'h16; // @[el2_lib.scala 324:41]
  wire  _T_3934 = _T_3882[5:0] == 6'h15; // @[el2_lib.scala 324:41]
  wire  _T_3932 = _T_3882[5:0] == 6'h14; // @[el2_lib.scala 324:41]
  wire [9:0] _T_4019 = {_T_3950,_T_3948,_T_3946,_T_3944,_T_3942,_T_3940,_T_3938,_T_3936,_T_3934,_T_3932}; // @[el2_lib.scala 327:69]
  wire  _T_3930 = _T_3882[5:0] == 6'h13; // @[el2_lib.scala 324:41]
  wire  _T_3928 = _T_3882[5:0] == 6'h12; // @[el2_lib.scala 324:41]
  wire  _T_3926 = _T_3882[5:0] == 6'h11; // @[el2_lib.scala 324:41]
  wire  _T_3924 = _T_3882[5:0] == 6'h10; // @[el2_lib.scala 324:41]
  wire  _T_3922 = _T_3882[5:0] == 6'hf; // @[el2_lib.scala 324:41]
  wire  _T_3920 = _T_3882[5:0] == 6'he; // @[el2_lib.scala 324:41]
  wire  _T_3918 = _T_3882[5:0] == 6'hd; // @[el2_lib.scala 324:41]
  wire  _T_3916 = _T_3882[5:0] == 6'hc; // @[el2_lib.scala 324:41]
  wire  _T_3914 = _T_3882[5:0] == 6'hb; // @[el2_lib.scala 324:41]
  wire  _T_3912 = _T_3882[5:0] == 6'ha; // @[el2_lib.scala 324:41]
  wire [9:0] _T_4009 = {_T_3930,_T_3928,_T_3926,_T_3924,_T_3922,_T_3920,_T_3918,_T_3916,_T_3914,_T_3912}; // @[el2_lib.scala 327:69]
  wire  _T_3910 = _T_3882[5:0] == 6'h9; // @[el2_lib.scala 324:41]
  wire  _T_3908 = _T_3882[5:0] == 6'h8; // @[el2_lib.scala 324:41]
  wire  _T_3906 = _T_3882[5:0] == 6'h7; // @[el2_lib.scala 324:41]
  wire  _T_3904 = _T_3882[5:0] == 6'h6; // @[el2_lib.scala 324:41]
  wire  _T_3902 = _T_3882[5:0] == 6'h5; // @[el2_lib.scala 324:41]
  wire  _T_3900 = _T_3882[5:0] == 6'h4; // @[el2_lib.scala 324:41]
  wire  _T_3898 = _T_3882[5:0] == 6'h3; // @[el2_lib.scala 324:41]
  wire  _T_3896 = _T_3882[5:0] == 6'h2; // @[el2_lib.scala 324:41]
  wire  _T_3894 = _T_3882[5:0] == 6'h1; // @[el2_lib.scala 324:41]
  wire [18:0] _T_4010 = {_T_4009,_T_3910,_T_3908,_T_3906,_T_3904,_T_3902,_T_3900,_T_3898,_T_3896,_T_3894}; // @[el2_lib.scala 327:69]
  wire [38:0] _T_4030 = {_T_4028,_T_4019,_T_4010}; // @[el2_lib.scala 327:69]
  wire [7:0] _T_3985 = {io_iccm_rd_data_ecc[74],io_iccm_rd_data_ecc[42:40],io_iccm_rd_data_ecc[73],io_iccm_rd_data_ecc[39],io_iccm_rd_data_ecc[72:71]}; // @[Cat.scala 29:58]
  wire [38:0] _T_3991 = {io_iccm_rd_data_ecc[77],io_iccm_rd_data_ecc[70:65],io_iccm_rd_data_ecc[76],io_iccm_rd_data_ecc[64:50],io_iccm_rd_data_ecc[75],io_iccm_rd_data_ecc[49:43],_T_3985}; // @[Cat.scala 29:58]
  wire [38:0] _T_4031 = _T_4030 ^ _T_3991; // @[el2_lib.scala 327:76]
  wire [38:0] _T_4032 = _T_3886 ? _T_4031 : _T_3991; // @[el2_lib.scala 327:31]
  wire [31:0] iccm_corrected_data_1 = {_T_4032[37:32],_T_4032[30:16],_T_4032[14:8],_T_4032[6:4],_T_4032[2]}; // @[Cat.scala 29:58]
  wire [31:0] iccm_dma_rdata_1_muxed = dma_mem_addr_ff[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 645:35]
  wire  _T_3505 = ~_T_3497[6]; // @[el2_lib.scala 320:55]
  wire  _T_3506 = _T_3499 & _T_3505; // @[el2_lib.scala 320:53]
  wire  _T_3890 = ~_T_3882[6]; // @[el2_lib.scala 320:55]
  wire  _T_3891 = _T_3884 & _T_3890; // @[el2_lib.scala 320:53]
  wire [1:0] iccm_double_ecc_error = {_T_3506,_T_3891}; // @[Cat.scala 29:58]
  wire  iccm_dma_ecc_error_in = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 647:53]
  wire [63:0] _T_3257 = {io_dma_mem_addr,io_dma_mem_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_3258 = {iccm_dma_rdata_1_muxed,_T_3647[37:32],_T_3647[30:16],_T_3647[14:8],_T_3647[6:4],_T_3647[2]}; // @[Cat.scala 29:58]
  reg [2:0] dma_mem_tag_ff; // @[el2_ifu_mem_ctl.scala 649:54]
  reg [2:0] iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 650:74]
  reg  iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 655:76]
  reg [63:0] iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 659:75]
  wire  _T_3263 = _T_2678 & _T_2667; // @[el2_ifu_mem_ctl.scala 662:65]
  wire  _T_3266 = _T_3244 & iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 663:50]
  reg [13:0] iccm_ecc_corr_index_ff; // @[Reg.scala 27:20]
  wire [14:0] _T_3267 = {iccm_ecc_corr_index_ff,1'h0}; // @[Cat.scala 29:58]
  wire [15:0] _T_3269 = _T_3266 ? {{1'd0}, _T_3267} : io_ifc_fetch_addr_bf[15:0]; // @[el2_ifu_mem_ctl.scala 663:8]
  wire [31:0] _T_3270 = _T_3263 ? io_dma_mem_addr : {{16'd0}, _T_3269}; // @[el2_ifu_mem_ctl.scala 662:25]
  wire  _T_3659 = _T_3497 == 7'h40; // @[el2_lib.scala 330:62]
  wire  _T_3660 = _T_3647[38] ^ _T_3659; // @[el2_lib.scala 330:44]
  wire [6:0] iccm_corrected_ecc_0 = {_T_3660,_T_3647[31],_T_3647[15],_T_3647[7],_T_3647[3],_T_3647[1:0]}; // @[Cat.scala 29:58]
  wire  _T_4044 = _T_3882 == 7'h40; // @[el2_lib.scala 330:62]
  wire  _T_4045 = _T_4032[38] ^ _T_4044; // @[el2_lib.scala 330:44]
  wire [6:0] iccm_corrected_ecc_1 = {_T_4045,_T_4032[31],_T_4032[15],_T_4032[7],_T_4032[3],_T_4032[1:0]}; // @[Cat.scala 29:58]
  wire  _T_4061 = _T_3 & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 675:58]
  wire [31:0] iccm_corrected_data_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_data_0 : iccm_corrected_data_1; // @[el2_ifu_mem_ctl.scala 677:38]
  wire [6:0] iccm_corrected_ecc_f_mux = iccm_single_ecc_error[0] ? iccm_corrected_ecc_0 : iccm_corrected_ecc_1; // @[el2_ifu_mem_ctl.scala 678:37]
  reg  iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 686:62]
  wire  _T_4069 = ~iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 680:76]
  wire  _T_4070 = io_iccm_rd_ecc_single_err & _T_4069; // @[el2_ifu_mem_ctl.scala 680:74]
  wire  _T_4072 = _T_4070 & _T_317; // @[el2_ifu_mem_ctl.scala 680:104]
  wire  iccm_ecc_write_status = _T_4072 | io_iccm_dma_sb_error; // @[el2_ifu_mem_ctl.scala 680:127]
  wire  _T_4073 = io_iccm_rd_ecc_single_err | iccm_rd_ecc_single_err_ff; // @[el2_ifu_mem_ctl.scala 681:67]
  wire  iccm_rd_ecc_single_err_hold_in = _T_4073 & _T_317; // @[el2_ifu_mem_ctl.scala 681:96]
  reg [13:0] iccm_rw_addr_f; // @[el2_ifu_mem_ctl.scala 685:51]
  wire [13:0] _T_4078 = iccm_rw_addr_f + 14'h1; // @[el2_ifu_mem_ctl.scala 684:102]
  wire [38:0] _T_4082 = {iccm_corrected_ecc_f_mux,iccm_corrected_data_f_mux}; // @[Cat.scala 29:58]
  wire  _T_4087 = ~io_ifc_fetch_uncacheable_bf; // @[el2_ifu_mem_ctl.scala 689:41]
  wire  _T_4088 = io_ifc_fetch_req_bf & _T_4087; // @[el2_ifu_mem_ctl.scala 689:39]
  wire  _T_4089 = ~io_ifc_iccm_access_bf; // @[el2_ifu_mem_ctl.scala 689:72]
  wire  _T_4090 = _T_4088 & _T_4089; // @[el2_ifu_mem_ctl.scala 689:70]
  wire  _T_4092 = ~miss_state_en; // @[el2_ifu_mem_ctl.scala 690:34]
  wire  _T_4093 = _T_2233 & _T_4092; // @[el2_ifu_mem_ctl.scala 690:32]
  wire  _T_4096 = _T_2249 & _T_4092; // @[el2_ifu_mem_ctl.scala 691:37]
  wire  _T_4097 = _T_4093 | _T_4096; // @[el2_ifu_mem_ctl.scala 690:88]
  wire  _T_4098 = miss_state == 3'h7; // @[el2_ifu_mem_ctl.scala 692:19]
  wire  _T_4100 = _T_4098 & _T_4092; // @[el2_ifu_mem_ctl.scala 692:41]
  wire  _T_4101 = _T_4097 | _T_4100; // @[el2_ifu_mem_ctl.scala 691:88]
  wire  _T_4102 = miss_state == 3'h3; // @[el2_ifu_mem_ctl.scala 693:19]
  wire  _T_4104 = _T_4102 & _T_4092; // @[el2_ifu_mem_ctl.scala 693:35]
  wire  _T_4105 = _T_4101 | _T_4104; // @[el2_ifu_mem_ctl.scala 692:88]
  wire  _T_4108 = _T_2248 & _T_4092; // @[el2_ifu_mem_ctl.scala 694:38]
  wire  _T_4109 = _T_4105 | _T_4108; // @[el2_ifu_mem_ctl.scala 693:88]
  wire  _T_4111 = _T_2249 & miss_state_en; // @[el2_ifu_mem_ctl.scala 695:37]
  wire  _T_4112 = miss_nxtstate == 3'h3; // @[el2_ifu_mem_ctl.scala 695:71]
  wire  _T_4113 = _T_4111 & _T_4112; // @[el2_ifu_mem_ctl.scala 695:54]
  wire  _T_4114 = _T_4109 | _T_4113; // @[el2_ifu_mem_ctl.scala 694:57]
  wire  _T_4115 = ~_T_4114; // @[el2_ifu_mem_ctl.scala 690:5]
  wire  _T_4116 = _T_4090 & _T_4115; // @[el2_ifu_mem_ctl.scala 689:96]
  wire  _T_4117 = io_ifc_fetch_req_bf & io_exu_flush_final; // @[el2_ifu_mem_ctl.scala 696:28]
  wire  _T_4119 = _T_4117 & _T_4087; // @[el2_ifu_mem_ctl.scala 696:50]
  wire  _T_4121 = _T_4119 & _T_4089; // @[el2_ifu_mem_ctl.scala 696:81]
  wire [1:0] _T_4124 = write_ic_16_bytes ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire  _T_10562 = bus_ifu_wr_en_ff_q & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 793:74]
  wire  bus_wren_1 = _T_10562 & miss_pending; // @[el2_ifu_mem_ctl.scala 793:98]
  wire  _T_10561 = bus_ifu_wr_en_ff_q & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 793:74]
  wire  bus_wren_0 = _T_10561 & miss_pending; // @[el2_ifu_mem_ctl.scala 793:98]
  wire [1:0] bus_ic_wr_en = {bus_wren_1,bus_wren_0}; // @[Cat.scala 29:58]
  wire  _T_4130 = ~_T_108; // @[el2_ifu_mem_ctl.scala 699:106]
  wire  _T_4131 = _T_2233 & _T_4130; // @[el2_ifu_mem_ctl.scala 699:104]
  wire  _T_4132 = _T_2249 | _T_4131; // @[el2_ifu_mem_ctl.scala 699:77]
  wire  _T_4136 = ~_T_51; // @[el2_ifu_mem_ctl.scala 699:172]
  wire  _T_4137 = _T_4132 & _T_4136; // @[el2_ifu_mem_ctl.scala 699:170]
  wire  _T_4138 = ~_T_4137; // @[el2_ifu_mem_ctl.scala 699:44]
  wire  _T_4142 = reset_ic_in | reset_ic_ff; // @[el2_ifu_mem_ctl.scala 702:64]
  wire  _T_4143 = ~_T_4142; // @[el2_ifu_mem_ctl.scala 702:50]
  wire  _T_4144 = _T_276 & _T_4143; // @[el2_ifu_mem_ctl.scala 702:48]
  wire  _T_4145 = ~reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 702:81]
  wire  ic_valid = _T_4144 & _T_4145; // @[el2_ifu_mem_ctl.scala 702:79]
  wire  _T_4147 = debug_c1_clken & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 703:82]
  reg [6:0] ifu_status_wr_addr_ff; // @[el2_ifu_mem_ctl.scala 706:14]
  wire  _T_4150 = io_ic_debug_wr_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 709:74]
  wire  _T_10559 = bus_ifu_wr_en_ff_q & last_beat; // @[el2_ifu_mem_ctl.scala 792:45]
  wire  way_status_wr_en = _T_10559 | ic_act_hit_f; // @[el2_ifu_mem_ctl.scala 792:58]
  wire  way_status_wr_en_w_debug = way_status_wr_en | _T_4150; // @[el2_ifu_mem_ctl.scala 709:53]
  reg  way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 711:14]
  wire  way_status_hit_new = io_ic_rd_hit[0]; // @[el2_ifu_mem_ctl.scala 788:41]
  reg  way_status_new_ff; // @[el2_ifu_mem_ctl.scala 719:14]
  wire  way_status_clken_0 = ifu_status_wr_addr_ff[6:3] == 4'h0; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_1 = ifu_status_wr_addr_ff[6:3] == 4'h1; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_2 = ifu_status_wr_addr_ff[6:3] == 4'h2; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_3 = ifu_status_wr_addr_ff[6:3] == 4'h3; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_4 = ifu_status_wr_addr_ff[6:3] == 4'h4; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_5 = ifu_status_wr_addr_ff[6:3] == 4'h5; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_6 = ifu_status_wr_addr_ff[6:3] == 4'h6; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_7 = ifu_status_wr_addr_ff[6:3] == 4'h7; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_8 = ifu_status_wr_addr_ff[6:3] == 4'h8; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_9 = ifu_status_wr_addr_ff[6:3] == 4'h9; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_10 = ifu_status_wr_addr_ff[6:3] == 4'ha; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_11 = ifu_status_wr_addr_ff[6:3] == 4'hb; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_12 = ifu_status_wr_addr_ff[6:3] == 4'hc; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_13 = ifu_status_wr_addr_ff[6:3] == 4'hd; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_14 = ifu_status_wr_addr_ff[6:3] == 4'he; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  way_status_clken_15 = ifu_status_wr_addr_ff[6:3] == 4'hf; // @[el2_ifu_mem_ctl.scala 721:132]
  wire  _T_4170 = ifu_status_wr_addr_ff[2:0] == 3'h0; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4171 = _T_4170 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4172 = _T_4171 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4175 = ifu_status_wr_addr_ff[2:0] == 3'h1; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4176 = _T_4175 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4177 = _T_4176 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4180 = ifu_status_wr_addr_ff[2:0] == 3'h2; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4181 = _T_4180 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4182 = _T_4181 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4185 = ifu_status_wr_addr_ff[2:0] == 3'h3; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4186 = _T_4185 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4187 = _T_4186 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4190 = ifu_status_wr_addr_ff[2:0] == 3'h4; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4191 = _T_4190 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4192 = _T_4191 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4195 = ifu_status_wr_addr_ff[2:0] == 3'h5; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4196 = _T_4195 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4197 = _T_4196 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4200 = ifu_status_wr_addr_ff[2:0] == 3'h6; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4201 = _T_4200 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4202 = _T_4201 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4205 = ifu_status_wr_addr_ff[2:0] == 3'h7; // @[el2_ifu_mem_ctl.scala 725:100]
  wire  _T_4206 = _T_4205 & way_status_wr_en_ff; // @[el2_ifu_mem_ctl.scala 725:108]
  wire  _T_4207 = _T_4206 & way_status_clken_0; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4212 = _T_4171 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4217 = _T_4176 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4222 = _T_4181 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4227 = _T_4186 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4232 = _T_4191 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4237 = _T_4196 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4242 = _T_4201 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4247 = _T_4206 & way_status_clken_1; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4252 = _T_4171 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4257 = _T_4176 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4262 = _T_4181 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4267 = _T_4186 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4272 = _T_4191 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4277 = _T_4196 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4282 = _T_4201 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4287 = _T_4206 & way_status_clken_2; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4292 = _T_4171 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4297 = _T_4176 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4302 = _T_4181 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4307 = _T_4186 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4312 = _T_4191 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4317 = _T_4196 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4322 = _T_4201 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4327 = _T_4206 & way_status_clken_3; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4332 = _T_4171 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4337 = _T_4176 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4342 = _T_4181 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4347 = _T_4186 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4352 = _T_4191 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4357 = _T_4196 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4362 = _T_4201 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4367 = _T_4206 & way_status_clken_4; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4372 = _T_4171 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4377 = _T_4176 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4382 = _T_4181 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4387 = _T_4186 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4392 = _T_4191 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4397 = _T_4196 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4402 = _T_4201 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4407 = _T_4206 & way_status_clken_5; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4412 = _T_4171 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4417 = _T_4176 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4422 = _T_4181 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4427 = _T_4186 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4432 = _T_4191 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4437 = _T_4196 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4442 = _T_4201 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4447 = _T_4206 & way_status_clken_6; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4452 = _T_4171 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4457 = _T_4176 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4462 = _T_4181 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4467 = _T_4186 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4472 = _T_4191 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4477 = _T_4196 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4482 = _T_4201 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4487 = _T_4206 & way_status_clken_7; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4492 = _T_4171 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4497 = _T_4176 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4502 = _T_4181 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4507 = _T_4186 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4512 = _T_4191 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4517 = _T_4196 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4522 = _T_4201 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4527 = _T_4206 & way_status_clken_8; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4532 = _T_4171 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4537 = _T_4176 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4542 = _T_4181 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4547 = _T_4186 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4552 = _T_4191 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4557 = _T_4196 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4562 = _T_4201 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4567 = _T_4206 & way_status_clken_9; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4572 = _T_4171 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4577 = _T_4176 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4582 = _T_4181 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4587 = _T_4186 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4592 = _T_4191 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4597 = _T_4196 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4602 = _T_4201 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4607 = _T_4206 & way_status_clken_10; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4612 = _T_4171 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4617 = _T_4176 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4622 = _T_4181 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4627 = _T_4186 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4632 = _T_4191 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4637 = _T_4196 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4642 = _T_4201 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4647 = _T_4206 & way_status_clken_11; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4652 = _T_4171 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4657 = _T_4176 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4662 = _T_4181 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4667 = _T_4186 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4672 = _T_4191 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4677 = _T_4196 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4682 = _T_4201 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4687 = _T_4206 & way_status_clken_12; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4692 = _T_4171 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4697 = _T_4176 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4702 = _T_4181 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4707 = _T_4186 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4712 = _T_4191 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4717 = _T_4196 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4722 = _T_4201 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4727 = _T_4206 & way_status_clken_13; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4732 = _T_4171 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4737 = _T_4176 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4742 = _T_4181 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4747 = _T_4186 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4752 = _T_4191 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4757 = _T_4196 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4762 = _T_4201 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4767 = _T_4206 & way_status_clken_14; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4772 = _T_4171 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4777 = _T_4176 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4782 = _T_4181 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4787 = _T_4186 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4792 = _T_4191 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4797 = _T_4196 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4802 = _T_4201 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_4807 = _T_4206 & way_status_clken_15; // @[el2_ifu_mem_ctl.scala 725:131]
  wire  _T_10565 = _T_100 & replace_way_mb_any_1; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_10566 = _T_10565 & miss_pending; // @[el2_ifu_mem_ctl.scala 795:108]
  wire  bus_wren_last_1 = _T_10566 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 795:123]
  wire  wren_reset_miss_1 = replace_way_mb_any_1 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 796:84]
  wire  _T_10568 = bus_wren_last_1 | wren_reset_miss_1; // @[el2_ifu_mem_ctl.scala 797:73]
  wire  _T_10563 = _T_100 & replace_way_mb_any_0; // @[el2_ifu_mem_ctl.scala 795:84]
  wire  _T_10564 = _T_10563 & miss_pending; // @[el2_ifu_mem_ctl.scala 795:108]
  wire  bus_wren_last_0 = _T_10564 & bus_last_data_beat; // @[el2_ifu_mem_ctl.scala 795:123]
  wire  wren_reset_miss_0 = replace_way_mb_any_0 & reset_tag_valid_for_miss; // @[el2_ifu_mem_ctl.scala 796:84]
  wire  _T_10567 = bus_wren_last_0 | wren_reset_miss_0; // @[el2_ifu_mem_ctl.scala 797:73]
  wire [1:0] ifu_tag_wren = {_T_10568,_T_10567}; // @[Cat.scala 29:58]
  wire [1:0] _T_10603 = _T_4150 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  wire [1:0] ic_debug_tag_wr_en = _T_10603 & io_ic_debug_way; // @[el2_ifu_mem_ctl.scala 831:90]
  wire [1:0] ifu_tag_wren_w_debug = ifu_tag_wren | ic_debug_tag_wr_en; // @[el2_ifu_mem_ctl.scala 738:45]
  reg [1:0] ifu_tag_wren_ff; // @[el2_ifu_mem_ctl.scala 740:14]
  reg  ic_valid_ff; // @[el2_ifu_mem_ctl.scala 744:14]
  wire  _T_5341 = ifu_ic_rw_int_addr_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5343 = _T_5341 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5345 = perr_ic_index_ff[6:5] == 2'h0; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5347 = _T_5345 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5348 = _T_5343 | _T_5347; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5349 = _T_5348 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5353 = _T_5341 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5357 = _T_5345 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5358 = _T_5353 | _T_5357; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5359 = _T_5358 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_0 = {_T_5359,_T_5349}; // @[Cat.scala 29:58]
  wire  _T_5361 = ifu_ic_rw_int_addr_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5363 = _T_5361 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5365 = perr_ic_index_ff[6:5] == 2'h1; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5367 = _T_5365 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5368 = _T_5363 | _T_5367; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5369 = _T_5368 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5373 = _T_5361 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5377 = _T_5365 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5378 = _T_5373 | _T_5377; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5379 = _T_5378 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_1 = {_T_5379,_T_5369}; // @[Cat.scala 29:58]
  wire  _T_5381 = ifu_ic_rw_int_addr_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5383 = _T_5381 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5385 = perr_ic_index_ff[6:5] == 2'h2; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5387 = _T_5385 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5388 = _T_5383 | _T_5387; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5389 = _T_5388 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5393 = _T_5381 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5397 = _T_5385 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5398 = _T_5393 | _T_5397; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5399 = _T_5398 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_2 = {_T_5399,_T_5389}; // @[Cat.scala 29:58]
  wire  _T_5401 = ifu_ic_rw_int_addr_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 748:78]
  wire  _T_5403 = _T_5401 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5405 = perr_ic_index_ff[6:5] == 2'h3; // @[el2_ifu_mem_ctl.scala 749:70]
  wire  _T_5407 = _T_5405 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5408 = _T_5403 | _T_5407; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5409 = _T_5408 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire  _T_5413 = _T_5401 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 748:87]
  wire  _T_5417 = _T_5405 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 749:79]
  wire  _T_5418 = _T_5413 | _T_5417; // @[el2_ifu_mem_ctl.scala 748:109]
  wire  _T_5419 = _T_5418 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 749:102]
  wire [1:0] tag_valid_clken_3 = {_T_5419,_T_5409}; // @[Cat.scala 29:58]
  wire  _T_5422 = ic_valid_ff & _T_195; // @[el2_ifu_mem_ctl.scala 757:66]
  wire  _T_5423 = ~perr_sel_invalidate; // @[el2_ifu_mem_ctl.scala 757:93]
  wire  _T_5424 = _T_5422 & _T_5423; // @[el2_ifu_mem_ctl.scala 757:91]
  wire  _T_5427 = _T_4949 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5428 = perr_ic_index_ff == 7'h0; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5430 = _T_5428 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5431 = _T_5427 | _T_5430; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5432 = _T_5431 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5434 = _T_5432 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5444 = _T_4950 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5445 = perr_ic_index_ff == 7'h1; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5447 = _T_5445 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5448 = _T_5444 | _T_5447; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5449 = _T_5448 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5451 = _T_5449 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5461 = _T_4951 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5462 = perr_ic_index_ff == 7'h2; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5464 = _T_5462 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5465 = _T_5461 | _T_5464; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5466 = _T_5465 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5468 = _T_5466 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5478 = _T_4952 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5479 = perr_ic_index_ff == 7'h3; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5481 = _T_5479 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5482 = _T_5478 | _T_5481; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5483 = _T_5482 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5485 = _T_5483 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5495 = _T_4953 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5496 = perr_ic_index_ff == 7'h4; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5498 = _T_5496 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5499 = _T_5495 | _T_5498; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5500 = _T_5499 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5502 = _T_5500 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5512 = _T_4954 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5513 = perr_ic_index_ff == 7'h5; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5515 = _T_5513 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5516 = _T_5512 | _T_5515; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5517 = _T_5516 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5519 = _T_5517 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5529 = _T_4955 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5530 = perr_ic_index_ff == 7'h6; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5532 = _T_5530 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5533 = _T_5529 | _T_5532; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5534 = _T_5533 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5536 = _T_5534 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5546 = _T_4956 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5547 = perr_ic_index_ff == 7'h7; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5549 = _T_5547 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5550 = _T_5546 | _T_5549; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5551 = _T_5550 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5553 = _T_5551 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5563 = _T_4957 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5564 = perr_ic_index_ff == 7'h8; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5566 = _T_5564 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5567 = _T_5563 | _T_5566; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5568 = _T_5567 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5570 = _T_5568 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5580 = _T_4958 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5581 = perr_ic_index_ff == 7'h9; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5583 = _T_5581 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5584 = _T_5580 | _T_5583; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5585 = _T_5584 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5587 = _T_5585 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5597 = _T_4959 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5598 = perr_ic_index_ff == 7'ha; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5600 = _T_5598 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5601 = _T_5597 | _T_5600; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5602 = _T_5601 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5604 = _T_5602 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5614 = _T_4960 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5615 = perr_ic_index_ff == 7'hb; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5617 = _T_5615 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5618 = _T_5614 | _T_5617; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5619 = _T_5618 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5621 = _T_5619 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5631 = _T_4961 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5632 = perr_ic_index_ff == 7'hc; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5634 = _T_5632 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5635 = _T_5631 | _T_5634; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5636 = _T_5635 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5638 = _T_5636 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5648 = _T_4962 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5649 = perr_ic_index_ff == 7'hd; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5651 = _T_5649 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5652 = _T_5648 | _T_5651; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5653 = _T_5652 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5655 = _T_5653 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5665 = _T_4963 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5666 = perr_ic_index_ff == 7'he; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5668 = _T_5666 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5669 = _T_5665 | _T_5668; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5670 = _T_5669 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5672 = _T_5670 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5682 = _T_4964 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5683 = perr_ic_index_ff == 7'hf; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5685 = _T_5683 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5686 = _T_5682 | _T_5685; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5687 = _T_5686 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5689 = _T_5687 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5699 = _T_4965 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5700 = perr_ic_index_ff == 7'h10; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5702 = _T_5700 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5703 = _T_5699 | _T_5702; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5704 = _T_5703 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5706 = _T_5704 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5716 = _T_4966 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5717 = perr_ic_index_ff == 7'h11; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5719 = _T_5717 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5720 = _T_5716 | _T_5719; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5721 = _T_5720 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5723 = _T_5721 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5733 = _T_4967 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5734 = perr_ic_index_ff == 7'h12; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5736 = _T_5734 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5737 = _T_5733 | _T_5736; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5738 = _T_5737 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5740 = _T_5738 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5750 = _T_4968 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5751 = perr_ic_index_ff == 7'h13; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5753 = _T_5751 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5754 = _T_5750 | _T_5753; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5755 = _T_5754 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5757 = _T_5755 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5767 = _T_4969 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5768 = perr_ic_index_ff == 7'h14; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5770 = _T_5768 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5771 = _T_5767 | _T_5770; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5772 = _T_5771 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5774 = _T_5772 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5784 = _T_4970 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5785 = perr_ic_index_ff == 7'h15; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5787 = _T_5785 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5788 = _T_5784 | _T_5787; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5789 = _T_5788 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5791 = _T_5789 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5801 = _T_4971 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5802 = perr_ic_index_ff == 7'h16; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5804 = _T_5802 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5805 = _T_5801 | _T_5804; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5806 = _T_5805 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5808 = _T_5806 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5818 = _T_4972 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5819 = perr_ic_index_ff == 7'h17; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5821 = _T_5819 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5822 = _T_5818 | _T_5821; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5823 = _T_5822 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5825 = _T_5823 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5835 = _T_4973 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5836 = perr_ic_index_ff == 7'h18; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5838 = _T_5836 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5839 = _T_5835 | _T_5838; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5840 = _T_5839 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5842 = _T_5840 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5852 = _T_4974 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5853 = perr_ic_index_ff == 7'h19; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5855 = _T_5853 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5856 = _T_5852 | _T_5855; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5857 = _T_5856 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5859 = _T_5857 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5869 = _T_4975 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5870 = perr_ic_index_ff == 7'h1a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5872 = _T_5870 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5873 = _T_5869 | _T_5872; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5874 = _T_5873 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5876 = _T_5874 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5886 = _T_4976 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5887 = perr_ic_index_ff == 7'h1b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5889 = _T_5887 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5890 = _T_5886 | _T_5889; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5891 = _T_5890 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5893 = _T_5891 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5903 = _T_4977 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5904 = perr_ic_index_ff == 7'h1c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5906 = _T_5904 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5907 = _T_5903 | _T_5906; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5908 = _T_5907 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5910 = _T_5908 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5920 = _T_4978 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5921 = perr_ic_index_ff == 7'h1d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5923 = _T_5921 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5924 = _T_5920 | _T_5923; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5925 = _T_5924 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5927 = _T_5925 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5937 = _T_4979 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5938 = perr_ic_index_ff == 7'h1e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5940 = _T_5938 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5941 = _T_5937 | _T_5940; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5942 = _T_5941 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5944 = _T_5942 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5954 = _T_4980 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5955 = perr_ic_index_ff == 7'h1f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_5957 = _T_5955 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5958 = _T_5954 | _T_5957; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5959 = _T_5958 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5961 = _T_5959 & tag_valid_clken_0[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5971 = _T_4949 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5974 = _T_5428 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5975 = _T_5971 | _T_5974; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5976 = _T_5975 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5978 = _T_5976 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_5988 = _T_4950 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_5991 = _T_5445 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_5992 = _T_5988 | _T_5991; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_5993 = _T_5992 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_5995 = _T_5993 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6005 = _T_4951 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6008 = _T_5462 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6009 = _T_6005 | _T_6008; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6010 = _T_6009 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6012 = _T_6010 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6022 = _T_4952 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6025 = _T_5479 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6026 = _T_6022 | _T_6025; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6027 = _T_6026 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6029 = _T_6027 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6039 = _T_4953 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6042 = _T_5496 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6043 = _T_6039 | _T_6042; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6044 = _T_6043 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6046 = _T_6044 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6056 = _T_4954 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6059 = _T_5513 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6060 = _T_6056 | _T_6059; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6061 = _T_6060 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6063 = _T_6061 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6073 = _T_4955 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6076 = _T_5530 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6077 = _T_6073 | _T_6076; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6078 = _T_6077 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6080 = _T_6078 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6090 = _T_4956 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6093 = _T_5547 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6094 = _T_6090 | _T_6093; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6095 = _T_6094 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6097 = _T_6095 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6107 = _T_4957 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6110 = _T_5564 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6111 = _T_6107 | _T_6110; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6112 = _T_6111 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6114 = _T_6112 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6124 = _T_4958 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6127 = _T_5581 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6128 = _T_6124 | _T_6127; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6129 = _T_6128 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6131 = _T_6129 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6141 = _T_4959 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6144 = _T_5598 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6145 = _T_6141 | _T_6144; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6146 = _T_6145 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6148 = _T_6146 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6158 = _T_4960 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6161 = _T_5615 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6162 = _T_6158 | _T_6161; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6163 = _T_6162 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6165 = _T_6163 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6175 = _T_4961 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6178 = _T_5632 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6179 = _T_6175 | _T_6178; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6180 = _T_6179 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6182 = _T_6180 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6192 = _T_4962 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6195 = _T_5649 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6196 = _T_6192 | _T_6195; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6197 = _T_6196 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6199 = _T_6197 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6209 = _T_4963 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6212 = _T_5666 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6213 = _T_6209 | _T_6212; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6214 = _T_6213 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6216 = _T_6214 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6226 = _T_4964 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6229 = _T_5683 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6230 = _T_6226 | _T_6229; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6231 = _T_6230 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6233 = _T_6231 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6243 = _T_4965 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6246 = _T_5700 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6247 = _T_6243 | _T_6246; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6248 = _T_6247 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6250 = _T_6248 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6260 = _T_4966 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6263 = _T_5717 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6264 = _T_6260 | _T_6263; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6265 = _T_6264 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6267 = _T_6265 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6277 = _T_4967 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6280 = _T_5734 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6281 = _T_6277 | _T_6280; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6282 = _T_6281 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6284 = _T_6282 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6294 = _T_4968 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6297 = _T_5751 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6298 = _T_6294 | _T_6297; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6299 = _T_6298 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6301 = _T_6299 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6311 = _T_4969 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6314 = _T_5768 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6315 = _T_6311 | _T_6314; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6316 = _T_6315 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6318 = _T_6316 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6328 = _T_4970 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6331 = _T_5785 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6332 = _T_6328 | _T_6331; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6333 = _T_6332 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6335 = _T_6333 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6345 = _T_4971 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6348 = _T_5802 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6349 = _T_6345 | _T_6348; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6350 = _T_6349 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6352 = _T_6350 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6362 = _T_4972 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6365 = _T_5819 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6366 = _T_6362 | _T_6365; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6367 = _T_6366 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6369 = _T_6367 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6379 = _T_4973 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6382 = _T_5836 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6383 = _T_6379 | _T_6382; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6384 = _T_6383 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6386 = _T_6384 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6396 = _T_4974 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6399 = _T_5853 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6400 = _T_6396 | _T_6399; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6401 = _T_6400 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6403 = _T_6401 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6413 = _T_4975 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6416 = _T_5870 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6417 = _T_6413 | _T_6416; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6418 = _T_6417 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6420 = _T_6418 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6430 = _T_4976 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6433 = _T_5887 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6434 = _T_6430 | _T_6433; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6435 = _T_6434 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6437 = _T_6435 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6447 = _T_4977 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6450 = _T_5904 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6451 = _T_6447 | _T_6450; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6452 = _T_6451 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6454 = _T_6452 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6464 = _T_4978 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6467 = _T_5921 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6468 = _T_6464 | _T_6467; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6469 = _T_6468 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6471 = _T_6469 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6481 = _T_4979 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6484 = _T_5938 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6485 = _T_6481 | _T_6484; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6486 = _T_6485 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6488 = _T_6486 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6498 = _T_4980 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6501 = _T_5955 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6502 = _T_6498 | _T_6501; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6503 = _T_6502 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6505 = _T_6503 & tag_valid_clken_0[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6515 = _T_4981 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6516 = perr_ic_index_ff == 7'h20; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6518 = _T_6516 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6519 = _T_6515 | _T_6518; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6520 = _T_6519 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6522 = _T_6520 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6532 = _T_4982 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6533 = perr_ic_index_ff == 7'h21; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6535 = _T_6533 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6536 = _T_6532 | _T_6535; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6537 = _T_6536 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6539 = _T_6537 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6549 = _T_4983 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6550 = perr_ic_index_ff == 7'h22; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6552 = _T_6550 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6553 = _T_6549 | _T_6552; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6554 = _T_6553 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6556 = _T_6554 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6566 = _T_4984 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6567 = perr_ic_index_ff == 7'h23; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6569 = _T_6567 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6570 = _T_6566 | _T_6569; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6571 = _T_6570 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6573 = _T_6571 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6583 = _T_4985 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6584 = perr_ic_index_ff == 7'h24; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6586 = _T_6584 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6587 = _T_6583 | _T_6586; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6588 = _T_6587 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6590 = _T_6588 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6600 = _T_4986 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6601 = perr_ic_index_ff == 7'h25; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6603 = _T_6601 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6604 = _T_6600 | _T_6603; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6605 = _T_6604 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6607 = _T_6605 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6617 = _T_4987 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6618 = perr_ic_index_ff == 7'h26; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6620 = _T_6618 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6621 = _T_6617 | _T_6620; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6622 = _T_6621 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6624 = _T_6622 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6634 = _T_4988 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6635 = perr_ic_index_ff == 7'h27; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6637 = _T_6635 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6638 = _T_6634 | _T_6637; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6639 = _T_6638 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6641 = _T_6639 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6651 = _T_4989 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6652 = perr_ic_index_ff == 7'h28; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6654 = _T_6652 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6655 = _T_6651 | _T_6654; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6656 = _T_6655 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6658 = _T_6656 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6668 = _T_4990 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6669 = perr_ic_index_ff == 7'h29; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6671 = _T_6669 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6672 = _T_6668 | _T_6671; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6673 = _T_6672 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6675 = _T_6673 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6685 = _T_4991 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6686 = perr_ic_index_ff == 7'h2a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6688 = _T_6686 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6689 = _T_6685 | _T_6688; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6690 = _T_6689 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6692 = _T_6690 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6702 = _T_4992 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6703 = perr_ic_index_ff == 7'h2b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6705 = _T_6703 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6706 = _T_6702 | _T_6705; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6707 = _T_6706 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6709 = _T_6707 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6719 = _T_4993 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6720 = perr_ic_index_ff == 7'h2c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6722 = _T_6720 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6723 = _T_6719 | _T_6722; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6724 = _T_6723 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6726 = _T_6724 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6736 = _T_4994 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6737 = perr_ic_index_ff == 7'h2d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6739 = _T_6737 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6740 = _T_6736 | _T_6739; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6741 = _T_6740 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6743 = _T_6741 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6753 = _T_4995 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6754 = perr_ic_index_ff == 7'h2e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6756 = _T_6754 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6757 = _T_6753 | _T_6756; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6758 = _T_6757 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6760 = _T_6758 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6770 = _T_4996 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6771 = perr_ic_index_ff == 7'h2f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6773 = _T_6771 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6774 = _T_6770 | _T_6773; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6775 = _T_6774 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6777 = _T_6775 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6787 = _T_4997 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6788 = perr_ic_index_ff == 7'h30; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6790 = _T_6788 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6791 = _T_6787 | _T_6790; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6792 = _T_6791 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6794 = _T_6792 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6804 = _T_4998 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6805 = perr_ic_index_ff == 7'h31; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6807 = _T_6805 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6808 = _T_6804 | _T_6807; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6809 = _T_6808 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6811 = _T_6809 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6821 = _T_4999 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6822 = perr_ic_index_ff == 7'h32; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6824 = _T_6822 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6825 = _T_6821 | _T_6824; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6826 = _T_6825 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6828 = _T_6826 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6838 = _T_5000 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6839 = perr_ic_index_ff == 7'h33; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6841 = _T_6839 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6842 = _T_6838 | _T_6841; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6843 = _T_6842 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6845 = _T_6843 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6855 = _T_5001 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6856 = perr_ic_index_ff == 7'h34; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6858 = _T_6856 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6859 = _T_6855 | _T_6858; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6860 = _T_6859 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6862 = _T_6860 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6872 = _T_5002 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6873 = perr_ic_index_ff == 7'h35; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6875 = _T_6873 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6876 = _T_6872 | _T_6875; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6877 = _T_6876 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6879 = _T_6877 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6889 = _T_5003 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6890 = perr_ic_index_ff == 7'h36; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6892 = _T_6890 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6893 = _T_6889 | _T_6892; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6894 = _T_6893 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6896 = _T_6894 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6906 = _T_5004 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6907 = perr_ic_index_ff == 7'h37; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6909 = _T_6907 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6910 = _T_6906 | _T_6909; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6911 = _T_6910 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6913 = _T_6911 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6923 = _T_5005 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6924 = perr_ic_index_ff == 7'h38; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6926 = _T_6924 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6927 = _T_6923 | _T_6926; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6928 = _T_6927 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6930 = _T_6928 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6940 = _T_5006 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6941 = perr_ic_index_ff == 7'h39; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6943 = _T_6941 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6944 = _T_6940 | _T_6943; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6945 = _T_6944 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6947 = _T_6945 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6957 = _T_5007 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6958 = perr_ic_index_ff == 7'h3a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6960 = _T_6958 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6961 = _T_6957 | _T_6960; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6962 = _T_6961 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6964 = _T_6962 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6974 = _T_5008 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6975 = perr_ic_index_ff == 7'h3b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6977 = _T_6975 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6978 = _T_6974 | _T_6977; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6979 = _T_6978 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6981 = _T_6979 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_6991 = _T_5009 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_6992 = perr_ic_index_ff == 7'h3c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_6994 = _T_6992 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_6995 = _T_6991 | _T_6994; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_6996 = _T_6995 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_6998 = _T_6996 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7008 = _T_5010 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7009 = perr_ic_index_ff == 7'h3d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7011 = _T_7009 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7012 = _T_7008 | _T_7011; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7013 = _T_7012 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7015 = _T_7013 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7025 = _T_5011 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7026 = perr_ic_index_ff == 7'h3e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7028 = _T_7026 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7029 = _T_7025 | _T_7028; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7030 = _T_7029 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7032 = _T_7030 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7042 = _T_5012 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7043 = perr_ic_index_ff == 7'h3f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7045 = _T_7043 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7046 = _T_7042 | _T_7045; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7047 = _T_7046 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7049 = _T_7047 & tag_valid_clken_1[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7059 = _T_4981 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7062 = _T_6516 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7063 = _T_7059 | _T_7062; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7064 = _T_7063 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7066 = _T_7064 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7076 = _T_4982 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7079 = _T_6533 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7080 = _T_7076 | _T_7079; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7081 = _T_7080 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7083 = _T_7081 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7093 = _T_4983 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7096 = _T_6550 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7097 = _T_7093 | _T_7096; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7098 = _T_7097 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7100 = _T_7098 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7110 = _T_4984 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7113 = _T_6567 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7114 = _T_7110 | _T_7113; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7115 = _T_7114 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7117 = _T_7115 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7127 = _T_4985 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7130 = _T_6584 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7131 = _T_7127 | _T_7130; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7132 = _T_7131 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7134 = _T_7132 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7144 = _T_4986 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7147 = _T_6601 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7148 = _T_7144 | _T_7147; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7149 = _T_7148 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7151 = _T_7149 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7161 = _T_4987 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7164 = _T_6618 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7165 = _T_7161 | _T_7164; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7166 = _T_7165 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7168 = _T_7166 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7178 = _T_4988 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7181 = _T_6635 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7182 = _T_7178 | _T_7181; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7183 = _T_7182 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7185 = _T_7183 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7195 = _T_4989 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7198 = _T_6652 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7199 = _T_7195 | _T_7198; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7200 = _T_7199 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7202 = _T_7200 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7212 = _T_4990 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7215 = _T_6669 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7216 = _T_7212 | _T_7215; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7217 = _T_7216 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7219 = _T_7217 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7229 = _T_4991 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7232 = _T_6686 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7233 = _T_7229 | _T_7232; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7234 = _T_7233 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7236 = _T_7234 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7246 = _T_4992 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7249 = _T_6703 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7250 = _T_7246 | _T_7249; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7251 = _T_7250 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7253 = _T_7251 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7263 = _T_4993 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7266 = _T_6720 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7267 = _T_7263 | _T_7266; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7268 = _T_7267 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7270 = _T_7268 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7280 = _T_4994 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7283 = _T_6737 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7284 = _T_7280 | _T_7283; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7285 = _T_7284 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7287 = _T_7285 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7297 = _T_4995 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7300 = _T_6754 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7301 = _T_7297 | _T_7300; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7302 = _T_7301 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7304 = _T_7302 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7314 = _T_4996 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7317 = _T_6771 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7318 = _T_7314 | _T_7317; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7319 = _T_7318 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7321 = _T_7319 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7331 = _T_4997 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7334 = _T_6788 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7335 = _T_7331 | _T_7334; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7336 = _T_7335 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7338 = _T_7336 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7348 = _T_4998 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7351 = _T_6805 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7352 = _T_7348 | _T_7351; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7353 = _T_7352 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7355 = _T_7353 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7365 = _T_4999 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7368 = _T_6822 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7369 = _T_7365 | _T_7368; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7370 = _T_7369 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7372 = _T_7370 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7382 = _T_5000 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7385 = _T_6839 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7386 = _T_7382 | _T_7385; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7387 = _T_7386 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7389 = _T_7387 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7399 = _T_5001 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7402 = _T_6856 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7403 = _T_7399 | _T_7402; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7404 = _T_7403 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7406 = _T_7404 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7416 = _T_5002 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7419 = _T_6873 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7420 = _T_7416 | _T_7419; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7421 = _T_7420 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7423 = _T_7421 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7433 = _T_5003 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7436 = _T_6890 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7437 = _T_7433 | _T_7436; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7438 = _T_7437 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7440 = _T_7438 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7450 = _T_5004 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7453 = _T_6907 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7454 = _T_7450 | _T_7453; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7455 = _T_7454 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7457 = _T_7455 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7467 = _T_5005 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7470 = _T_6924 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7471 = _T_7467 | _T_7470; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7472 = _T_7471 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7474 = _T_7472 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7484 = _T_5006 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7487 = _T_6941 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7488 = _T_7484 | _T_7487; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7489 = _T_7488 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7491 = _T_7489 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7501 = _T_5007 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7504 = _T_6958 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7505 = _T_7501 | _T_7504; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7506 = _T_7505 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7508 = _T_7506 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7518 = _T_5008 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7521 = _T_6975 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7522 = _T_7518 | _T_7521; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7523 = _T_7522 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7525 = _T_7523 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7535 = _T_5009 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7538 = _T_6992 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7539 = _T_7535 | _T_7538; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7540 = _T_7539 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7542 = _T_7540 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7552 = _T_5010 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7555 = _T_7009 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7556 = _T_7552 | _T_7555; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7557 = _T_7556 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7559 = _T_7557 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7569 = _T_5011 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7572 = _T_7026 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7573 = _T_7569 | _T_7572; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7574 = _T_7573 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7576 = _T_7574 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7586 = _T_5012 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7589 = _T_7043 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7590 = _T_7586 | _T_7589; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7591 = _T_7590 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7593 = _T_7591 & tag_valid_clken_1[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7603 = _T_5013 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7604 = perr_ic_index_ff == 7'h40; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7606 = _T_7604 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7607 = _T_7603 | _T_7606; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7608 = _T_7607 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7610 = _T_7608 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7620 = _T_5014 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7621 = perr_ic_index_ff == 7'h41; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7623 = _T_7621 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7624 = _T_7620 | _T_7623; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7625 = _T_7624 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7627 = _T_7625 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7637 = _T_5015 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7638 = perr_ic_index_ff == 7'h42; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7640 = _T_7638 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7641 = _T_7637 | _T_7640; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7642 = _T_7641 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7644 = _T_7642 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7654 = _T_5016 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7655 = perr_ic_index_ff == 7'h43; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7657 = _T_7655 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7658 = _T_7654 | _T_7657; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7659 = _T_7658 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7661 = _T_7659 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7671 = _T_5017 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7672 = perr_ic_index_ff == 7'h44; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7674 = _T_7672 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7675 = _T_7671 | _T_7674; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7676 = _T_7675 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7678 = _T_7676 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7688 = _T_5018 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7689 = perr_ic_index_ff == 7'h45; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7691 = _T_7689 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7692 = _T_7688 | _T_7691; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7693 = _T_7692 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7695 = _T_7693 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7705 = _T_5019 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7706 = perr_ic_index_ff == 7'h46; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7708 = _T_7706 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7709 = _T_7705 | _T_7708; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7710 = _T_7709 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7712 = _T_7710 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7722 = _T_5020 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7723 = perr_ic_index_ff == 7'h47; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7725 = _T_7723 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7726 = _T_7722 | _T_7725; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7727 = _T_7726 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7729 = _T_7727 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7739 = _T_5021 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7740 = perr_ic_index_ff == 7'h48; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7742 = _T_7740 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7743 = _T_7739 | _T_7742; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7744 = _T_7743 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7746 = _T_7744 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7756 = _T_5022 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7757 = perr_ic_index_ff == 7'h49; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7759 = _T_7757 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7760 = _T_7756 | _T_7759; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7761 = _T_7760 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7763 = _T_7761 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7773 = _T_5023 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7774 = perr_ic_index_ff == 7'h4a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7776 = _T_7774 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7777 = _T_7773 | _T_7776; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7778 = _T_7777 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7780 = _T_7778 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7790 = _T_5024 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7791 = perr_ic_index_ff == 7'h4b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7793 = _T_7791 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7794 = _T_7790 | _T_7793; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7795 = _T_7794 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7797 = _T_7795 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7807 = _T_5025 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7808 = perr_ic_index_ff == 7'h4c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7810 = _T_7808 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7811 = _T_7807 | _T_7810; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7812 = _T_7811 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7814 = _T_7812 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7824 = _T_5026 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7825 = perr_ic_index_ff == 7'h4d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7827 = _T_7825 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7828 = _T_7824 | _T_7827; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7829 = _T_7828 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7831 = _T_7829 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7841 = _T_5027 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7842 = perr_ic_index_ff == 7'h4e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7844 = _T_7842 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7845 = _T_7841 | _T_7844; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7846 = _T_7845 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7848 = _T_7846 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7858 = _T_5028 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7859 = perr_ic_index_ff == 7'h4f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7861 = _T_7859 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7862 = _T_7858 | _T_7861; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7863 = _T_7862 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7865 = _T_7863 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7875 = _T_5029 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7876 = perr_ic_index_ff == 7'h50; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7878 = _T_7876 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7879 = _T_7875 | _T_7878; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7880 = _T_7879 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7882 = _T_7880 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7892 = _T_5030 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7893 = perr_ic_index_ff == 7'h51; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7895 = _T_7893 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7896 = _T_7892 | _T_7895; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7897 = _T_7896 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7899 = _T_7897 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7909 = _T_5031 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7910 = perr_ic_index_ff == 7'h52; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7912 = _T_7910 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7913 = _T_7909 | _T_7912; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7914 = _T_7913 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7916 = _T_7914 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7926 = _T_5032 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7927 = perr_ic_index_ff == 7'h53; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7929 = _T_7927 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7930 = _T_7926 | _T_7929; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7931 = _T_7930 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7933 = _T_7931 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7943 = _T_5033 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7944 = perr_ic_index_ff == 7'h54; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7946 = _T_7944 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7947 = _T_7943 | _T_7946; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7948 = _T_7947 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7950 = _T_7948 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7960 = _T_5034 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7961 = perr_ic_index_ff == 7'h55; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7963 = _T_7961 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7964 = _T_7960 | _T_7963; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7965 = _T_7964 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7967 = _T_7965 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7977 = _T_5035 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7978 = perr_ic_index_ff == 7'h56; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7980 = _T_7978 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7981 = _T_7977 | _T_7980; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7982 = _T_7981 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_7984 = _T_7982 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_7994 = _T_5036 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_7995 = perr_ic_index_ff == 7'h57; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_7997 = _T_7995 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_7998 = _T_7994 | _T_7997; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_7999 = _T_7998 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8001 = _T_7999 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8011 = _T_5037 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8012 = perr_ic_index_ff == 7'h58; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8014 = _T_8012 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8015 = _T_8011 | _T_8014; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8016 = _T_8015 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8018 = _T_8016 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8028 = _T_5038 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8029 = perr_ic_index_ff == 7'h59; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8031 = _T_8029 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8032 = _T_8028 | _T_8031; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8033 = _T_8032 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8035 = _T_8033 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8045 = _T_5039 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8046 = perr_ic_index_ff == 7'h5a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8048 = _T_8046 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8049 = _T_8045 | _T_8048; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8050 = _T_8049 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8052 = _T_8050 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8062 = _T_5040 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8063 = perr_ic_index_ff == 7'h5b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8065 = _T_8063 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8066 = _T_8062 | _T_8065; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8067 = _T_8066 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8069 = _T_8067 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8079 = _T_5041 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8080 = perr_ic_index_ff == 7'h5c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8082 = _T_8080 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8083 = _T_8079 | _T_8082; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8084 = _T_8083 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8086 = _T_8084 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8096 = _T_5042 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8097 = perr_ic_index_ff == 7'h5d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8099 = _T_8097 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8100 = _T_8096 | _T_8099; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8101 = _T_8100 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8103 = _T_8101 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8113 = _T_5043 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8114 = perr_ic_index_ff == 7'h5e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8116 = _T_8114 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8117 = _T_8113 | _T_8116; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8118 = _T_8117 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8120 = _T_8118 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8130 = _T_5044 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8131 = perr_ic_index_ff == 7'h5f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8133 = _T_8131 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8134 = _T_8130 | _T_8133; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8135 = _T_8134 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8137 = _T_8135 & tag_valid_clken_2[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8147 = _T_5013 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8150 = _T_7604 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8151 = _T_8147 | _T_8150; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8152 = _T_8151 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8154 = _T_8152 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8164 = _T_5014 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8167 = _T_7621 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8168 = _T_8164 | _T_8167; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8169 = _T_8168 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8171 = _T_8169 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8181 = _T_5015 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8184 = _T_7638 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8185 = _T_8181 | _T_8184; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8186 = _T_8185 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8188 = _T_8186 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8198 = _T_5016 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8201 = _T_7655 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8202 = _T_8198 | _T_8201; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8203 = _T_8202 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8205 = _T_8203 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8215 = _T_5017 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8218 = _T_7672 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8219 = _T_8215 | _T_8218; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8220 = _T_8219 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8222 = _T_8220 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8232 = _T_5018 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8235 = _T_7689 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8236 = _T_8232 | _T_8235; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8237 = _T_8236 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8239 = _T_8237 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8249 = _T_5019 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8252 = _T_7706 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8253 = _T_8249 | _T_8252; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8254 = _T_8253 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8256 = _T_8254 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8266 = _T_5020 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8269 = _T_7723 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8270 = _T_8266 | _T_8269; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8271 = _T_8270 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8273 = _T_8271 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8283 = _T_5021 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8286 = _T_7740 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8287 = _T_8283 | _T_8286; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8288 = _T_8287 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8290 = _T_8288 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8300 = _T_5022 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8303 = _T_7757 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8304 = _T_8300 | _T_8303; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8305 = _T_8304 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8307 = _T_8305 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8317 = _T_5023 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8320 = _T_7774 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8321 = _T_8317 | _T_8320; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8322 = _T_8321 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8324 = _T_8322 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8334 = _T_5024 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8337 = _T_7791 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8338 = _T_8334 | _T_8337; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8339 = _T_8338 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8341 = _T_8339 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8351 = _T_5025 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8354 = _T_7808 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8355 = _T_8351 | _T_8354; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8356 = _T_8355 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8358 = _T_8356 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8368 = _T_5026 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8371 = _T_7825 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8372 = _T_8368 | _T_8371; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8373 = _T_8372 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8375 = _T_8373 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8385 = _T_5027 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8388 = _T_7842 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8389 = _T_8385 | _T_8388; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8390 = _T_8389 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8392 = _T_8390 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8402 = _T_5028 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8405 = _T_7859 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8406 = _T_8402 | _T_8405; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8407 = _T_8406 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8409 = _T_8407 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8419 = _T_5029 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8422 = _T_7876 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8423 = _T_8419 | _T_8422; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8424 = _T_8423 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8426 = _T_8424 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8436 = _T_5030 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8439 = _T_7893 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8440 = _T_8436 | _T_8439; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8441 = _T_8440 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8443 = _T_8441 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8453 = _T_5031 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8456 = _T_7910 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8457 = _T_8453 | _T_8456; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8458 = _T_8457 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8460 = _T_8458 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8470 = _T_5032 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8473 = _T_7927 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8474 = _T_8470 | _T_8473; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8475 = _T_8474 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8477 = _T_8475 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8487 = _T_5033 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8490 = _T_7944 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8491 = _T_8487 | _T_8490; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8492 = _T_8491 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8494 = _T_8492 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8504 = _T_5034 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8507 = _T_7961 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8508 = _T_8504 | _T_8507; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8509 = _T_8508 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8511 = _T_8509 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8521 = _T_5035 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8524 = _T_7978 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8525 = _T_8521 | _T_8524; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8526 = _T_8525 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8528 = _T_8526 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8538 = _T_5036 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8541 = _T_7995 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8542 = _T_8538 | _T_8541; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8543 = _T_8542 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8545 = _T_8543 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8555 = _T_5037 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8558 = _T_8012 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8559 = _T_8555 | _T_8558; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8560 = _T_8559 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8562 = _T_8560 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8572 = _T_5038 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8575 = _T_8029 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8576 = _T_8572 | _T_8575; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8577 = _T_8576 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8579 = _T_8577 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8589 = _T_5039 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8592 = _T_8046 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8593 = _T_8589 | _T_8592; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8594 = _T_8593 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8596 = _T_8594 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8606 = _T_5040 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8609 = _T_8063 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8610 = _T_8606 | _T_8609; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8611 = _T_8610 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8613 = _T_8611 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8623 = _T_5041 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8626 = _T_8080 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8627 = _T_8623 | _T_8626; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8628 = _T_8627 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8630 = _T_8628 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8640 = _T_5042 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8643 = _T_8097 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8644 = _T_8640 | _T_8643; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8645 = _T_8644 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8647 = _T_8645 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8657 = _T_5043 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8660 = _T_8114 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8661 = _T_8657 | _T_8660; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8662 = _T_8661 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8664 = _T_8662 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8674 = _T_5044 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8677 = _T_8131 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8678 = _T_8674 | _T_8677; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8679 = _T_8678 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8681 = _T_8679 & tag_valid_clken_2[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8691 = _T_5045 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8692 = perr_ic_index_ff == 7'h60; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8694 = _T_8692 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8695 = _T_8691 | _T_8694; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8696 = _T_8695 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8698 = _T_8696 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8708 = _T_5046 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8709 = perr_ic_index_ff == 7'h61; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8711 = _T_8709 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8712 = _T_8708 | _T_8711; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8713 = _T_8712 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8715 = _T_8713 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8725 = _T_5047 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8726 = perr_ic_index_ff == 7'h62; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8728 = _T_8726 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8729 = _T_8725 | _T_8728; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8730 = _T_8729 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8732 = _T_8730 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8742 = _T_5048 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8743 = perr_ic_index_ff == 7'h63; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8745 = _T_8743 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8746 = _T_8742 | _T_8745; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8747 = _T_8746 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8749 = _T_8747 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8759 = _T_5049 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8760 = perr_ic_index_ff == 7'h64; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8762 = _T_8760 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8763 = _T_8759 | _T_8762; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8764 = _T_8763 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8766 = _T_8764 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8776 = _T_5050 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8777 = perr_ic_index_ff == 7'h65; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8779 = _T_8777 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8780 = _T_8776 | _T_8779; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8781 = _T_8780 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8783 = _T_8781 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8793 = _T_5051 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8794 = perr_ic_index_ff == 7'h66; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8796 = _T_8794 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8797 = _T_8793 | _T_8796; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8798 = _T_8797 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8800 = _T_8798 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8810 = _T_5052 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8811 = perr_ic_index_ff == 7'h67; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8813 = _T_8811 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8814 = _T_8810 | _T_8813; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8815 = _T_8814 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8817 = _T_8815 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8827 = _T_5053 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8828 = perr_ic_index_ff == 7'h68; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8830 = _T_8828 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8831 = _T_8827 | _T_8830; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8832 = _T_8831 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8834 = _T_8832 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8844 = _T_5054 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8845 = perr_ic_index_ff == 7'h69; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8847 = _T_8845 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8848 = _T_8844 | _T_8847; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8849 = _T_8848 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8851 = _T_8849 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8861 = _T_5055 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8862 = perr_ic_index_ff == 7'h6a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8864 = _T_8862 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8865 = _T_8861 | _T_8864; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8866 = _T_8865 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8868 = _T_8866 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8878 = _T_5056 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8879 = perr_ic_index_ff == 7'h6b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8881 = _T_8879 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8882 = _T_8878 | _T_8881; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8883 = _T_8882 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8885 = _T_8883 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8895 = _T_5057 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8896 = perr_ic_index_ff == 7'h6c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8898 = _T_8896 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8899 = _T_8895 | _T_8898; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8900 = _T_8899 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8902 = _T_8900 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8912 = _T_5058 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8913 = perr_ic_index_ff == 7'h6d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8915 = _T_8913 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8916 = _T_8912 | _T_8915; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8917 = _T_8916 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8919 = _T_8917 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8929 = _T_5059 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8930 = perr_ic_index_ff == 7'h6e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8932 = _T_8930 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8933 = _T_8929 | _T_8932; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8934 = _T_8933 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8936 = _T_8934 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8946 = _T_5060 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8947 = perr_ic_index_ff == 7'h6f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8949 = _T_8947 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8950 = _T_8946 | _T_8949; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8951 = _T_8950 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8953 = _T_8951 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8963 = _T_5061 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8964 = perr_ic_index_ff == 7'h70; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8966 = _T_8964 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8967 = _T_8963 | _T_8966; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8968 = _T_8967 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8970 = _T_8968 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8980 = _T_5062 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8981 = perr_ic_index_ff == 7'h71; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_8983 = _T_8981 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_8984 = _T_8980 | _T_8983; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_8985 = _T_8984 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_8987 = _T_8985 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_8997 = _T_5063 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_8998 = perr_ic_index_ff == 7'h72; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9000 = _T_8998 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9001 = _T_8997 | _T_9000; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9002 = _T_9001 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9004 = _T_9002 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9014 = _T_5064 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9015 = perr_ic_index_ff == 7'h73; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9017 = _T_9015 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9018 = _T_9014 | _T_9017; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9019 = _T_9018 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9021 = _T_9019 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9031 = _T_5065 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9032 = perr_ic_index_ff == 7'h74; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9034 = _T_9032 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9035 = _T_9031 | _T_9034; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9036 = _T_9035 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9038 = _T_9036 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9048 = _T_5066 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9049 = perr_ic_index_ff == 7'h75; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9051 = _T_9049 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9052 = _T_9048 | _T_9051; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9053 = _T_9052 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9055 = _T_9053 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9065 = _T_5067 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9066 = perr_ic_index_ff == 7'h76; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9068 = _T_9066 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9069 = _T_9065 | _T_9068; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9070 = _T_9069 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9072 = _T_9070 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9082 = _T_5068 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9083 = perr_ic_index_ff == 7'h77; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9085 = _T_9083 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9086 = _T_9082 | _T_9085; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9087 = _T_9086 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9089 = _T_9087 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9099 = _T_5069 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9100 = perr_ic_index_ff == 7'h78; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9102 = _T_9100 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9103 = _T_9099 | _T_9102; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9104 = _T_9103 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9106 = _T_9104 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9116 = _T_5070 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9117 = perr_ic_index_ff == 7'h79; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9119 = _T_9117 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9120 = _T_9116 | _T_9119; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9121 = _T_9120 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9123 = _T_9121 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9133 = _T_5071 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9134 = perr_ic_index_ff == 7'h7a; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9136 = _T_9134 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9137 = _T_9133 | _T_9136; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9138 = _T_9137 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9140 = _T_9138 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9150 = _T_5072 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9151 = perr_ic_index_ff == 7'h7b; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9153 = _T_9151 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9154 = _T_9150 | _T_9153; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9155 = _T_9154 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9157 = _T_9155 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9167 = _T_5073 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9168 = perr_ic_index_ff == 7'h7c; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9170 = _T_9168 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9171 = _T_9167 | _T_9170; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9172 = _T_9171 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9174 = _T_9172 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9184 = _T_5074 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9185 = perr_ic_index_ff == 7'h7d; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9187 = _T_9185 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9188 = _T_9184 | _T_9187; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9189 = _T_9188 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9191 = _T_9189 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9201 = _T_5075 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9202 = perr_ic_index_ff == 7'h7e; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9204 = _T_9202 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9205 = _T_9201 | _T_9204; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9206 = _T_9205 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9208 = _T_9206 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9218 = _T_5076 & ifu_tag_wren_ff[0]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9219 = perr_ic_index_ff == 7'h7f; // @[el2_ifu_mem_ctl.scala 758:102]
  wire  _T_9221 = _T_9219 & perr_err_inv_way[0]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9222 = _T_9218 | _T_9221; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9223 = _T_9222 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9225 = _T_9223 & tag_valid_clken_3[0]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9235 = _T_5045 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9238 = _T_8692 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9239 = _T_9235 | _T_9238; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9240 = _T_9239 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9242 = _T_9240 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9252 = _T_5046 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9255 = _T_8709 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9256 = _T_9252 | _T_9255; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9257 = _T_9256 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9259 = _T_9257 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9269 = _T_5047 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9272 = _T_8726 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9273 = _T_9269 | _T_9272; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9274 = _T_9273 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9276 = _T_9274 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9286 = _T_5048 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9289 = _T_8743 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9290 = _T_9286 | _T_9289; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9291 = _T_9290 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9293 = _T_9291 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9303 = _T_5049 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9306 = _T_8760 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9307 = _T_9303 | _T_9306; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9308 = _T_9307 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9310 = _T_9308 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9320 = _T_5050 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9323 = _T_8777 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9324 = _T_9320 | _T_9323; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9325 = _T_9324 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9327 = _T_9325 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9337 = _T_5051 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9340 = _T_8794 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9341 = _T_9337 | _T_9340; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9342 = _T_9341 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9344 = _T_9342 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9354 = _T_5052 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9357 = _T_8811 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9358 = _T_9354 | _T_9357; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9359 = _T_9358 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9361 = _T_9359 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9371 = _T_5053 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9374 = _T_8828 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9375 = _T_9371 | _T_9374; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9376 = _T_9375 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9378 = _T_9376 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9388 = _T_5054 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9391 = _T_8845 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9392 = _T_9388 | _T_9391; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9393 = _T_9392 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9395 = _T_9393 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9405 = _T_5055 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9408 = _T_8862 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9409 = _T_9405 | _T_9408; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9410 = _T_9409 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9412 = _T_9410 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9422 = _T_5056 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9425 = _T_8879 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9426 = _T_9422 | _T_9425; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9427 = _T_9426 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9429 = _T_9427 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9439 = _T_5057 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9442 = _T_8896 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9443 = _T_9439 | _T_9442; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9444 = _T_9443 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9446 = _T_9444 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9456 = _T_5058 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9459 = _T_8913 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9460 = _T_9456 | _T_9459; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9461 = _T_9460 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9463 = _T_9461 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9473 = _T_5059 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9476 = _T_8930 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9477 = _T_9473 | _T_9476; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9478 = _T_9477 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9480 = _T_9478 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9490 = _T_5060 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9493 = _T_8947 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9494 = _T_9490 | _T_9493; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9495 = _T_9494 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9497 = _T_9495 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9507 = _T_5061 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9510 = _T_8964 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9511 = _T_9507 | _T_9510; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9512 = _T_9511 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9514 = _T_9512 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9524 = _T_5062 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9527 = _T_8981 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9528 = _T_9524 | _T_9527; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9529 = _T_9528 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9531 = _T_9529 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9541 = _T_5063 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9544 = _T_8998 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9545 = _T_9541 | _T_9544; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9546 = _T_9545 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9548 = _T_9546 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9558 = _T_5064 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9561 = _T_9015 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9562 = _T_9558 | _T_9561; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9563 = _T_9562 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9565 = _T_9563 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9575 = _T_5065 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9578 = _T_9032 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9579 = _T_9575 | _T_9578; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9580 = _T_9579 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9582 = _T_9580 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9592 = _T_5066 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9595 = _T_9049 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9596 = _T_9592 | _T_9595; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9597 = _T_9596 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9599 = _T_9597 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9609 = _T_5067 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9612 = _T_9066 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9613 = _T_9609 | _T_9612; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9614 = _T_9613 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9616 = _T_9614 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9626 = _T_5068 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9629 = _T_9083 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9630 = _T_9626 | _T_9629; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9631 = _T_9630 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9633 = _T_9631 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9643 = _T_5069 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9646 = _T_9100 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9647 = _T_9643 | _T_9646; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9648 = _T_9647 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9650 = _T_9648 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9660 = _T_5070 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9663 = _T_9117 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9664 = _T_9660 | _T_9663; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9665 = _T_9664 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9667 = _T_9665 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9677 = _T_5071 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9680 = _T_9134 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9681 = _T_9677 | _T_9680; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9682 = _T_9681 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9684 = _T_9682 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9694 = _T_5072 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9697 = _T_9151 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9698 = _T_9694 | _T_9697; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9699 = _T_9698 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9701 = _T_9699 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9711 = _T_5073 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9714 = _T_9168 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9715 = _T_9711 | _T_9714; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9716 = _T_9715 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9718 = _T_9716 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9728 = _T_5074 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9731 = _T_9185 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9732 = _T_9728 | _T_9731; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9733 = _T_9732 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9735 = _T_9733 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9745 = _T_5075 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9748 = _T_9202 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9749 = _T_9745 | _T_9748; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9750 = _T_9749 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9752 = _T_9750 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_9762 = _T_5076 & ifu_tag_wren_ff[1]; // @[el2_ifu_mem_ctl.scala 758:59]
  wire  _T_9765 = _T_9219 & perr_err_inv_way[1]; // @[el2_ifu_mem_ctl.scala 758:124]
  wire  _T_9766 = _T_9762 | _T_9765; // @[el2_ifu_mem_ctl.scala 758:81]
  wire  _T_9767 = _T_9766 | reset_all_tags; // @[el2_ifu_mem_ctl.scala 758:147]
  wire  _T_9769 = _T_9767 & tag_valid_clken_3[1]; // @[el2_ifu_mem_ctl.scala 758:165]
  wire  _T_10571 = ~fetch_uncacheable_ff; // @[el2_ifu_mem_ctl.scala 813:63]
  wire  _T_10572 = _T_10571 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 813:85]
  wire [1:0] _T_10574 = _T_10572 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  _T_10581; // @[el2_ifu_mem_ctl.scala 818:57]
  reg  _T_10582; // @[el2_ifu_mem_ctl.scala 819:56]
  reg  _T_10583; // @[el2_ifu_mem_ctl.scala 820:59]
  wire  _T_10584 = ~ifu_bus_arready_ff; // @[el2_ifu_mem_ctl.scala 821:80]
  wire  _T_10585 = ifu_bus_arvalid_ff & _T_10584; // @[el2_ifu_mem_ctl.scala 821:78]
  wire  _T_10586 = _T_10585 & miss_pending; // @[el2_ifu_mem_ctl.scala 821:100]
  reg  _T_10587; // @[el2_ifu_mem_ctl.scala 821:58]
  reg  _T_10588; // @[el2_ifu_mem_ctl.scala 822:58]
  wire  _T_10591 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h3; // @[el2_ifu_mem_ctl.scala 829:71]
  wire  _T_10593 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h2; // @[el2_ifu_mem_ctl.scala 829:124]
  wire  _T_10595 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h1; // @[el2_ifu_mem_ctl.scala 830:50]
  wire  _T_10597 = io_dec_tlu_ic_diag_pkt_icache_dicawics[15:14] == 2'h0; // @[el2_ifu_mem_ctl.scala 830:103]
  wire [3:0] _T_10600 = {_T_10591,_T_10593,_T_10595,_T_10597}; // @[Cat.scala 29:58]
  wire  ic_debug_ict_array_sel_in = io_ic_debug_rd_en & io_ic_debug_tag_array; // @[el2_ifu_mem_ctl.scala 832:53]
  reg  _T_10611; // @[Reg.scala 27:20]
  assign io_ifu_miss_state_idle = miss_state == 3'h0; // @[el2_ifu_mem_ctl.scala 328:26]
  assign io_ifu_ic_mb_empty = _T_326 | _T_231; // @[el2_ifu_mem_ctl.scala 327:22]
  assign io_ic_dma_active = _T_11 | io_dec_tlu_flush_err_wb; // @[el2_ifu_mem_ctl.scala 192:20]
  assign io_ic_write_stall = write_ic_16_bytes & _T_4138; // @[el2_ifu_mem_ctl.scala 699:21]
  assign io_ifu_pmu_ic_miss = _T_10581; // @[el2_ifu_mem_ctl.scala 818:22]
  assign io_ifu_pmu_ic_hit = _T_10582; // @[el2_ifu_mem_ctl.scala 819:21]
  assign io_ifu_pmu_bus_error = _T_10583; // @[el2_ifu_mem_ctl.scala 820:24]
  assign io_ifu_pmu_bus_busy = _T_10587; // @[el2_ifu_mem_ctl.scala 821:23]
  assign io_ifu_pmu_bus_trxn = _T_10588; // @[el2_ifu_mem_ctl.scala 822:23]
  assign io_ifu_axi_awvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 142:22]
  assign io_ifu_axi_awid = 3'h0; // @[el2_ifu_mem_ctl.scala 141:19]
  assign io_ifu_axi_awaddr = 32'h0; // @[el2_ifu_mem_ctl.scala 136:21]
  assign io_ifu_axi_awregion = 4'h0; // @[el2_ifu_mem_ctl.scala 140:23]
  assign io_ifu_axi_awlen = 8'h0; // @[el2_ifu_mem_ctl.scala 138:20]
  assign io_ifu_axi_awsize = 3'h0; // @[el2_ifu_mem_ctl.scala 149:21]
  assign io_ifu_axi_awburst = 2'h0; // @[el2_ifu_mem_ctl.scala 151:22]
  assign io_ifu_axi_awlock = 1'h0; // @[el2_ifu_mem_ctl.scala 146:21]
  assign io_ifu_axi_awcache = 4'h0; // @[el2_ifu_mem_ctl.scala 144:22]
  assign io_ifu_axi_awprot = 3'h0; // @[el2_ifu_mem_ctl.scala 137:21]
  assign io_ifu_axi_awqos = 4'h0; // @[el2_ifu_mem_ctl.scala 135:20]
  assign io_ifu_axi_wvalid = 1'h0; // @[el2_ifu_mem_ctl.scala 133:21]
  assign io_ifu_axi_wdata = 64'h0; // @[el2_ifu_mem_ctl.scala 134:20]
  assign io_ifu_axi_wstrb = 8'h0; // @[el2_ifu_mem_ctl.scala 143:20]
  assign io_ifu_axi_wlast = 1'h0; // @[el2_ifu_mem_ctl.scala 152:20]
  assign io_ifu_axi_bready = 1'h0; // @[el2_ifu_mem_ctl.scala 147:21]
  assign io_ifu_axi_arvalid = ifu_bus_cmd_valid; // @[el2_ifu_mem_ctl.scala 560:22]
  assign io_ifu_axi_arid = bus_rd_addr_count & _T_2572; // @[el2_ifu_mem_ctl.scala 561:19]
  assign io_ifu_axi_araddr = _T_2574 & _T_2576; // @[el2_ifu_mem_ctl.scala 562:21]
  assign io_ifu_axi_arregion = ifu_ic_req_addr_f[28:25]; // @[el2_ifu_mem_ctl.scala 565:23]
  assign io_ifu_axi_arlen = 8'h0; // @[el2_ifu_mem_ctl.scala 148:20]
  assign io_ifu_axi_arsize = 3'h3; // @[el2_ifu_mem_ctl.scala 563:21]
  assign io_ifu_axi_arburst = 2'h1; // @[el2_ifu_mem_ctl.scala 566:22]
  assign io_ifu_axi_arlock = 1'h0; // @[el2_ifu_mem_ctl.scala 139:21]
  assign io_ifu_axi_arcache = 4'hf; // @[el2_ifu_mem_ctl.scala 564:22]
  assign io_ifu_axi_arprot = 3'h0; // @[el2_ifu_mem_ctl.scala 150:21]
  assign io_ifu_axi_arqos = 4'h0; // @[el2_ifu_mem_ctl.scala 145:20]
  assign io_ifu_axi_rready = 1'h1; // @[el2_ifu_mem_ctl.scala 567:21]
  assign io_iccm_dma_ecc_error = |iccm_double_ecc_error; // @[el2_ifu_mem_ctl.scala 658:25]
  assign io_iccm_dma_rvalid = iccm_dma_rvalid_temp; // @[el2_ifu_mem_ctl.scala 656:22]
  assign io_iccm_dma_rdata = iccm_dma_rdata_temp; // @[el2_ifu_mem_ctl.scala 660:21]
  assign io_iccm_dma_rtag = iccm_dma_rtag_temp; // @[el2_ifu_mem_ctl.scala 651:20]
  assign io_iccm_ready = _T_2675 & _T_2669; // @[el2_ifu_mem_ctl.scala 630:17]
  assign io_ic_rw_addr = _T_338 | _T_339; // @[el2_ifu_mem_ctl.scala 337:17]
  assign io_ic_wr_en = bus_ic_wr_en & _T_4124; // @[el2_ifu_mem_ctl.scala 698:15]
  assign io_ic_rd_en = _T_4116 | _T_4121; // @[el2_ifu_mem_ctl.scala 689:15]
  assign io_ic_wr_data_0 = ic_wr_16bytes_data[70:0]; // @[el2_ifu_mem_ctl.scala 344:17]
  assign io_ic_wr_data_1 = ic_wr_16bytes_data[141:71]; // @[el2_ifu_mem_ctl.scala 344:17]
  assign io_ic_debug_wr_data = io_dec_tlu_ic_diag_pkt_icache_wrdata; // @[el2_ifu_mem_ctl.scala 345:23]
  assign io_ifu_ic_debug_rd_data = _T_1209; // @[el2_ifu_mem_ctl.scala 353:27]
  assign io_ic_debug_addr = io_dec_tlu_ic_diag_pkt_icache_dicawics[9:0]; // @[el2_ifu_mem_ctl.scala 825:20]
  assign io_ic_debug_rd_en = io_dec_tlu_ic_diag_pkt_icache_rd_valid; // @[el2_ifu_mem_ctl.scala 827:21]
  assign io_ic_debug_wr_en = io_dec_tlu_ic_diag_pkt_icache_wr_valid; // @[el2_ifu_mem_ctl.scala 828:21]
  assign io_ic_debug_tag_array = io_dec_tlu_ic_diag_pkt_icache_dicawics[16]; // @[el2_ifu_mem_ctl.scala 826:25]
  assign io_ic_debug_way = _T_10600[1:0]; // @[el2_ifu_mem_ctl.scala 829:19]
  assign io_ic_tag_valid = ic_tag_valid_unq & _T_10574; // @[el2_ifu_mem_ctl.scala 813:19]
  assign io_iccm_rw_addr = _T_3270[14:0]; // @[el2_ifu_mem_ctl.scala 662:19]
  assign io_iccm_wren = _T_2679 | iccm_correct_ecc; // @[el2_ifu_mem_ctl.scala 632:16]
  assign io_iccm_rden = _T_2683 | _T_2684; // @[el2_ifu_mem_ctl.scala 633:16]
  assign io_iccm_wr_data = _T_3245 ? _T_3246 : _T_3253; // @[el2_ifu_mem_ctl.scala 639:19]
  assign io_iccm_wr_size = _T_2689 & io_dma_mem_sz; // @[el2_ifu_mem_ctl.scala 635:19]
  assign io_ic_hit_f = _T_263 | _T_264; // @[el2_ifu_mem_ctl.scala 289:15]
  assign io_ic_access_fault_f = _T_2457 & _T_317; // @[el2_ifu_mem_ctl.scala 385:24]
  assign io_ic_access_fault_type_f = io_iccm_rd_ecc_double_err ? 2'h1 : _T_1271; // @[el2_ifu_mem_ctl.scala 386:29]
  assign io_iccm_rd_ecc_single_err = _T_4061 & ifc_fetch_req_f; // @[el2_ifu_mem_ctl.scala 675:29]
  assign io_iccm_rd_ecc_double_err = iccm_dma_ecc_error_in & ifc_iccm_access_f; // @[el2_ifu_mem_ctl.scala 676:29]
  assign io_ic_error_start = _T_1197 | ic_rd_parity_final_err; // @[el2_ifu_mem_ctl.scala 347:21]
  assign io_ifu_async_error_start = io_iccm_rd_ecc_single_err | io_ic_error_start; // @[el2_ifu_mem_ctl.scala 191:28]
  assign io_iccm_dma_sb_error = _T_3 & dma_iccm_req_f; // @[el2_ifu_mem_ctl.scala 190:24]
  assign io_ic_fetch_val_f = {_T_1279,fetch_req_f_qual}; // @[el2_ifu_mem_ctl.scala 389:21]
  assign io_ic_data_f = io_ic_rd_data[31:0]; // @[el2_ifu_mem_ctl.scala 382:16]
  assign io_ic_premux_data = ic_premux_data_temp[63:0]; // @[el2_ifu_mem_ctl.scala 379:21]
  assign io_ic_sel_premux_data = fetch_req_iccm_f | sel_byp_data; // @[el2_ifu_mem_ctl.scala 380:25]
  assign io_ifu_ic_debug_rd_data_valid = _T_10611; // @[el2_ifu_mem_ctl.scala 836:33]
  assign io_iccm_buf_correct_ecc = iccm_correct_ecc & _T_2462; // @[el2_ifu_mem_ctl.scala 479:27]
  assign io_iccm_correction_state = _T_2490 ? 1'h0 : _GEN_60; // @[el2_ifu_mem_ctl.scala 514:28 el2_ifu_mem_ctl.scala 527:32 el2_ifu_mem_ctl.scala 534:32 el2_ifu_mem_ctl.scala 541:32]
  assign io_test = {_T_2873,_T_2870}; // @[el2_ifu_mem_ctl.scala 636:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flush_final_f = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ifc_fetch_req_f_raw = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  miss_state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  scnd_miss_req_q = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  ifu_fetch_addr_int_f = _RAND_4[30:0];
  _RAND_5 = {1{`RANDOM}};
  ifc_iccm_access_f = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  iccm_dma_rvalid_in = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dma_iccm_req_f = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  perr_state = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  err_stop_state = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  reset_all_tags = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ifc_region_acc_fault_final_f = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  ifu_bus_rvalid_unq_ff = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  bus_ifu_bus_clk_en_ff = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  uncacheable_miss_ff = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  bus_data_beat_count = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ic_miss_buff_data_valid = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  imb_ff = _RAND_17[30:0];
  _RAND_18 = {1{`RANDOM}};
  last_data_recieved_ff = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  sel_mb_addr_ff = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  way_status_mb_scnd_ff = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  ifu_ic_rw_int_addr_ff = _RAND_21[6:0];
  _RAND_22 = {1{`RANDOM}};
  way_status_out_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  way_status_out_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  way_status_out_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  way_status_out_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  way_status_out_4 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  way_status_out_5 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  way_status_out_6 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  way_status_out_7 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  way_status_out_8 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  way_status_out_9 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  way_status_out_10 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  way_status_out_11 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  way_status_out_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  way_status_out_13 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  way_status_out_14 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  way_status_out_15 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  way_status_out_16 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  way_status_out_17 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  way_status_out_18 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  way_status_out_19 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  way_status_out_20 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  way_status_out_21 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  way_status_out_22 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  way_status_out_23 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  way_status_out_24 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  way_status_out_25 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  way_status_out_26 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  way_status_out_27 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  way_status_out_28 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  way_status_out_29 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  way_status_out_30 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  way_status_out_31 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  way_status_out_32 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  way_status_out_33 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  way_status_out_34 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  way_status_out_35 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  way_status_out_36 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  way_status_out_37 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  way_status_out_38 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  way_status_out_39 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  way_status_out_40 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  way_status_out_41 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  way_status_out_42 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  way_status_out_43 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  way_status_out_44 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  way_status_out_45 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  way_status_out_46 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  way_status_out_47 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  way_status_out_48 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  way_status_out_49 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  way_status_out_50 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  way_status_out_51 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  way_status_out_52 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  way_status_out_53 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  way_status_out_54 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  way_status_out_55 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  way_status_out_56 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  way_status_out_57 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  way_status_out_58 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  way_status_out_59 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  way_status_out_60 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  way_status_out_61 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  way_status_out_62 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  way_status_out_63 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  way_status_out_64 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  way_status_out_65 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  way_status_out_66 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  way_status_out_67 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  way_status_out_68 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  way_status_out_69 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  way_status_out_70 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  way_status_out_71 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  way_status_out_72 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  way_status_out_73 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  way_status_out_74 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  way_status_out_75 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  way_status_out_76 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  way_status_out_77 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  way_status_out_78 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  way_status_out_79 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  way_status_out_80 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  way_status_out_81 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  way_status_out_82 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  way_status_out_83 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  way_status_out_84 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  way_status_out_85 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  way_status_out_86 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  way_status_out_87 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  way_status_out_88 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  way_status_out_89 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  way_status_out_90 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  way_status_out_91 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  way_status_out_92 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  way_status_out_93 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  way_status_out_94 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  way_status_out_95 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  way_status_out_96 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  way_status_out_97 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  way_status_out_98 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  way_status_out_99 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  way_status_out_100 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  way_status_out_101 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  way_status_out_102 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  way_status_out_103 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  way_status_out_104 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  way_status_out_105 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  way_status_out_106 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  way_status_out_107 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  way_status_out_108 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  way_status_out_109 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  way_status_out_110 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  way_status_out_111 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  way_status_out_112 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  way_status_out_113 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  way_status_out_114 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  way_status_out_115 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  way_status_out_116 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  way_status_out_117 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  way_status_out_118 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  way_status_out_119 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  way_status_out_120 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  way_status_out_121 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  way_status_out_122 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  way_status_out_123 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  way_status_out_124 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  way_status_out_125 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  way_status_out_126 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  way_status_out_127 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  tagv_mb_scnd_ff = _RAND_150[1:0];
  _RAND_151 = {1{`RANDOM}};
  uncacheable_miss_scnd_ff = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  imb_scnd_ff = _RAND_152[30:0];
  _RAND_153 = {1{`RANDOM}};
  ifu_bus_rid_ff = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  ifu_bus_rresp_ff = _RAND_154[1:0];
  _RAND_155 = {1{`RANDOM}};
  ifu_wr_data_comb_err_ff = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  way_status_mb_ff = _RAND_156[0:0];
  _RAND_157 = {1{`RANDOM}};
  tagv_mb_ff = _RAND_157[1:0];
  _RAND_158 = {1{`RANDOM}};
  reset_ic_ff = _RAND_158[0:0];
  _RAND_159 = {1{`RANDOM}};
  fetch_uncacheable_ff = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  miss_addr = _RAND_160[25:0];
  _RAND_161 = {1{`RANDOM}};
  ifc_region_acc_fault_f = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  bus_rd_addr_count = _RAND_162[2:0];
  _RAND_163 = {1{`RANDOM}};
  ic_act_miss_f_delayed = _RAND_163[0:0];
  _RAND_164 = {2{`RANDOM}};
  ifu_bus_rdata_ff = _RAND_164[63:0];
  _RAND_165 = {1{`RANDOM}};
  ic_miss_buff_data_0 = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  ic_miss_buff_data_1 = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  ic_miss_buff_data_2 = _RAND_167[31:0];
  _RAND_168 = {1{`RANDOM}};
  ic_miss_buff_data_3 = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  ic_miss_buff_data_4 = _RAND_169[31:0];
  _RAND_170 = {1{`RANDOM}};
  ic_miss_buff_data_5 = _RAND_170[31:0];
  _RAND_171 = {1{`RANDOM}};
  ic_miss_buff_data_6 = _RAND_171[31:0];
  _RAND_172 = {1{`RANDOM}};
  ic_miss_buff_data_7 = _RAND_172[31:0];
  _RAND_173 = {1{`RANDOM}};
  ic_miss_buff_data_8 = _RAND_173[31:0];
  _RAND_174 = {1{`RANDOM}};
  ic_miss_buff_data_9 = _RAND_174[31:0];
  _RAND_175 = {1{`RANDOM}};
  ic_miss_buff_data_10 = _RAND_175[31:0];
  _RAND_176 = {1{`RANDOM}};
  ic_miss_buff_data_11 = _RAND_176[31:0];
  _RAND_177 = {1{`RANDOM}};
  ic_miss_buff_data_12 = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  ic_miss_buff_data_13 = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  ic_miss_buff_data_14 = _RAND_179[31:0];
  _RAND_180 = {1{`RANDOM}};
  ic_miss_buff_data_15 = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  ic_crit_wd_rdy_new_ff = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  ic_miss_buff_data_error = _RAND_182[7:0];
  _RAND_183 = {1{`RANDOM}};
  ic_debug_ict_array_sel_ff = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  ic_tag_valid_out_1_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  ic_tag_valid_out_1_1 = _RAND_185[0:0];
  _RAND_186 = {1{`RANDOM}};
  ic_tag_valid_out_1_2 = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  ic_tag_valid_out_1_3 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  ic_tag_valid_out_1_4 = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  ic_tag_valid_out_1_5 = _RAND_189[0:0];
  _RAND_190 = {1{`RANDOM}};
  ic_tag_valid_out_1_6 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  ic_tag_valid_out_1_7 = _RAND_191[0:0];
  _RAND_192 = {1{`RANDOM}};
  ic_tag_valid_out_1_8 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  ic_tag_valid_out_1_9 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  ic_tag_valid_out_1_10 = _RAND_194[0:0];
  _RAND_195 = {1{`RANDOM}};
  ic_tag_valid_out_1_11 = _RAND_195[0:0];
  _RAND_196 = {1{`RANDOM}};
  ic_tag_valid_out_1_12 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  ic_tag_valid_out_1_13 = _RAND_197[0:0];
  _RAND_198 = {1{`RANDOM}};
  ic_tag_valid_out_1_14 = _RAND_198[0:0];
  _RAND_199 = {1{`RANDOM}};
  ic_tag_valid_out_1_15 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  ic_tag_valid_out_1_16 = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  ic_tag_valid_out_1_17 = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  ic_tag_valid_out_1_18 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  ic_tag_valid_out_1_19 = _RAND_203[0:0];
  _RAND_204 = {1{`RANDOM}};
  ic_tag_valid_out_1_20 = _RAND_204[0:0];
  _RAND_205 = {1{`RANDOM}};
  ic_tag_valid_out_1_21 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  ic_tag_valid_out_1_22 = _RAND_206[0:0];
  _RAND_207 = {1{`RANDOM}};
  ic_tag_valid_out_1_23 = _RAND_207[0:0];
  _RAND_208 = {1{`RANDOM}};
  ic_tag_valid_out_1_24 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  ic_tag_valid_out_1_25 = _RAND_209[0:0];
  _RAND_210 = {1{`RANDOM}};
  ic_tag_valid_out_1_26 = _RAND_210[0:0];
  _RAND_211 = {1{`RANDOM}};
  ic_tag_valid_out_1_27 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  ic_tag_valid_out_1_28 = _RAND_212[0:0];
  _RAND_213 = {1{`RANDOM}};
  ic_tag_valid_out_1_29 = _RAND_213[0:0];
  _RAND_214 = {1{`RANDOM}};
  ic_tag_valid_out_1_30 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  ic_tag_valid_out_1_31 = _RAND_215[0:0];
  _RAND_216 = {1{`RANDOM}};
  ic_tag_valid_out_1_32 = _RAND_216[0:0];
  _RAND_217 = {1{`RANDOM}};
  ic_tag_valid_out_1_33 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  ic_tag_valid_out_1_34 = _RAND_218[0:0];
  _RAND_219 = {1{`RANDOM}};
  ic_tag_valid_out_1_35 = _RAND_219[0:0];
  _RAND_220 = {1{`RANDOM}};
  ic_tag_valid_out_1_36 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  ic_tag_valid_out_1_37 = _RAND_221[0:0];
  _RAND_222 = {1{`RANDOM}};
  ic_tag_valid_out_1_38 = _RAND_222[0:0];
  _RAND_223 = {1{`RANDOM}};
  ic_tag_valid_out_1_39 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  ic_tag_valid_out_1_40 = _RAND_224[0:0];
  _RAND_225 = {1{`RANDOM}};
  ic_tag_valid_out_1_41 = _RAND_225[0:0];
  _RAND_226 = {1{`RANDOM}};
  ic_tag_valid_out_1_42 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  ic_tag_valid_out_1_43 = _RAND_227[0:0];
  _RAND_228 = {1{`RANDOM}};
  ic_tag_valid_out_1_44 = _RAND_228[0:0];
  _RAND_229 = {1{`RANDOM}};
  ic_tag_valid_out_1_45 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  ic_tag_valid_out_1_46 = _RAND_230[0:0];
  _RAND_231 = {1{`RANDOM}};
  ic_tag_valid_out_1_47 = _RAND_231[0:0];
  _RAND_232 = {1{`RANDOM}};
  ic_tag_valid_out_1_48 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  ic_tag_valid_out_1_49 = _RAND_233[0:0];
  _RAND_234 = {1{`RANDOM}};
  ic_tag_valid_out_1_50 = _RAND_234[0:0];
  _RAND_235 = {1{`RANDOM}};
  ic_tag_valid_out_1_51 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  ic_tag_valid_out_1_52 = _RAND_236[0:0];
  _RAND_237 = {1{`RANDOM}};
  ic_tag_valid_out_1_53 = _RAND_237[0:0];
  _RAND_238 = {1{`RANDOM}};
  ic_tag_valid_out_1_54 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  ic_tag_valid_out_1_55 = _RAND_239[0:0];
  _RAND_240 = {1{`RANDOM}};
  ic_tag_valid_out_1_56 = _RAND_240[0:0];
  _RAND_241 = {1{`RANDOM}};
  ic_tag_valid_out_1_57 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  ic_tag_valid_out_1_58 = _RAND_242[0:0];
  _RAND_243 = {1{`RANDOM}};
  ic_tag_valid_out_1_59 = _RAND_243[0:0];
  _RAND_244 = {1{`RANDOM}};
  ic_tag_valid_out_1_60 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  ic_tag_valid_out_1_61 = _RAND_245[0:0];
  _RAND_246 = {1{`RANDOM}};
  ic_tag_valid_out_1_62 = _RAND_246[0:0];
  _RAND_247 = {1{`RANDOM}};
  ic_tag_valid_out_1_63 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  ic_tag_valid_out_1_64 = _RAND_248[0:0];
  _RAND_249 = {1{`RANDOM}};
  ic_tag_valid_out_1_65 = _RAND_249[0:0];
  _RAND_250 = {1{`RANDOM}};
  ic_tag_valid_out_1_66 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  ic_tag_valid_out_1_67 = _RAND_251[0:0];
  _RAND_252 = {1{`RANDOM}};
  ic_tag_valid_out_1_68 = _RAND_252[0:0];
  _RAND_253 = {1{`RANDOM}};
  ic_tag_valid_out_1_69 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  ic_tag_valid_out_1_70 = _RAND_254[0:0];
  _RAND_255 = {1{`RANDOM}};
  ic_tag_valid_out_1_71 = _RAND_255[0:0];
  _RAND_256 = {1{`RANDOM}};
  ic_tag_valid_out_1_72 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  ic_tag_valid_out_1_73 = _RAND_257[0:0];
  _RAND_258 = {1{`RANDOM}};
  ic_tag_valid_out_1_74 = _RAND_258[0:0];
  _RAND_259 = {1{`RANDOM}};
  ic_tag_valid_out_1_75 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  ic_tag_valid_out_1_76 = _RAND_260[0:0];
  _RAND_261 = {1{`RANDOM}};
  ic_tag_valid_out_1_77 = _RAND_261[0:0];
  _RAND_262 = {1{`RANDOM}};
  ic_tag_valid_out_1_78 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  ic_tag_valid_out_1_79 = _RAND_263[0:0];
  _RAND_264 = {1{`RANDOM}};
  ic_tag_valid_out_1_80 = _RAND_264[0:0];
  _RAND_265 = {1{`RANDOM}};
  ic_tag_valid_out_1_81 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  ic_tag_valid_out_1_82 = _RAND_266[0:0];
  _RAND_267 = {1{`RANDOM}};
  ic_tag_valid_out_1_83 = _RAND_267[0:0];
  _RAND_268 = {1{`RANDOM}};
  ic_tag_valid_out_1_84 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  ic_tag_valid_out_1_85 = _RAND_269[0:0];
  _RAND_270 = {1{`RANDOM}};
  ic_tag_valid_out_1_86 = _RAND_270[0:0];
  _RAND_271 = {1{`RANDOM}};
  ic_tag_valid_out_1_87 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  ic_tag_valid_out_1_88 = _RAND_272[0:0];
  _RAND_273 = {1{`RANDOM}};
  ic_tag_valid_out_1_89 = _RAND_273[0:0];
  _RAND_274 = {1{`RANDOM}};
  ic_tag_valid_out_1_90 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  ic_tag_valid_out_1_91 = _RAND_275[0:0];
  _RAND_276 = {1{`RANDOM}};
  ic_tag_valid_out_1_92 = _RAND_276[0:0];
  _RAND_277 = {1{`RANDOM}};
  ic_tag_valid_out_1_93 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  ic_tag_valid_out_1_94 = _RAND_278[0:0];
  _RAND_279 = {1{`RANDOM}};
  ic_tag_valid_out_1_95 = _RAND_279[0:0];
  _RAND_280 = {1{`RANDOM}};
  ic_tag_valid_out_1_96 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  ic_tag_valid_out_1_97 = _RAND_281[0:0];
  _RAND_282 = {1{`RANDOM}};
  ic_tag_valid_out_1_98 = _RAND_282[0:0];
  _RAND_283 = {1{`RANDOM}};
  ic_tag_valid_out_1_99 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  ic_tag_valid_out_1_100 = _RAND_284[0:0];
  _RAND_285 = {1{`RANDOM}};
  ic_tag_valid_out_1_101 = _RAND_285[0:0];
  _RAND_286 = {1{`RANDOM}};
  ic_tag_valid_out_1_102 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  ic_tag_valid_out_1_103 = _RAND_287[0:0];
  _RAND_288 = {1{`RANDOM}};
  ic_tag_valid_out_1_104 = _RAND_288[0:0];
  _RAND_289 = {1{`RANDOM}};
  ic_tag_valid_out_1_105 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  ic_tag_valid_out_1_106 = _RAND_290[0:0];
  _RAND_291 = {1{`RANDOM}};
  ic_tag_valid_out_1_107 = _RAND_291[0:0];
  _RAND_292 = {1{`RANDOM}};
  ic_tag_valid_out_1_108 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  ic_tag_valid_out_1_109 = _RAND_293[0:0];
  _RAND_294 = {1{`RANDOM}};
  ic_tag_valid_out_1_110 = _RAND_294[0:0];
  _RAND_295 = {1{`RANDOM}};
  ic_tag_valid_out_1_111 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  ic_tag_valid_out_1_112 = _RAND_296[0:0];
  _RAND_297 = {1{`RANDOM}};
  ic_tag_valid_out_1_113 = _RAND_297[0:0];
  _RAND_298 = {1{`RANDOM}};
  ic_tag_valid_out_1_114 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  ic_tag_valid_out_1_115 = _RAND_299[0:0];
  _RAND_300 = {1{`RANDOM}};
  ic_tag_valid_out_1_116 = _RAND_300[0:0];
  _RAND_301 = {1{`RANDOM}};
  ic_tag_valid_out_1_117 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  ic_tag_valid_out_1_118 = _RAND_302[0:0];
  _RAND_303 = {1{`RANDOM}};
  ic_tag_valid_out_1_119 = _RAND_303[0:0];
  _RAND_304 = {1{`RANDOM}};
  ic_tag_valid_out_1_120 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  ic_tag_valid_out_1_121 = _RAND_305[0:0];
  _RAND_306 = {1{`RANDOM}};
  ic_tag_valid_out_1_122 = _RAND_306[0:0];
  _RAND_307 = {1{`RANDOM}};
  ic_tag_valid_out_1_123 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  ic_tag_valid_out_1_124 = _RAND_308[0:0];
  _RAND_309 = {1{`RANDOM}};
  ic_tag_valid_out_1_125 = _RAND_309[0:0];
  _RAND_310 = {1{`RANDOM}};
  ic_tag_valid_out_1_126 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  ic_tag_valid_out_1_127 = _RAND_311[0:0];
  _RAND_312 = {1{`RANDOM}};
  ic_tag_valid_out_0_0 = _RAND_312[0:0];
  _RAND_313 = {1{`RANDOM}};
  ic_tag_valid_out_0_1 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  ic_tag_valid_out_0_2 = _RAND_314[0:0];
  _RAND_315 = {1{`RANDOM}};
  ic_tag_valid_out_0_3 = _RAND_315[0:0];
  _RAND_316 = {1{`RANDOM}};
  ic_tag_valid_out_0_4 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  ic_tag_valid_out_0_5 = _RAND_317[0:0];
  _RAND_318 = {1{`RANDOM}};
  ic_tag_valid_out_0_6 = _RAND_318[0:0];
  _RAND_319 = {1{`RANDOM}};
  ic_tag_valid_out_0_7 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  ic_tag_valid_out_0_8 = _RAND_320[0:0];
  _RAND_321 = {1{`RANDOM}};
  ic_tag_valid_out_0_9 = _RAND_321[0:0];
  _RAND_322 = {1{`RANDOM}};
  ic_tag_valid_out_0_10 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  ic_tag_valid_out_0_11 = _RAND_323[0:0];
  _RAND_324 = {1{`RANDOM}};
  ic_tag_valid_out_0_12 = _RAND_324[0:0];
  _RAND_325 = {1{`RANDOM}};
  ic_tag_valid_out_0_13 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  ic_tag_valid_out_0_14 = _RAND_326[0:0];
  _RAND_327 = {1{`RANDOM}};
  ic_tag_valid_out_0_15 = _RAND_327[0:0];
  _RAND_328 = {1{`RANDOM}};
  ic_tag_valid_out_0_16 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  ic_tag_valid_out_0_17 = _RAND_329[0:0];
  _RAND_330 = {1{`RANDOM}};
  ic_tag_valid_out_0_18 = _RAND_330[0:0];
  _RAND_331 = {1{`RANDOM}};
  ic_tag_valid_out_0_19 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  ic_tag_valid_out_0_20 = _RAND_332[0:0];
  _RAND_333 = {1{`RANDOM}};
  ic_tag_valid_out_0_21 = _RAND_333[0:0];
  _RAND_334 = {1{`RANDOM}};
  ic_tag_valid_out_0_22 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  ic_tag_valid_out_0_23 = _RAND_335[0:0];
  _RAND_336 = {1{`RANDOM}};
  ic_tag_valid_out_0_24 = _RAND_336[0:0];
  _RAND_337 = {1{`RANDOM}};
  ic_tag_valid_out_0_25 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  ic_tag_valid_out_0_26 = _RAND_338[0:0];
  _RAND_339 = {1{`RANDOM}};
  ic_tag_valid_out_0_27 = _RAND_339[0:0];
  _RAND_340 = {1{`RANDOM}};
  ic_tag_valid_out_0_28 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  ic_tag_valid_out_0_29 = _RAND_341[0:0];
  _RAND_342 = {1{`RANDOM}};
  ic_tag_valid_out_0_30 = _RAND_342[0:0];
  _RAND_343 = {1{`RANDOM}};
  ic_tag_valid_out_0_31 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  ic_tag_valid_out_0_32 = _RAND_344[0:0];
  _RAND_345 = {1{`RANDOM}};
  ic_tag_valid_out_0_33 = _RAND_345[0:0];
  _RAND_346 = {1{`RANDOM}};
  ic_tag_valid_out_0_34 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  ic_tag_valid_out_0_35 = _RAND_347[0:0];
  _RAND_348 = {1{`RANDOM}};
  ic_tag_valid_out_0_36 = _RAND_348[0:0];
  _RAND_349 = {1{`RANDOM}};
  ic_tag_valid_out_0_37 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  ic_tag_valid_out_0_38 = _RAND_350[0:0];
  _RAND_351 = {1{`RANDOM}};
  ic_tag_valid_out_0_39 = _RAND_351[0:0];
  _RAND_352 = {1{`RANDOM}};
  ic_tag_valid_out_0_40 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  ic_tag_valid_out_0_41 = _RAND_353[0:0];
  _RAND_354 = {1{`RANDOM}};
  ic_tag_valid_out_0_42 = _RAND_354[0:0];
  _RAND_355 = {1{`RANDOM}};
  ic_tag_valid_out_0_43 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  ic_tag_valid_out_0_44 = _RAND_356[0:0];
  _RAND_357 = {1{`RANDOM}};
  ic_tag_valid_out_0_45 = _RAND_357[0:0];
  _RAND_358 = {1{`RANDOM}};
  ic_tag_valid_out_0_46 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  ic_tag_valid_out_0_47 = _RAND_359[0:0];
  _RAND_360 = {1{`RANDOM}};
  ic_tag_valid_out_0_48 = _RAND_360[0:0];
  _RAND_361 = {1{`RANDOM}};
  ic_tag_valid_out_0_49 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  ic_tag_valid_out_0_50 = _RAND_362[0:0];
  _RAND_363 = {1{`RANDOM}};
  ic_tag_valid_out_0_51 = _RAND_363[0:0];
  _RAND_364 = {1{`RANDOM}};
  ic_tag_valid_out_0_52 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  ic_tag_valid_out_0_53 = _RAND_365[0:0];
  _RAND_366 = {1{`RANDOM}};
  ic_tag_valid_out_0_54 = _RAND_366[0:0];
  _RAND_367 = {1{`RANDOM}};
  ic_tag_valid_out_0_55 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  ic_tag_valid_out_0_56 = _RAND_368[0:0];
  _RAND_369 = {1{`RANDOM}};
  ic_tag_valid_out_0_57 = _RAND_369[0:0];
  _RAND_370 = {1{`RANDOM}};
  ic_tag_valid_out_0_58 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  ic_tag_valid_out_0_59 = _RAND_371[0:0];
  _RAND_372 = {1{`RANDOM}};
  ic_tag_valid_out_0_60 = _RAND_372[0:0];
  _RAND_373 = {1{`RANDOM}};
  ic_tag_valid_out_0_61 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  ic_tag_valid_out_0_62 = _RAND_374[0:0];
  _RAND_375 = {1{`RANDOM}};
  ic_tag_valid_out_0_63 = _RAND_375[0:0];
  _RAND_376 = {1{`RANDOM}};
  ic_tag_valid_out_0_64 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  ic_tag_valid_out_0_65 = _RAND_377[0:0];
  _RAND_378 = {1{`RANDOM}};
  ic_tag_valid_out_0_66 = _RAND_378[0:0];
  _RAND_379 = {1{`RANDOM}};
  ic_tag_valid_out_0_67 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  ic_tag_valid_out_0_68 = _RAND_380[0:0];
  _RAND_381 = {1{`RANDOM}};
  ic_tag_valid_out_0_69 = _RAND_381[0:0];
  _RAND_382 = {1{`RANDOM}};
  ic_tag_valid_out_0_70 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  ic_tag_valid_out_0_71 = _RAND_383[0:0];
  _RAND_384 = {1{`RANDOM}};
  ic_tag_valid_out_0_72 = _RAND_384[0:0];
  _RAND_385 = {1{`RANDOM}};
  ic_tag_valid_out_0_73 = _RAND_385[0:0];
  _RAND_386 = {1{`RANDOM}};
  ic_tag_valid_out_0_74 = _RAND_386[0:0];
  _RAND_387 = {1{`RANDOM}};
  ic_tag_valid_out_0_75 = _RAND_387[0:0];
  _RAND_388 = {1{`RANDOM}};
  ic_tag_valid_out_0_76 = _RAND_388[0:0];
  _RAND_389 = {1{`RANDOM}};
  ic_tag_valid_out_0_77 = _RAND_389[0:0];
  _RAND_390 = {1{`RANDOM}};
  ic_tag_valid_out_0_78 = _RAND_390[0:0];
  _RAND_391 = {1{`RANDOM}};
  ic_tag_valid_out_0_79 = _RAND_391[0:0];
  _RAND_392 = {1{`RANDOM}};
  ic_tag_valid_out_0_80 = _RAND_392[0:0];
  _RAND_393 = {1{`RANDOM}};
  ic_tag_valid_out_0_81 = _RAND_393[0:0];
  _RAND_394 = {1{`RANDOM}};
  ic_tag_valid_out_0_82 = _RAND_394[0:0];
  _RAND_395 = {1{`RANDOM}};
  ic_tag_valid_out_0_83 = _RAND_395[0:0];
  _RAND_396 = {1{`RANDOM}};
  ic_tag_valid_out_0_84 = _RAND_396[0:0];
  _RAND_397 = {1{`RANDOM}};
  ic_tag_valid_out_0_85 = _RAND_397[0:0];
  _RAND_398 = {1{`RANDOM}};
  ic_tag_valid_out_0_86 = _RAND_398[0:0];
  _RAND_399 = {1{`RANDOM}};
  ic_tag_valid_out_0_87 = _RAND_399[0:0];
  _RAND_400 = {1{`RANDOM}};
  ic_tag_valid_out_0_88 = _RAND_400[0:0];
  _RAND_401 = {1{`RANDOM}};
  ic_tag_valid_out_0_89 = _RAND_401[0:0];
  _RAND_402 = {1{`RANDOM}};
  ic_tag_valid_out_0_90 = _RAND_402[0:0];
  _RAND_403 = {1{`RANDOM}};
  ic_tag_valid_out_0_91 = _RAND_403[0:0];
  _RAND_404 = {1{`RANDOM}};
  ic_tag_valid_out_0_92 = _RAND_404[0:0];
  _RAND_405 = {1{`RANDOM}};
  ic_tag_valid_out_0_93 = _RAND_405[0:0];
  _RAND_406 = {1{`RANDOM}};
  ic_tag_valid_out_0_94 = _RAND_406[0:0];
  _RAND_407 = {1{`RANDOM}};
  ic_tag_valid_out_0_95 = _RAND_407[0:0];
  _RAND_408 = {1{`RANDOM}};
  ic_tag_valid_out_0_96 = _RAND_408[0:0];
  _RAND_409 = {1{`RANDOM}};
  ic_tag_valid_out_0_97 = _RAND_409[0:0];
  _RAND_410 = {1{`RANDOM}};
  ic_tag_valid_out_0_98 = _RAND_410[0:0];
  _RAND_411 = {1{`RANDOM}};
  ic_tag_valid_out_0_99 = _RAND_411[0:0];
  _RAND_412 = {1{`RANDOM}};
  ic_tag_valid_out_0_100 = _RAND_412[0:0];
  _RAND_413 = {1{`RANDOM}};
  ic_tag_valid_out_0_101 = _RAND_413[0:0];
  _RAND_414 = {1{`RANDOM}};
  ic_tag_valid_out_0_102 = _RAND_414[0:0];
  _RAND_415 = {1{`RANDOM}};
  ic_tag_valid_out_0_103 = _RAND_415[0:0];
  _RAND_416 = {1{`RANDOM}};
  ic_tag_valid_out_0_104 = _RAND_416[0:0];
  _RAND_417 = {1{`RANDOM}};
  ic_tag_valid_out_0_105 = _RAND_417[0:0];
  _RAND_418 = {1{`RANDOM}};
  ic_tag_valid_out_0_106 = _RAND_418[0:0];
  _RAND_419 = {1{`RANDOM}};
  ic_tag_valid_out_0_107 = _RAND_419[0:0];
  _RAND_420 = {1{`RANDOM}};
  ic_tag_valid_out_0_108 = _RAND_420[0:0];
  _RAND_421 = {1{`RANDOM}};
  ic_tag_valid_out_0_109 = _RAND_421[0:0];
  _RAND_422 = {1{`RANDOM}};
  ic_tag_valid_out_0_110 = _RAND_422[0:0];
  _RAND_423 = {1{`RANDOM}};
  ic_tag_valid_out_0_111 = _RAND_423[0:0];
  _RAND_424 = {1{`RANDOM}};
  ic_tag_valid_out_0_112 = _RAND_424[0:0];
  _RAND_425 = {1{`RANDOM}};
  ic_tag_valid_out_0_113 = _RAND_425[0:0];
  _RAND_426 = {1{`RANDOM}};
  ic_tag_valid_out_0_114 = _RAND_426[0:0];
  _RAND_427 = {1{`RANDOM}};
  ic_tag_valid_out_0_115 = _RAND_427[0:0];
  _RAND_428 = {1{`RANDOM}};
  ic_tag_valid_out_0_116 = _RAND_428[0:0];
  _RAND_429 = {1{`RANDOM}};
  ic_tag_valid_out_0_117 = _RAND_429[0:0];
  _RAND_430 = {1{`RANDOM}};
  ic_tag_valid_out_0_118 = _RAND_430[0:0];
  _RAND_431 = {1{`RANDOM}};
  ic_tag_valid_out_0_119 = _RAND_431[0:0];
  _RAND_432 = {1{`RANDOM}};
  ic_tag_valid_out_0_120 = _RAND_432[0:0];
  _RAND_433 = {1{`RANDOM}};
  ic_tag_valid_out_0_121 = _RAND_433[0:0];
  _RAND_434 = {1{`RANDOM}};
  ic_tag_valid_out_0_122 = _RAND_434[0:0];
  _RAND_435 = {1{`RANDOM}};
  ic_tag_valid_out_0_123 = _RAND_435[0:0];
  _RAND_436 = {1{`RANDOM}};
  ic_tag_valid_out_0_124 = _RAND_436[0:0];
  _RAND_437 = {1{`RANDOM}};
  ic_tag_valid_out_0_125 = _RAND_437[0:0];
  _RAND_438 = {1{`RANDOM}};
  ic_tag_valid_out_0_126 = _RAND_438[0:0];
  _RAND_439 = {1{`RANDOM}};
  ic_tag_valid_out_0_127 = _RAND_439[0:0];
  _RAND_440 = {1{`RANDOM}};
  ic_debug_way_ff = _RAND_440[1:0];
  _RAND_441 = {1{`RANDOM}};
  ic_debug_rd_en_ff = _RAND_441[0:0];
  _RAND_442 = {3{`RANDOM}};
  _T_1209 = _RAND_442[70:0];
  _RAND_443 = {1{`RANDOM}};
  perr_ic_index_ff = _RAND_443[6:0];
  _RAND_444 = {1{`RANDOM}};
  dma_sb_err_state_ff = _RAND_444[0:0];
  _RAND_445 = {1{`RANDOM}};
  ifu_bus_cmd_valid = _RAND_445[0:0];
  _RAND_446 = {1{`RANDOM}};
  bus_cmd_beat_count = _RAND_446[2:0];
  _RAND_447 = {1{`RANDOM}};
  ifu_bus_arready_unq_ff = _RAND_447[0:0];
  _RAND_448 = {1{`RANDOM}};
  ifu_bus_arvalid_ff = _RAND_448[0:0];
  _RAND_449 = {1{`RANDOM}};
  ifc_dma_access_ok_prev = _RAND_449[0:0];
  _RAND_450 = {2{`RANDOM}};
  iccm_ecc_corr_data_ff = _RAND_450[38:0];
  _RAND_451 = {1{`RANDOM}};
  dma_mem_addr_ff = _RAND_451[1:0];
  _RAND_452 = {1{`RANDOM}};
  dma_mem_tag_ff = _RAND_452[2:0];
  _RAND_453 = {1{`RANDOM}};
  iccm_dma_rtag_temp = _RAND_453[2:0];
  _RAND_454 = {1{`RANDOM}};
  iccm_dma_rvalid_temp = _RAND_454[0:0];
  _RAND_455 = {2{`RANDOM}};
  iccm_dma_rdata_temp = _RAND_455[63:0];
  _RAND_456 = {1{`RANDOM}};
  iccm_ecc_corr_index_ff = _RAND_456[13:0];
  _RAND_457 = {1{`RANDOM}};
  iccm_rd_ecc_single_err_ff = _RAND_457[0:0];
  _RAND_458 = {1{`RANDOM}};
  iccm_rw_addr_f = _RAND_458[13:0];
  _RAND_459 = {1{`RANDOM}};
  ifu_status_wr_addr_ff = _RAND_459[6:0];
  _RAND_460 = {1{`RANDOM}};
  way_status_wr_en_ff = _RAND_460[0:0];
  _RAND_461 = {1{`RANDOM}};
  way_status_new_ff = _RAND_461[0:0];
  _RAND_462 = {1{`RANDOM}};
  ifu_tag_wren_ff = _RAND_462[1:0];
  _RAND_463 = {1{`RANDOM}};
  ic_valid_ff = _RAND_463[0:0];
  _RAND_464 = {1{`RANDOM}};
  _T_10581 = _RAND_464[0:0];
  _RAND_465 = {1{`RANDOM}};
  _T_10582 = _RAND_465[0:0];
  _RAND_466 = {1{`RANDOM}};
  _T_10583 = _RAND_466[0:0];
  _RAND_467 = {1{`RANDOM}};
  _T_10587 = _RAND_467[0:0];
  _RAND_468 = {1{`RANDOM}};
  _T_10588 = _RAND_468[0:0];
  _RAND_469 = {1{`RANDOM}};
  _T_10611 = _RAND_469[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flush_final_f <= 1'h0;
    end else begin
      flush_final_f <= io_exu_flush_final;
    end
    if (reset) begin
      ifc_fetch_req_f_raw <= 1'h0;
    end else begin
      ifc_fetch_req_f_raw <= ifc_fetch_req_qual_bf;
    end
    if (reset) begin
      miss_state <= 3'h0;
    end else if (miss_state_en) begin
      if (_T_24) begin
        if (_T_26) begin
          miss_state <= 3'h1;
        end else begin
          miss_state <= 3'h2;
        end
      end else if (_T_31) begin
        if (_T_36) begin
          miss_state <= 3'h0;
        end else if (_T_40) begin
          miss_state <= 3'h3;
        end else if (_T_47) begin
          miss_state <= 3'h4;
        end else if (_T_51) begin
          miss_state <= 3'h0;
        end else if (_T_61) begin
          miss_state <= 3'h6;
        end else if (_T_71) begin
          miss_state <= 3'h6;
        end else if (_T_79) begin
          miss_state <= 3'h0;
        end else if (_T_84) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_102) begin
        miss_state <= 3'h0;
      end else if (_T_106) begin
        if (_T_113) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_121) begin
        if (_T_126) begin
          miss_state <= 3'h2;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_132) begin
        if (_T_137) begin
          miss_state <= 3'h5;
        end else if (_T_143) begin
          miss_state <= 3'h7;
        end else begin
          miss_state <= 3'h0;
        end
      end else if (_T_151) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h1;
        end
      end else if (_T_160) begin
        if (io_dec_tlu_force_halt) begin
          miss_state <= 3'h0;
        end else if (io_exu_flush_final) begin
          if (_T_32) begin
            miss_state <= 3'h0;
          end else begin
            miss_state <= 3'h2;
          end
        end else begin
          miss_state <= 3'h0;
        end
      end else begin
        miss_state <= 3'h0;
      end
    end
    if (reset) begin
      ifu_fetch_addr_int_f <= 31'h0;
    end else begin
      ifu_fetch_addr_int_f <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifc_iccm_access_f <= 1'h0;
    end else begin
      ifc_iccm_access_f <= io_ifc_iccm_access_bf;
    end
    if (reset) begin
      ifc_region_acc_fault_final_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_final_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      ifu_bus_rvalid_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rvalid_unq_ff <= io_ifu_axi_rvalid;
    end
    if (reset) begin
      uncacheable_miss_ff <= 1'h0;
    end else if (scnd_miss_req) begin
      uncacheable_miss_ff <= uncacheable_miss_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      uncacheable_miss_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (scnd_miss_req) begin
      imb_ff <= imb_scnd_ff;
    end else if (!(sel_hold_imb)) begin
      imb_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      way_status_mb_scnd_ff <= 1'h0;
    end else if (!(_T_19)) begin
      way_status_mb_scnd_ff <= way_status;
    end
    if (reset) begin
      way_status_out_0 <= 1'h0;
    end else if (_T_4172) begin
      way_status_out_0 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_1 <= 1'h0;
    end else if (_T_4177) begin
      way_status_out_1 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_2 <= 1'h0;
    end else if (_T_4182) begin
      way_status_out_2 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_3 <= 1'h0;
    end else if (_T_4187) begin
      way_status_out_3 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_4 <= 1'h0;
    end else if (_T_4192) begin
      way_status_out_4 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_5 <= 1'h0;
    end else if (_T_4197) begin
      way_status_out_5 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_6 <= 1'h0;
    end else if (_T_4202) begin
      way_status_out_6 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_7 <= 1'h0;
    end else if (_T_4207) begin
      way_status_out_7 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_8 <= 1'h0;
    end else if (_T_4212) begin
      way_status_out_8 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_9 <= 1'h0;
    end else if (_T_4217) begin
      way_status_out_9 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_10 <= 1'h0;
    end else if (_T_4222) begin
      way_status_out_10 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_11 <= 1'h0;
    end else if (_T_4227) begin
      way_status_out_11 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_12 <= 1'h0;
    end else if (_T_4232) begin
      way_status_out_12 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_13 <= 1'h0;
    end else if (_T_4237) begin
      way_status_out_13 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_14 <= 1'h0;
    end else if (_T_4242) begin
      way_status_out_14 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_15 <= 1'h0;
    end else if (_T_4247) begin
      way_status_out_15 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_16 <= 1'h0;
    end else if (_T_4252) begin
      way_status_out_16 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_17 <= 1'h0;
    end else if (_T_4257) begin
      way_status_out_17 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_18 <= 1'h0;
    end else if (_T_4262) begin
      way_status_out_18 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_19 <= 1'h0;
    end else if (_T_4267) begin
      way_status_out_19 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_20 <= 1'h0;
    end else if (_T_4272) begin
      way_status_out_20 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_21 <= 1'h0;
    end else if (_T_4277) begin
      way_status_out_21 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_22 <= 1'h0;
    end else if (_T_4282) begin
      way_status_out_22 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_23 <= 1'h0;
    end else if (_T_4287) begin
      way_status_out_23 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_24 <= 1'h0;
    end else if (_T_4292) begin
      way_status_out_24 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_25 <= 1'h0;
    end else if (_T_4297) begin
      way_status_out_25 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_26 <= 1'h0;
    end else if (_T_4302) begin
      way_status_out_26 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_27 <= 1'h0;
    end else if (_T_4307) begin
      way_status_out_27 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_28 <= 1'h0;
    end else if (_T_4312) begin
      way_status_out_28 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_29 <= 1'h0;
    end else if (_T_4317) begin
      way_status_out_29 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_30 <= 1'h0;
    end else if (_T_4322) begin
      way_status_out_30 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_31 <= 1'h0;
    end else if (_T_4327) begin
      way_status_out_31 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_32 <= 1'h0;
    end else if (_T_4332) begin
      way_status_out_32 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_33 <= 1'h0;
    end else if (_T_4337) begin
      way_status_out_33 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_34 <= 1'h0;
    end else if (_T_4342) begin
      way_status_out_34 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_35 <= 1'h0;
    end else if (_T_4347) begin
      way_status_out_35 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_36 <= 1'h0;
    end else if (_T_4352) begin
      way_status_out_36 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_37 <= 1'h0;
    end else if (_T_4357) begin
      way_status_out_37 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_38 <= 1'h0;
    end else if (_T_4362) begin
      way_status_out_38 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_39 <= 1'h0;
    end else if (_T_4367) begin
      way_status_out_39 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_40 <= 1'h0;
    end else if (_T_4372) begin
      way_status_out_40 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_41 <= 1'h0;
    end else if (_T_4377) begin
      way_status_out_41 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_42 <= 1'h0;
    end else if (_T_4382) begin
      way_status_out_42 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_43 <= 1'h0;
    end else if (_T_4387) begin
      way_status_out_43 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_44 <= 1'h0;
    end else if (_T_4392) begin
      way_status_out_44 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_45 <= 1'h0;
    end else if (_T_4397) begin
      way_status_out_45 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_46 <= 1'h0;
    end else if (_T_4402) begin
      way_status_out_46 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_47 <= 1'h0;
    end else if (_T_4407) begin
      way_status_out_47 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_48 <= 1'h0;
    end else if (_T_4412) begin
      way_status_out_48 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_49 <= 1'h0;
    end else if (_T_4417) begin
      way_status_out_49 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_50 <= 1'h0;
    end else if (_T_4422) begin
      way_status_out_50 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_51 <= 1'h0;
    end else if (_T_4427) begin
      way_status_out_51 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_52 <= 1'h0;
    end else if (_T_4432) begin
      way_status_out_52 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_53 <= 1'h0;
    end else if (_T_4437) begin
      way_status_out_53 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_54 <= 1'h0;
    end else if (_T_4442) begin
      way_status_out_54 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_55 <= 1'h0;
    end else if (_T_4447) begin
      way_status_out_55 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_56 <= 1'h0;
    end else if (_T_4452) begin
      way_status_out_56 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_57 <= 1'h0;
    end else if (_T_4457) begin
      way_status_out_57 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_58 <= 1'h0;
    end else if (_T_4462) begin
      way_status_out_58 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_59 <= 1'h0;
    end else if (_T_4467) begin
      way_status_out_59 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_60 <= 1'h0;
    end else if (_T_4472) begin
      way_status_out_60 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_61 <= 1'h0;
    end else if (_T_4477) begin
      way_status_out_61 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_62 <= 1'h0;
    end else if (_T_4482) begin
      way_status_out_62 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_63 <= 1'h0;
    end else if (_T_4487) begin
      way_status_out_63 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_64 <= 1'h0;
    end else if (_T_4492) begin
      way_status_out_64 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_65 <= 1'h0;
    end else if (_T_4497) begin
      way_status_out_65 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_66 <= 1'h0;
    end else if (_T_4502) begin
      way_status_out_66 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_67 <= 1'h0;
    end else if (_T_4507) begin
      way_status_out_67 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_68 <= 1'h0;
    end else if (_T_4512) begin
      way_status_out_68 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_69 <= 1'h0;
    end else if (_T_4517) begin
      way_status_out_69 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_70 <= 1'h0;
    end else if (_T_4522) begin
      way_status_out_70 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_71 <= 1'h0;
    end else if (_T_4527) begin
      way_status_out_71 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_72 <= 1'h0;
    end else if (_T_4532) begin
      way_status_out_72 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_73 <= 1'h0;
    end else if (_T_4537) begin
      way_status_out_73 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_74 <= 1'h0;
    end else if (_T_4542) begin
      way_status_out_74 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_75 <= 1'h0;
    end else if (_T_4547) begin
      way_status_out_75 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_76 <= 1'h0;
    end else if (_T_4552) begin
      way_status_out_76 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_77 <= 1'h0;
    end else if (_T_4557) begin
      way_status_out_77 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_78 <= 1'h0;
    end else if (_T_4562) begin
      way_status_out_78 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_79 <= 1'h0;
    end else if (_T_4567) begin
      way_status_out_79 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_80 <= 1'h0;
    end else if (_T_4572) begin
      way_status_out_80 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_81 <= 1'h0;
    end else if (_T_4577) begin
      way_status_out_81 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_82 <= 1'h0;
    end else if (_T_4582) begin
      way_status_out_82 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_83 <= 1'h0;
    end else if (_T_4587) begin
      way_status_out_83 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_84 <= 1'h0;
    end else if (_T_4592) begin
      way_status_out_84 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_85 <= 1'h0;
    end else if (_T_4597) begin
      way_status_out_85 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_86 <= 1'h0;
    end else if (_T_4602) begin
      way_status_out_86 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_87 <= 1'h0;
    end else if (_T_4607) begin
      way_status_out_87 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_88 <= 1'h0;
    end else if (_T_4612) begin
      way_status_out_88 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_89 <= 1'h0;
    end else if (_T_4617) begin
      way_status_out_89 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_90 <= 1'h0;
    end else if (_T_4622) begin
      way_status_out_90 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_91 <= 1'h0;
    end else if (_T_4627) begin
      way_status_out_91 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_92 <= 1'h0;
    end else if (_T_4632) begin
      way_status_out_92 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_93 <= 1'h0;
    end else if (_T_4637) begin
      way_status_out_93 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_94 <= 1'h0;
    end else if (_T_4642) begin
      way_status_out_94 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_95 <= 1'h0;
    end else if (_T_4647) begin
      way_status_out_95 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_96 <= 1'h0;
    end else if (_T_4652) begin
      way_status_out_96 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_97 <= 1'h0;
    end else if (_T_4657) begin
      way_status_out_97 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_98 <= 1'h0;
    end else if (_T_4662) begin
      way_status_out_98 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_99 <= 1'h0;
    end else if (_T_4667) begin
      way_status_out_99 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_100 <= 1'h0;
    end else if (_T_4672) begin
      way_status_out_100 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_101 <= 1'h0;
    end else if (_T_4677) begin
      way_status_out_101 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_102 <= 1'h0;
    end else if (_T_4682) begin
      way_status_out_102 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_103 <= 1'h0;
    end else if (_T_4687) begin
      way_status_out_103 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_104 <= 1'h0;
    end else if (_T_4692) begin
      way_status_out_104 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_105 <= 1'h0;
    end else if (_T_4697) begin
      way_status_out_105 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_106 <= 1'h0;
    end else if (_T_4702) begin
      way_status_out_106 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_107 <= 1'h0;
    end else if (_T_4707) begin
      way_status_out_107 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_108 <= 1'h0;
    end else if (_T_4712) begin
      way_status_out_108 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_109 <= 1'h0;
    end else if (_T_4717) begin
      way_status_out_109 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_110 <= 1'h0;
    end else if (_T_4722) begin
      way_status_out_110 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_111 <= 1'h0;
    end else if (_T_4727) begin
      way_status_out_111 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_112 <= 1'h0;
    end else if (_T_4732) begin
      way_status_out_112 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_113 <= 1'h0;
    end else if (_T_4737) begin
      way_status_out_113 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_114 <= 1'h0;
    end else if (_T_4742) begin
      way_status_out_114 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_115 <= 1'h0;
    end else if (_T_4747) begin
      way_status_out_115 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_116 <= 1'h0;
    end else if (_T_4752) begin
      way_status_out_116 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_117 <= 1'h0;
    end else if (_T_4757) begin
      way_status_out_117 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_118 <= 1'h0;
    end else if (_T_4762) begin
      way_status_out_118 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_119 <= 1'h0;
    end else if (_T_4767) begin
      way_status_out_119 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_120 <= 1'h0;
    end else if (_T_4772) begin
      way_status_out_120 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_121 <= 1'h0;
    end else if (_T_4777) begin
      way_status_out_121 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_122 <= 1'h0;
    end else if (_T_4782) begin
      way_status_out_122 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_123 <= 1'h0;
    end else if (_T_4787) begin
      way_status_out_123 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_124 <= 1'h0;
    end else if (_T_4792) begin
      way_status_out_124 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_125 <= 1'h0;
    end else if (_T_4797) begin
      way_status_out_125 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_126 <= 1'h0;
    end else if (_T_4802) begin
      way_status_out_126 <= way_status_new_ff;
    end
    if (reset) begin
      way_status_out_127 <= 1'h0;
    end else if (_T_4807) begin
      way_status_out_127 <= way_status_new_ff;
    end
    if (reset) begin
      tagv_mb_scnd_ff <= 2'h0;
    end else if (!(_T_19)) begin
      tagv_mb_scnd_ff <= _T_198;
    end
    if (reset) begin
      uncacheable_miss_scnd_ff <= 1'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      uncacheable_miss_scnd_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      imb_scnd_ff <= 31'h0;
    end else if (!(sel_hold_imb_scnd)) begin
      imb_scnd_ff <= io_ifc_fetch_addr_bf;
    end
    if (reset) begin
      ifu_bus_rid_ff <= 3'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rid_ff <= io_ifu_axi_rid;
    end
    if (reset) begin
      ifu_bus_rresp_ff <= 2'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rresp_ff <= io_ifu_axi_rresp;
    end
    if (reset) begin
      way_status_mb_ff <= 1'h0;
    end else if (_T_278) begin
      way_status_mb_ff <= way_status_mb_scnd_ff;
    end else if (_T_280) begin
      way_status_mb_ff <= replace_way_mb_any_0;
    end else if (!(miss_pending)) begin
      way_status_mb_ff <= way_status;
    end
    if (reset) begin
      tagv_mb_ff <= 2'h0;
    end else if (scnd_miss_req) begin
      tagv_mb_ff <= _T_290;
    end else if (!(miss_pending)) begin
      tagv_mb_ff <= _T_295;
    end
    reset_ic_ff <= _T_298 & _T_299;
    if (reset) begin
      fetch_uncacheable_ff <= 1'h0;
    end else begin
      fetch_uncacheable_ff <= io_ifc_fetch_uncacheable_bf;
    end
    if (reset) begin
      miss_addr <= 26'h0;
    end else if (_T_231) begin
      miss_addr <= imb_ff[30:5];
    end else if (scnd_miss_req_q) begin
      miss_addr <= imb_scnd_ff[30:5];
    end
    if (reset) begin
      ifc_region_acc_fault_f <= 1'h0;
    end else begin
      ifc_region_acc_fault_f <= io_ifc_region_acc_fault_bf;
    end
    if (reset) begin
      bus_rd_addr_count <= 3'h0;
    end else if (_T_2615) begin
      if (_T_231) begin
        bus_rd_addr_count <= imb_ff[4:2];
      end else if (scnd_miss_req_q) begin
        bus_rd_addr_count <= imb_scnd_ff[4:2];
      end else if (bus_cmd_sent) begin
        bus_rd_addr_count <= _T_2611;
      end
    end
    if (reset) begin
      ifu_bus_rdata_ff <= 64'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_rdata_ff <= io_ifu_axi_rdata;
    end
    if (reset) begin
      ic_miss_buff_data_0 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_0 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_1 <= 32'h0;
    end else if (write_fill_data_0) begin
      ic_miss_buff_data_1 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_2 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_2 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_3 <= 32'h0;
    end else if (write_fill_data_1) begin
      ic_miss_buff_data_3 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_4 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_4 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_5 <= 32'h0;
    end else if (write_fill_data_2) begin
      ic_miss_buff_data_5 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_6 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_6 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_7 <= 32'h0;
    end else if (write_fill_data_3) begin
      ic_miss_buff_data_7 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_8 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_8 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_9 <= 32'h0;
    end else if (write_fill_data_4) begin
      ic_miss_buff_data_9 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_10 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_10 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_11 <= 32'h0;
    end else if (write_fill_data_5) begin
      ic_miss_buff_data_11 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_12 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_12 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_13 <= 32'h0;
    end else if (write_fill_data_6) begin
      ic_miss_buff_data_13 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_miss_buff_data_14 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_14 <= io_ifu_axi_rdata[31:0];
    end
    if (reset) begin
      ic_miss_buff_data_15 <= 32'h0;
    end else if (write_fill_data_7) begin
      ic_miss_buff_data_15 <= io_ifu_axi_rdata[63:32];
    end
    if (reset) begin
      ic_debug_ict_array_sel_ff <= 1'h0;
    end else if (debug_c1_clken) begin
      ic_debug_ict_array_sel_ff <= ic_debug_ict_array_sel_in;
    end
    if (reset) begin
      ic_tag_valid_out_1_0 <= 1'h0;
    end else if (_T_5978) begin
      ic_tag_valid_out_1_0 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_1 <= 1'h0;
    end else if (_T_5995) begin
      ic_tag_valid_out_1_1 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_2 <= 1'h0;
    end else if (_T_6012) begin
      ic_tag_valid_out_1_2 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_3 <= 1'h0;
    end else if (_T_6029) begin
      ic_tag_valid_out_1_3 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_4 <= 1'h0;
    end else if (_T_6046) begin
      ic_tag_valid_out_1_4 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_5 <= 1'h0;
    end else if (_T_6063) begin
      ic_tag_valid_out_1_5 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_6 <= 1'h0;
    end else if (_T_6080) begin
      ic_tag_valid_out_1_6 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_7 <= 1'h0;
    end else if (_T_6097) begin
      ic_tag_valid_out_1_7 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_8 <= 1'h0;
    end else if (_T_6114) begin
      ic_tag_valid_out_1_8 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_9 <= 1'h0;
    end else if (_T_6131) begin
      ic_tag_valid_out_1_9 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_10 <= 1'h0;
    end else if (_T_6148) begin
      ic_tag_valid_out_1_10 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_11 <= 1'h0;
    end else if (_T_6165) begin
      ic_tag_valid_out_1_11 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_12 <= 1'h0;
    end else if (_T_6182) begin
      ic_tag_valid_out_1_12 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_13 <= 1'h0;
    end else if (_T_6199) begin
      ic_tag_valid_out_1_13 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_14 <= 1'h0;
    end else if (_T_6216) begin
      ic_tag_valid_out_1_14 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_15 <= 1'h0;
    end else if (_T_6233) begin
      ic_tag_valid_out_1_15 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_16 <= 1'h0;
    end else if (_T_6250) begin
      ic_tag_valid_out_1_16 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_17 <= 1'h0;
    end else if (_T_6267) begin
      ic_tag_valid_out_1_17 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_18 <= 1'h0;
    end else if (_T_6284) begin
      ic_tag_valid_out_1_18 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_19 <= 1'h0;
    end else if (_T_6301) begin
      ic_tag_valid_out_1_19 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_20 <= 1'h0;
    end else if (_T_6318) begin
      ic_tag_valid_out_1_20 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_21 <= 1'h0;
    end else if (_T_6335) begin
      ic_tag_valid_out_1_21 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_22 <= 1'h0;
    end else if (_T_6352) begin
      ic_tag_valid_out_1_22 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_23 <= 1'h0;
    end else if (_T_6369) begin
      ic_tag_valid_out_1_23 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_24 <= 1'h0;
    end else if (_T_6386) begin
      ic_tag_valid_out_1_24 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_25 <= 1'h0;
    end else if (_T_6403) begin
      ic_tag_valid_out_1_25 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_26 <= 1'h0;
    end else if (_T_6420) begin
      ic_tag_valid_out_1_26 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_27 <= 1'h0;
    end else if (_T_6437) begin
      ic_tag_valid_out_1_27 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_28 <= 1'h0;
    end else if (_T_6454) begin
      ic_tag_valid_out_1_28 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_29 <= 1'h0;
    end else if (_T_6471) begin
      ic_tag_valid_out_1_29 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_30 <= 1'h0;
    end else if (_T_6488) begin
      ic_tag_valid_out_1_30 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_31 <= 1'h0;
    end else if (_T_6505) begin
      ic_tag_valid_out_1_31 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_32 <= 1'h0;
    end else if (_T_7066) begin
      ic_tag_valid_out_1_32 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_33 <= 1'h0;
    end else if (_T_7083) begin
      ic_tag_valid_out_1_33 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_34 <= 1'h0;
    end else if (_T_7100) begin
      ic_tag_valid_out_1_34 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_35 <= 1'h0;
    end else if (_T_7117) begin
      ic_tag_valid_out_1_35 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_36 <= 1'h0;
    end else if (_T_7134) begin
      ic_tag_valid_out_1_36 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_37 <= 1'h0;
    end else if (_T_7151) begin
      ic_tag_valid_out_1_37 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_38 <= 1'h0;
    end else if (_T_7168) begin
      ic_tag_valid_out_1_38 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_39 <= 1'h0;
    end else if (_T_7185) begin
      ic_tag_valid_out_1_39 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_40 <= 1'h0;
    end else if (_T_7202) begin
      ic_tag_valid_out_1_40 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_41 <= 1'h0;
    end else if (_T_7219) begin
      ic_tag_valid_out_1_41 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_42 <= 1'h0;
    end else if (_T_7236) begin
      ic_tag_valid_out_1_42 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_43 <= 1'h0;
    end else if (_T_7253) begin
      ic_tag_valid_out_1_43 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_44 <= 1'h0;
    end else if (_T_7270) begin
      ic_tag_valid_out_1_44 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_45 <= 1'h0;
    end else if (_T_7287) begin
      ic_tag_valid_out_1_45 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_46 <= 1'h0;
    end else if (_T_7304) begin
      ic_tag_valid_out_1_46 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_47 <= 1'h0;
    end else if (_T_7321) begin
      ic_tag_valid_out_1_47 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_48 <= 1'h0;
    end else if (_T_7338) begin
      ic_tag_valid_out_1_48 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_49 <= 1'h0;
    end else if (_T_7355) begin
      ic_tag_valid_out_1_49 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_50 <= 1'h0;
    end else if (_T_7372) begin
      ic_tag_valid_out_1_50 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_51 <= 1'h0;
    end else if (_T_7389) begin
      ic_tag_valid_out_1_51 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_52 <= 1'h0;
    end else if (_T_7406) begin
      ic_tag_valid_out_1_52 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_53 <= 1'h0;
    end else if (_T_7423) begin
      ic_tag_valid_out_1_53 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_54 <= 1'h0;
    end else if (_T_7440) begin
      ic_tag_valid_out_1_54 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_55 <= 1'h0;
    end else if (_T_7457) begin
      ic_tag_valid_out_1_55 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_56 <= 1'h0;
    end else if (_T_7474) begin
      ic_tag_valid_out_1_56 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_57 <= 1'h0;
    end else if (_T_7491) begin
      ic_tag_valid_out_1_57 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_58 <= 1'h0;
    end else if (_T_7508) begin
      ic_tag_valid_out_1_58 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_59 <= 1'h0;
    end else if (_T_7525) begin
      ic_tag_valid_out_1_59 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_60 <= 1'h0;
    end else if (_T_7542) begin
      ic_tag_valid_out_1_60 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_61 <= 1'h0;
    end else if (_T_7559) begin
      ic_tag_valid_out_1_61 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_62 <= 1'h0;
    end else if (_T_7576) begin
      ic_tag_valid_out_1_62 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_63 <= 1'h0;
    end else if (_T_7593) begin
      ic_tag_valid_out_1_63 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_64 <= 1'h0;
    end else if (_T_8154) begin
      ic_tag_valid_out_1_64 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_65 <= 1'h0;
    end else if (_T_8171) begin
      ic_tag_valid_out_1_65 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_66 <= 1'h0;
    end else if (_T_8188) begin
      ic_tag_valid_out_1_66 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_67 <= 1'h0;
    end else if (_T_8205) begin
      ic_tag_valid_out_1_67 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_68 <= 1'h0;
    end else if (_T_8222) begin
      ic_tag_valid_out_1_68 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_69 <= 1'h0;
    end else if (_T_8239) begin
      ic_tag_valid_out_1_69 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_70 <= 1'h0;
    end else if (_T_8256) begin
      ic_tag_valid_out_1_70 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_71 <= 1'h0;
    end else if (_T_8273) begin
      ic_tag_valid_out_1_71 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_72 <= 1'h0;
    end else if (_T_8290) begin
      ic_tag_valid_out_1_72 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_73 <= 1'h0;
    end else if (_T_8307) begin
      ic_tag_valid_out_1_73 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_74 <= 1'h0;
    end else if (_T_8324) begin
      ic_tag_valid_out_1_74 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_75 <= 1'h0;
    end else if (_T_8341) begin
      ic_tag_valid_out_1_75 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_76 <= 1'h0;
    end else if (_T_8358) begin
      ic_tag_valid_out_1_76 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_77 <= 1'h0;
    end else if (_T_8375) begin
      ic_tag_valid_out_1_77 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_78 <= 1'h0;
    end else if (_T_8392) begin
      ic_tag_valid_out_1_78 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_79 <= 1'h0;
    end else if (_T_8409) begin
      ic_tag_valid_out_1_79 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_80 <= 1'h0;
    end else if (_T_8426) begin
      ic_tag_valid_out_1_80 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_81 <= 1'h0;
    end else if (_T_8443) begin
      ic_tag_valid_out_1_81 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_82 <= 1'h0;
    end else if (_T_8460) begin
      ic_tag_valid_out_1_82 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_83 <= 1'h0;
    end else if (_T_8477) begin
      ic_tag_valid_out_1_83 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_84 <= 1'h0;
    end else if (_T_8494) begin
      ic_tag_valid_out_1_84 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_85 <= 1'h0;
    end else if (_T_8511) begin
      ic_tag_valid_out_1_85 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_86 <= 1'h0;
    end else if (_T_8528) begin
      ic_tag_valid_out_1_86 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_87 <= 1'h0;
    end else if (_T_8545) begin
      ic_tag_valid_out_1_87 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_88 <= 1'h0;
    end else if (_T_8562) begin
      ic_tag_valid_out_1_88 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_89 <= 1'h0;
    end else if (_T_8579) begin
      ic_tag_valid_out_1_89 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_90 <= 1'h0;
    end else if (_T_8596) begin
      ic_tag_valid_out_1_90 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_91 <= 1'h0;
    end else if (_T_8613) begin
      ic_tag_valid_out_1_91 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_92 <= 1'h0;
    end else if (_T_8630) begin
      ic_tag_valid_out_1_92 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_93 <= 1'h0;
    end else if (_T_8647) begin
      ic_tag_valid_out_1_93 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_94 <= 1'h0;
    end else if (_T_8664) begin
      ic_tag_valid_out_1_94 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_95 <= 1'h0;
    end else if (_T_8681) begin
      ic_tag_valid_out_1_95 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_96 <= 1'h0;
    end else if (_T_9242) begin
      ic_tag_valid_out_1_96 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_97 <= 1'h0;
    end else if (_T_9259) begin
      ic_tag_valid_out_1_97 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_98 <= 1'h0;
    end else if (_T_9276) begin
      ic_tag_valid_out_1_98 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_99 <= 1'h0;
    end else if (_T_9293) begin
      ic_tag_valid_out_1_99 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_100 <= 1'h0;
    end else if (_T_9310) begin
      ic_tag_valid_out_1_100 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_101 <= 1'h0;
    end else if (_T_9327) begin
      ic_tag_valid_out_1_101 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_102 <= 1'h0;
    end else if (_T_9344) begin
      ic_tag_valid_out_1_102 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_103 <= 1'h0;
    end else if (_T_9361) begin
      ic_tag_valid_out_1_103 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_104 <= 1'h0;
    end else if (_T_9378) begin
      ic_tag_valid_out_1_104 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_105 <= 1'h0;
    end else if (_T_9395) begin
      ic_tag_valid_out_1_105 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_106 <= 1'h0;
    end else if (_T_9412) begin
      ic_tag_valid_out_1_106 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_107 <= 1'h0;
    end else if (_T_9429) begin
      ic_tag_valid_out_1_107 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_108 <= 1'h0;
    end else if (_T_9446) begin
      ic_tag_valid_out_1_108 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_109 <= 1'h0;
    end else if (_T_9463) begin
      ic_tag_valid_out_1_109 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_110 <= 1'h0;
    end else if (_T_9480) begin
      ic_tag_valid_out_1_110 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_111 <= 1'h0;
    end else if (_T_9497) begin
      ic_tag_valid_out_1_111 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_112 <= 1'h0;
    end else if (_T_9514) begin
      ic_tag_valid_out_1_112 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_113 <= 1'h0;
    end else if (_T_9531) begin
      ic_tag_valid_out_1_113 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_114 <= 1'h0;
    end else if (_T_9548) begin
      ic_tag_valid_out_1_114 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_115 <= 1'h0;
    end else if (_T_9565) begin
      ic_tag_valid_out_1_115 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_116 <= 1'h0;
    end else if (_T_9582) begin
      ic_tag_valid_out_1_116 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_117 <= 1'h0;
    end else if (_T_9599) begin
      ic_tag_valid_out_1_117 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_118 <= 1'h0;
    end else if (_T_9616) begin
      ic_tag_valid_out_1_118 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_119 <= 1'h0;
    end else if (_T_9633) begin
      ic_tag_valid_out_1_119 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_120 <= 1'h0;
    end else if (_T_9650) begin
      ic_tag_valid_out_1_120 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_121 <= 1'h0;
    end else if (_T_9667) begin
      ic_tag_valid_out_1_121 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_122 <= 1'h0;
    end else if (_T_9684) begin
      ic_tag_valid_out_1_122 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_123 <= 1'h0;
    end else if (_T_9701) begin
      ic_tag_valid_out_1_123 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_124 <= 1'h0;
    end else if (_T_9718) begin
      ic_tag_valid_out_1_124 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_125 <= 1'h0;
    end else if (_T_9735) begin
      ic_tag_valid_out_1_125 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_126 <= 1'h0;
    end else if (_T_9752) begin
      ic_tag_valid_out_1_126 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_1_127 <= 1'h0;
    end else if (_T_9769) begin
      ic_tag_valid_out_1_127 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_0 <= 1'h0;
    end else if (_T_5434) begin
      ic_tag_valid_out_0_0 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_1 <= 1'h0;
    end else if (_T_5451) begin
      ic_tag_valid_out_0_1 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_2 <= 1'h0;
    end else if (_T_5468) begin
      ic_tag_valid_out_0_2 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_3 <= 1'h0;
    end else if (_T_5485) begin
      ic_tag_valid_out_0_3 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_4 <= 1'h0;
    end else if (_T_5502) begin
      ic_tag_valid_out_0_4 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_5 <= 1'h0;
    end else if (_T_5519) begin
      ic_tag_valid_out_0_5 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_6 <= 1'h0;
    end else if (_T_5536) begin
      ic_tag_valid_out_0_6 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_7 <= 1'h0;
    end else if (_T_5553) begin
      ic_tag_valid_out_0_7 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_8 <= 1'h0;
    end else if (_T_5570) begin
      ic_tag_valid_out_0_8 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_9 <= 1'h0;
    end else if (_T_5587) begin
      ic_tag_valid_out_0_9 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_10 <= 1'h0;
    end else if (_T_5604) begin
      ic_tag_valid_out_0_10 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_11 <= 1'h0;
    end else if (_T_5621) begin
      ic_tag_valid_out_0_11 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_12 <= 1'h0;
    end else if (_T_5638) begin
      ic_tag_valid_out_0_12 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_13 <= 1'h0;
    end else if (_T_5655) begin
      ic_tag_valid_out_0_13 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_14 <= 1'h0;
    end else if (_T_5672) begin
      ic_tag_valid_out_0_14 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_15 <= 1'h0;
    end else if (_T_5689) begin
      ic_tag_valid_out_0_15 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_16 <= 1'h0;
    end else if (_T_5706) begin
      ic_tag_valid_out_0_16 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_17 <= 1'h0;
    end else if (_T_5723) begin
      ic_tag_valid_out_0_17 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_18 <= 1'h0;
    end else if (_T_5740) begin
      ic_tag_valid_out_0_18 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_19 <= 1'h0;
    end else if (_T_5757) begin
      ic_tag_valid_out_0_19 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_20 <= 1'h0;
    end else if (_T_5774) begin
      ic_tag_valid_out_0_20 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_21 <= 1'h0;
    end else if (_T_5791) begin
      ic_tag_valid_out_0_21 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_22 <= 1'h0;
    end else if (_T_5808) begin
      ic_tag_valid_out_0_22 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_23 <= 1'h0;
    end else if (_T_5825) begin
      ic_tag_valid_out_0_23 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_24 <= 1'h0;
    end else if (_T_5842) begin
      ic_tag_valid_out_0_24 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_25 <= 1'h0;
    end else if (_T_5859) begin
      ic_tag_valid_out_0_25 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_26 <= 1'h0;
    end else if (_T_5876) begin
      ic_tag_valid_out_0_26 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_27 <= 1'h0;
    end else if (_T_5893) begin
      ic_tag_valid_out_0_27 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_28 <= 1'h0;
    end else if (_T_5910) begin
      ic_tag_valid_out_0_28 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_29 <= 1'h0;
    end else if (_T_5927) begin
      ic_tag_valid_out_0_29 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_30 <= 1'h0;
    end else if (_T_5944) begin
      ic_tag_valid_out_0_30 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_31 <= 1'h0;
    end else if (_T_5961) begin
      ic_tag_valid_out_0_31 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_32 <= 1'h0;
    end else if (_T_6522) begin
      ic_tag_valid_out_0_32 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_33 <= 1'h0;
    end else if (_T_6539) begin
      ic_tag_valid_out_0_33 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_34 <= 1'h0;
    end else if (_T_6556) begin
      ic_tag_valid_out_0_34 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_35 <= 1'h0;
    end else if (_T_6573) begin
      ic_tag_valid_out_0_35 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_36 <= 1'h0;
    end else if (_T_6590) begin
      ic_tag_valid_out_0_36 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_37 <= 1'h0;
    end else if (_T_6607) begin
      ic_tag_valid_out_0_37 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_38 <= 1'h0;
    end else if (_T_6624) begin
      ic_tag_valid_out_0_38 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_39 <= 1'h0;
    end else if (_T_6641) begin
      ic_tag_valid_out_0_39 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_40 <= 1'h0;
    end else if (_T_6658) begin
      ic_tag_valid_out_0_40 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_41 <= 1'h0;
    end else if (_T_6675) begin
      ic_tag_valid_out_0_41 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_42 <= 1'h0;
    end else if (_T_6692) begin
      ic_tag_valid_out_0_42 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_43 <= 1'h0;
    end else if (_T_6709) begin
      ic_tag_valid_out_0_43 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_44 <= 1'h0;
    end else if (_T_6726) begin
      ic_tag_valid_out_0_44 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_45 <= 1'h0;
    end else if (_T_6743) begin
      ic_tag_valid_out_0_45 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_46 <= 1'h0;
    end else if (_T_6760) begin
      ic_tag_valid_out_0_46 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_47 <= 1'h0;
    end else if (_T_6777) begin
      ic_tag_valid_out_0_47 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_48 <= 1'h0;
    end else if (_T_6794) begin
      ic_tag_valid_out_0_48 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_49 <= 1'h0;
    end else if (_T_6811) begin
      ic_tag_valid_out_0_49 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_50 <= 1'h0;
    end else if (_T_6828) begin
      ic_tag_valid_out_0_50 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_51 <= 1'h0;
    end else if (_T_6845) begin
      ic_tag_valid_out_0_51 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_52 <= 1'h0;
    end else if (_T_6862) begin
      ic_tag_valid_out_0_52 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_53 <= 1'h0;
    end else if (_T_6879) begin
      ic_tag_valid_out_0_53 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_54 <= 1'h0;
    end else if (_T_6896) begin
      ic_tag_valid_out_0_54 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_55 <= 1'h0;
    end else if (_T_6913) begin
      ic_tag_valid_out_0_55 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_56 <= 1'h0;
    end else if (_T_6930) begin
      ic_tag_valid_out_0_56 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_57 <= 1'h0;
    end else if (_T_6947) begin
      ic_tag_valid_out_0_57 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_58 <= 1'h0;
    end else if (_T_6964) begin
      ic_tag_valid_out_0_58 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_59 <= 1'h0;
    end else if (_T_6981) begin
      ic_tag_valid_out_0_59 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_60 <= 1'h0;
    end else if (_T_6998) begin
      ic_tag_valid_out_0_60 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_61 <= 1'h0;
    end else if (_T_7015) begin
      ic_tag_valid_out_0_61 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_62 <= 1'h0;
    end else if (_T_7032) begin
      ic_tag_valid_out_0_62 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_63 <= 1'h0;
    end else if (_T_7049) begin
      ic_tag_valid_out_0_63 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_64 <= 1'h0;
    end else if (_T_7610) begin
      ic_tag_valid_out_0_64 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_65 <= 1'h0;
    end else if (_T_7627) begin
      ic_tag_valid_out_0_65 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_66 <= 1'h0;
    end else if (_T_7644) begin
      ic_tag_valid_out_0_66 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_67 <= 1'h0;
    end else if (_T_7661) begin
      ic_tag_valid_out_0_67 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_68 <= 1'h0;
    end else if (_T_7678) begin
      ic_tag_valid_out_0_68 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_69 <= 1'h0;
    end else if (_T_7695) begin
      ic_tag_valid_out_0_69 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_70 <= 1'h0;
    end else if (_T_7712) begin
      ic_tag_valid_out_0_70 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_71 <= 1'h0;
    end else if (_T_7729) begin
      ic_tag_valid_out_0_71 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_72 <= 1'h0;
    end else if (_T_7746) begin
      ic_tag_valid_out_0_72 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_73 <= 1'h0;
    end else if (_T_7763) begin
      ic_tag_valid_out_0_73 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_74 <= 1'h0;
    end else if (_T_7780) begin
      ic_tag_valid_out_0_74 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_75 <= 1'h0;
    end else if (_T_7797) begin
      ic_tag_valid_out_0_75 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_76 <= 1'h0;
    end else if (_T_7814) begin
      ic_tag_valid_out_0_76 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_77 <= 1'h0;
    end else if (_T_7831) begin
      ic_tag_valid_out_0_77 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_78 <= 1'h0;
    end else if (_T_7848) begin
      ic_tag_valid_out_0_78 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_79 <= 1'h0;
    end else if (_T_7865) begin
      ic_tag_valid_out_0_79 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_80 <= 1'h0;
    end else if (_T_7882) begin
      ic_tag_valid_out_0_80 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_81 <= 1'h0;
    end else if (_T_7899) begin
      ic_tag_valid_out_0_81 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_82 <= 1'h0;
    end else if (_T_7916) begin
      ic_tag_valid_out_0_82 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_83 <= 1'h0;
    end else if (_T_7933) begin
      ic_tag_valid_out_0_83 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_84 <= 1'h0;
    end else if (_T_7950) begin
      ic_tag_valid_out_0_84 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_85 <= 1'h0;
    end else if (_T_7967) begin
      ic_tag_valid_out_0_85 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_86 <= 1'h0;
    end else if (_T_7984) begin
      ic_tag_valid_out_0_86 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_87 <= 1'h0;
    end else if (_T_8001) begin
      ic_tag_valid_out_0_87 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_88 <= 1'h0;
    end else if (_T_8018) begin
      ic_tag_valid_out_0_88 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_89 <= 1'h0;
    end else if (_T_8035) begin
      ic_tag_valid_out_0_89 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_90 <= 1'h0;
    end else if (_T_8052) begin
      ic_tag_valid_out_0_90 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_91 <= 1'h0;
    end else if (_T_8069) begin
      ic_tag_valid_out_0_91 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_92 <= 1'h0;
    end else if (_T_8086) begin
      ic_tag_valid_out_0_92 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_93 <= 1'h0;
    end else if (_T_8103) begin
      ic_tag_valid_out_0_93 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_94 <= 1'h0;
    end else if (_T_8120) begin
      ic_tag_valid_out_0_94 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_95 <= 1'h0;
    end else if (_T_8137) begin
      ic_tag_valid_out_0_95 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_96 <= 1'h0;
    end else if (_T_8698) begin
      ic_tag_valid_out_0_96 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_97 <= 1'h0;
    end else if (_T_8715) begin
      ic_tag_valid_out_0_97 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_98 <= 1'h0;
    end else if (_T_8732) begin
      ic_tag_valid_out_0_98 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_99 <= 1'h0;
    end else if (_T_8749) begin
      ic_tag_valid_out_0_99 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_100 <= 1'h0;
    end else if (_T_8766) begin
      ic_tag_valid_out_0_100 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_101 <= 1'h0;
    end else if (_T_8783) begin
      ic_tag_valid_out_0_101 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_102 <= 1'h0;
    end else if (_T_8800) begin
      ic_tag_valid_out_0_102 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_103 <= 1'h0;
    end else if (_T_8817) begin
      ic_tag_valid_out_0_103 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_104 <= 1'h0;
    end else if (_T_8834) begin
      ic_tag_valid_out_0_104 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_105 <= 1'h0;
    end else if (_T_8851) begin
      ic_tag_valid_out_0_105 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_106 <= 1'h0;
    end else if (_T_8868) begin
      ic_tag_valid_out_0_106 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_107 <= 1'h0;
    end else if (_T_8885) begin
      ic_tag_valid_out_0_107 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_108 <= 1'h0;
    end else if (_T_8902) begin
      ic_tag_valid_out_0_108 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_109 <= 1'h0;
    end else if (_T_8919) begin
      ic_tag_valid_out_0_109 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_110 <= 1'h0;
    end else if (_T_8936) begin
      ic_tag_valid_out_0_110 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_111 <= 1'h0;
    end else if (_T_8953) begin
      ic_tag_valid_out_0_111 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_112 <= 1'h0;
    end else if (_T_8970) begin
      ic_tag_valid_out_0_112 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_113 <= 1'h0;
    end else if (_T_8987) begin
      ic_tag_valid_out_0_113 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_114 <= 1'h0;
    end else if (_T_9004) begin
      ic_tag_valid_out_0_114 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_115 <= 1'h0;
    end else if (_T_9021) begin
      ic_tag_valid_out_0_115 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_116 <= 1'h0;
    end else if (_T_9038) begin
      ic_tag_valid_out_0_116 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_117 <= 1'h0;
    end else if (_T_9055) begin
      ic_tag_valid_out_0_117 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_118 <= 1'h0;
    end else if (_T_9072) begin
      ic_tag_valid_out_0_118 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_119 <= 1'h0;
    end else if (_T_9089) begin
      ic_tag_valid_out_0_119 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_120 <= 1'h0;
    end else if (_T_9106) begin
      ic_tag_valid_out_0_120 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_121 <= 1'h0;
    end else if (_T_9123) begin
      ic_tag_valid_out_0_121 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_122 <= 1'h0;
    end else if (_T_9140) begin
      ic_tag_valid_out_0_122 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_123 <= 1'h0;
    end else if (_T_9157) begin
      ic_tag_valid_out_0_123 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_124 <= 1'h0;
    end else if (_T_9174) begin
      ic_tag_valid_out_0_124 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_125 <= 1'h0;
    end else if (_T_9191) begin
      ic_tag_valid_out_0_125 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_126 <= 1'h0;
    end else if (_T_9208) begin
      ic_tag_valid_out_0_126 <= _T_5424;
    end
    if (reset) begin
      ic_tag_valid_out_0_127 <= 1'h0;
    end else if (_T_9225) begin
      ic_tag_valid_out_0_127 <= _T_5424;
    end
    if (reset) begin
      ic_debug_way_ff <= 2'h0;
    end else if (debug_c1_clken) begin
      ic_debug_way_ff <= io_ic_debug_way;
    end
    if (reset) begin
      _T_1209 <= 71'h0;
    end else if (ic_debug_rd_en_ff) begin
      if (ic_debug_ict_array_sel_ff) begin
        _T_1209 <= {{5'd0}, _T_1208};
      end else begin
        _T_1209 <= io_ic_debug_rd_data;
      end
    end
    if (reset) begin
      ifu_bus_cmd_valid <= 1'h0;
    end else if (_T_2564) begin
      ifu_bus_cmd_valid <= ifc_bus_ic_req_ff_in;
    end
    if (reset) begin
      bus_cmd_beat_count <= 3'h0;
    end else if (_T_2639) begin
      bus_cmd_beat_count <= bus_new_cmd_beat_count;
    end
    if (reset) begin
      ifu_bus_arready_unq_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arready_unq_ff <= io_ifu_axi_arready;
    end
    if (reset) begin
      ifu_bus_arvalid_ff <= 1'h0;
    end else if (io_ifu_bus_clk_en) begin
      ifu_bus_arvalid_ff <= io_ifu_axi_arvalid;
    end
  end
  always @(posedge io_free_clk) begin
    if (reset) begin
      scnd_miss_req_q <= 1'h0;
    end else begin
      scnd_miss_req_q <= scnd_miss_req_in;
    end
    if (reset) begin
      iccm_dma_rvalid_in <= 1'h0;
    end else begin
      iccm_dma_rvalid_in <= _T_2683;
    end
    if (reset) begin
      dma_iccm_req_f <= 1'h0;
    end else begin
      dma_iccm_req_f <= io_dma_iccm_req;
    end
    if (reset) begin
      perr_state <= 3'h0;
    end else if (perr_state_en) begin
      if (_T_2465) begin
        if (io_iccm_dma_sb_error) begin
          perr_state <= 3'h4;
        end else if (_T_2467) begin
          perr_state <= 3'h1;
        end else begin
          perr_state <= 3'h2;
        end
      end else if (_T_2477) begin
        perr_state <= 3'h0;
      end else if (_T_2480) begin
        if (_T_2482) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else if (_T_2486) begin
        if (io_dec_tlu_force_halt) begin
          perr_state <= 3'h0;
        end else begin
          perr_state <= 3'h3;
        end
      end else begin
        perr_state <= 3'h0;
      end
    end
    if (reset) begin
      err_stop_state <= 2'h0;
    end else if (err_stop_state_en) begin
      if (_T_2490) begin
        err_stop_state <= 2'h1;
      end else if (_T_2495) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (_T_2518) begin
          err_stop_state <= 2'h3;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h2;
        end else begin
          err_stop_state <= 2'h1;
        end
      end else if (_T_2522) begin
        if (_T_2497) begin
          err_stop_state <= 2'h0;
        end else if (io_ifu_fetch_val[0]) begin
          err_stop_state <= 2'h3;
        end else begin
          err_stop_state <= 2'h2;
        end
      end else if (_T_2539) begin
        if (_T_2543) begin
          err_stop_state <= 2'h0;
        end else if (io_dec_tlu_flush_err_wb) begin
          err_stop_state <= 2'h1;
        end else begin
          err_stop_state <= 2'h3;
        end
      end else begin
        err_stop_state <= 2'h0;
      end
    end
    if (reset) begin
      bus_ifu_bus_clk_en_ff <= 1'h0;
    end else begin
      bus_ifu_bus_clk_en_ff <= io_ifu_bus_clk_en;
    end
    if (reset) begin
      bus_data_beat_count <= 3'h0;
    end else begin
      bus_data_beat_count <= bus_new_data_beat_count;
    end
    if (reset) begin
      ic_miss_buff_data_valid <= 8'h0;
    end else begin
      ic_miss_buff_data_valid <= _T_1368;
    end
    if (reset) begin
      last_data_recieved_ff <= 1'h0;
    end else begin
      last_data_recieved_ff <= last_data_recieved_in;
    end
    if (reset) begin
      sel_mb_addr_ff <= 1'h0;
    end else begin
      sel_mb_addr_ff <= sel_mb_addr;
    end
    if (reset) begin
      ifu_ic_rw_int_addr_ff <= 7'h0;
    end else if (_T_4147) begin
      ifu_ic_rw_int_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_ic_rw_int_addr_ff <= ifu_ic_rw_int_addr[11:5];
    end
    if (reset) begin
      ifu_wr_data_comb_err_ff <= 1'h0;
    end else begin
      ifu_wr_data_comb_err_ff <= ifu_wr_cumulative_err;
    end
    if (reset) begin
      ic_act_miss_f_delayed <= 1'h0;
    end else begin
      ic_act_miss_f_delayed <= ic_act_miss_f;
    end
    if (reset) begin
      ic_crit_wd_rdy_new_ff <= 1'h0;
    end else begin
      ic_crit_wd_rdy_new_ff <= ic_crit_wd_rdy_new_in;
    end
    if (reset) begin
      ic_miss_buff_data_error <= 8'h0;
    end else begin
      ic_miss_buff_data_error <= _T_1408;
    end
    if (reset) begin
      ic_debug_rd_en_ff <= 1'h0;
    end else begin
      ic_debug_rd_en_ff <= io_ic_debug_rd_en;
    end
    if (reset) begin
      ifc_dma_access_ok_prev <= 1'h0;
    end else begin
      ifc_dma_access_ok_prev <= ifc_dma_access_ok_d;
    end
    if (reset) begin
      iccm_ecc_corr_data_ff <= 39'h0;
    end else if (iccm_ecc_write_status) begin
      iccm_ecc_corr_data_ff <= _T_4082;
    end
    if (reset) begin
      dma_mem_addr_ff <= 2'h0;
    end else begin
      dma_mem_addr_ff <= io_dma_mem_addr[3:2];
    end
    if (reset) begin
      dma_mem_tag_ff <= 3'h0;
    end else begin
      dma_mem_tag_ff <= io_dma_mem_tag;
    end
    if (reset) begin
      iccm_dma_rtag_temp <= 3'h0;
    end else begin
      iccm_dma_rtag_temp <= dma_mem_tag_ff;
    end
    if (reset) begin
      iccm_dma_rvalid_temp <= 1'h0;
    end else begin
      iccm_dma_rvalid_temp <= iccm_dma_rvalid_in;
    end
    if (reset) begin
      iccm_dma_rdata_temp <= 64'h0;
    end else if (iccm_dma_ecc_error_in) begin
      iccm_dma_rdata_temp <= _T_3257;
    end else begin
      iccm_dma_rdata_temp <= _T_3258;
    end
    if (reset) begin
      iccm_ecc_corr_index_ff <= 14'h0;
    end else if (iccm_ecc_write_status) begin
      if (iccm_single_ecc_error[0]) begin
        iccm_ecc_corr_index_ff <= iccm_rw_addr_f;
      end else begin
        iccm_ecc_corr_index_ff <= _T_4078;
      end
    end
    if (reset) begin
      iccm_rd_ecc_single_err_ff <= 1'h0;
    end else begin
      iccm_rd_ecc_single_err_ff <= iccm_rd_ecc_single_err_hold_in;
    end
    if (reset) begin
      iccm_rw_addr_f <= 14'h0;
    end else begin
      iccm_rw_addr_f <= io_iccm_rw_addr[14:1];
    end
    if (reset) begin
      ifu_status_wr_addr_ff <= 7'h0;
    end else if (_T_4147) begin
      ifu_status_wr_addr_ff <= io_ic_debug_addr[9:3];
    end else begin
      ifu_status_wr_addr_ff <= ifu_status_wr_addr[11:5];
    end
    if (reset) begin
      way_status_wr_en_ff <= 1'h0;
    end else begin
      way_status_wr_en_ff <= way_status_wr_en_w_debug;
    end
    if (reset) begin
      way_status_new_ff <= 1'h0;
    end else if (_T_4150) begin
      way_status_new_ff <= io_ic_debug_wr_data[4];
    end else if (_T_10559) begin
      way_status_new_ff <= replace_way_mb_any_0;
    end else begin
      way_status_new_ff <= way_status_hit_new;
    end
    if (reset) begin
      ifu_tag_wren_ff <= 2'h0;
    end else begin
      ifu_tag_wren_ff <= ifu_tag_wren_w_debug;
    end
    if (reset) begin
      ic_valid_ff <= 1'h0;
    end else if (_T_4150) begin
      ic_valid_ff <= io_ic_debug_wr_data[0];
    end else begin
      ic_valid_ff <= ic_valid;
    end
    if (reset) begin
      _T_10611 <= 1'h0;
    end else if (ic_debug_rd_en_ff) begin
      _T_10611 <= ic_debug_rd_en_ff;
    end
  end
  always @(posedge io_active_clk) begin
    if (reset) begin
      reset_all_tags <= 1'h0;
    end else begin
      reset_all_tags <= io_dec_tlu_fence_i_wb;
    end
    if (reset) begin
      perr_ic_index_ff <= 7'h0;
    end else if (perr_sb_write_status) begin
      perr_ic_index_ff <= ifu_ic_rw_int_addr_ff;
    end
    if (reset) begin
      dma_sb_err_state_ff <= 1'h0;
    end else begin
      dma_sb_err_state_ff <= _T_7;
    end
    if (reset) begin
      _T_10581 <= 1'h0;
    end else begin
      _T_10581 <= ic_act_miss_f;
    end
    if (reset) begin
      _T_10582 <= 1'h0;
    end else begin
      _T_10582 <= ic_act_hit_f;
    end
    if (reset) begin
      _T_10583 <= 1'h0;
    end else begin
      _T_10583 <= ifc_bus_acc_fault_f;
    end
    if (reset) begin
      _T_10587 <= 1'h0;
    end else begin
      _T_10587 <= _T_10586;
    end
    if (reset) begin
      _T_10588 <= 1'h0;
    end else begin
      _T_10588 <= bus_cmd_sent;
    end
  end
endmodule
